`timescale 1ns / 1ps

//

module divider_8x8(CLK, A, B, OUT);
input wire CLK;
input wire [7:0] A;
input wire [7:0] B;
output reg [7:0] OUT;

always @(posedge CLK)
case ({A, B})
    16'b00000000_00000000 : OUT <= 0;  //0 / 0 = 0
    16'b00000000_00000001 : OUT <= 0;  //0 / 1 = 0
    16'b00000000_00000010 : OUT <= 0;  //0 / 2 = 0
    16'b00000000_00000011 : OUT <= 0;  //0 / 3 = 0
    16'b00000000_00000100 : OUT <= 0;  //0 / 4 = 0
    16'b00000000_00000101 : OUT <= 0;  //0 / 5 = 0
    16'b00000000_00000110 : OUT <= 0;  //0 / 6 = 0
    16'b00000000_00000111 : OUT <= 0;  //0 / 7 = 0
    16'b00000000_00001000 : OUT <= 0;  //0 / 8 = 0
    16'b00000000_00001001 : OUT <= 0;  //0 / 9 = 0
    16'b00000000_00001010 : OUT <= 0;  //0 / 10 = 0
    16'b00000000_00001011 : OUT <= 0;  //0 / 11 = 0
    16'b00000000_00001100 : OUT <= 0;  //0 / 12 = 0
    16'b00000000_00001101 : OUT <= 0;  //0 / 13 = 0
    16'b00000000_00001110 : OUT <= 0;  //0 / 14 = 0
    16'b00000000_00001111 : OUT <= 0;  //0 / 15 = 0
    16'b00000000_00010000 : OUT <= 0;  //0 / 16 = 0
    16'b00000000_00010001 : OUT <= 0;  //0 / 17 = 0
    16'b00000000_00010010 : OUT <= 0;  //0 / 18 = 0
    16'b00000000_00010011 : OUT <= 0;  //0 / 19 = 0
    16'b00000000_00010100 : OUT <= 0;  //0 / 20 = 0
    16'b00000000_00010101 : OUT <= 0;  //0 / 21 = 0
    16'b00000000_00010110 : OUT <= 0;  //0 / 22 = 0
    16'b00000000_00010111 : OUT <= 0;  //0 / 23 = 0
    16'b00000000_00011000 : OUT <= 0;  //0 / 24 = 0
    16'b00000000_00011001 : OUT <= 0;  //0 / 25 = 0
    16'b00000000_00011010 : OUT <= 0;  //0 / 26 = 0
    16'b00000000_00011011 : OUT <= 0;  //0 / 27 = 0
    16'b00000000_00011100 : OUT <= 0;  //0 / 28 = 0
    16'b00000000_00011101 : OUT <= 0;  //0 / 29 = 0
    16'b00000000_00011110 : OUT <= 0;  //0 / 30 = 0
    16'b00000000_00011111 : OUT <= 0;  //0 / 31 = 0
    16'b00000000_00100000 : OUT <= 0;  //0 / 32 = 0
    16'b00000000_00100001 : OUT <= 0;  //0 / 33 = 0
    16'b00000000_00100010 : OUT <= 0;  //0 / 34 = 0
    16'b00000000_00100011 : OUT <= 0;  //0 / 35 = 0
    16'b00000000_00100100 : OUT <= 0;  //0 / 36 = 0
    16'b00000000_00100101 : OUT <= 0;  //0 / 37 = 0
    16'b00000000_00100110 : OUT <= 0;  //0 / 38 = 0
    16'b00000000_00100111 : OUT <= 0;  //0 / 39 = 0
    16'b00000000_00101000 : OUT <= 0;  //0 / 40 = 0
    16'b00000000_00101001 : OUT <= 0;  //0 / 41 = 0
    16'b00000000_00101010 : OUT <= 0;  //0 / 42 = 0
    16'b00000000_00101011 : OUT <= 0;  //0 / 43 = 0
    16'b00000000_00101100 : OUT <= 0;  //0 / 44 = 0
    16'b00000000_00101101 : OUT <= 0;  //0 / 45 = 0
    16'b00000000_00101110 : OUT <= 0;  //0 / 46 = 0
    16'b00000000_00101111 : OUT <= 0;  //0 / 47 = 0
    16'b00000000_00110000 : OUT <= 0;  //0 / 48 = 0
    16'b00000000_00110001 : OUT <= 0;  //0 / 49 = 0
    16'b00000000_00110010 : OUT <= 0;  //0 / 50 = 0
    16'b00000000_00110011 : OUT <= 0;  //0 / 51 = 0
    16'b00000000_00110100 : OUT <= 0;  //0 / 52 = 0
    16'b00000000_00110101 : OUT <= 0;  //0 / 53 = 0
    16'b00000000_00110110 : OUT <= 0;  //0 / 54 = 0
    16'b00000000_00110111 : OUT <= 0;  //0 / 55 = 0
    16'b00000000_00111000 : OUT <= 0;  //0 / 56 = 0
    16'b00000000_00111001 : OUT <= 0;  //0 / 57 = 0
    16'b00000000_00111010 : OUT <= 0;  //0 / 58 = 0
    16'b00000000_00111011 : OUT <= 0;  //0 / 59 = 0
    16'b00000000_00111100 : OUT <= 0;  //0 / 60 = 0
    16'b00000000_00111101 : OUT <= 0;  //0 / 61 = 0
    16'b00000000_00111110 : OUT <= 0;  //0 / 62 = 0
    16'b00000000_00111111 : OUT <= 0;  //0 / 63 = 0
    16'b00000000_01000000 : OUT <= 0;  //0 / 64 = 0
    16'b00000000_01000001 : OUT <= 0;  //0 / 65 = 0
    16'b00000000_01000010 : OUT <= 0;  //0 / 66 = 0
    16'b00000000_01000011 : OUT <= 0;  //0 / 67 = 0
    16'b00000000_01000100 : OUT <= 0;  //0 / 68 = 0
    16'b00000000_01000101 : OUT <= 0;  //0 / 69 = 0
    16'b00000000_01000110 : OUT <= 0;  //0 / 70 = 0
    16'b00000000_01000111 : OUT <= 0;  //0 / 71 = 0
    16'b00000000_01001000 : OUT <= 0;  //0 / 72 = 0
    16'b00000000_01001001 : OUT <= 0;  //0 / 73 = 0
    16'b00000000_01001010 : OUT <= 0;  //0 / 74 = 0
    16'b00000000_01001011 : OUT <= 0;  //0 / 75 = 0
    16'b00000000_01001100 : OUT <= 0;  //0 / 76 = 0
    16'b00000000_01001101 : OUT <= 0;  //0 / 77 = 0
    16'b00000000_01001110 : OUT <= 0;  //0 / 78 = 0
    16'b00000000_01001111 : OUT <= 0;  //0 / 79 = 0
    16'b00000000_01010000 : OUT <= 0;  //0 / 80 = 0
    16'b00000000_01010001 : OUT <= 0;  //0 / 81 = 0
    16'b00000000_01010010 : OUT <= 0;  //0 / 82 = 0
    16'b00000000_01010011 : OUT <= 0;  //0 / 83 = 0
    16'b00000000_01010100 : OUT <= 0;  //0 / 84 = 0
    16'b00000000_01010101 : OUT <= 0;  //0 / 85 = 0
    16'b00000000_01010110 : OUT <= 0;  //0 / 86 = 0
    16'b00000000_01010111 : OUT <= 0;  //0 / 87 = 0
    16'b00000000_01011000 : OUT <= 0;  //0 / 88 = 0
    16'b00000000_01011001 : OUT <= 0;  //0 / 89 = 0
    16'b00000000_01011010 : OUT <= 0;  //0 / 90 = 0
    16'b00000000_01011011 : OUT <= 0;  //0 / 91 = 0
    16'b00000000_01011100 : OUT <= 0;  //0 / 92 = 0
    16'b00000000_01011101 : OUT <= 0;  //0 / 93 = 0
    16'b00000000_01011110 : OUT <= 0;  //0 / 94 = 0
    16'b00000000_01011111 : OUT <= 0;  //0 / 95 = 0
    16'b00000000_01100000 : OUT <= 0;  //0 / 96 = 0
    16'b00000000_01100001 : OUT <= 0;  //0 / 97 = 0
    16'b00000000_01100010 : OUT <= 0;  //0 / 98 = 0
    16'b00000000_01100011 : OUT <= 0;  //0 / 99 = 0
    16'b00000000_01100100 : OUT <= 0;  //0 / 100 = 0
    16'b00000000_01100101 : OUT <= 0;  //0 / 101 = 0
    16'b00000000_01100110 : OUT <= 0;  //0 / 102 = 0
    16'b00000000_01100111 : OUT <= 0;  //0 / 103 = 0
    16'b00000000_01101000 : OUT <= 0;  //0 / 104 = 0
    16'b00000000_01101001 : OUT <= 0;  //0 / 105 = 0
    16'b00000000_01101010 : OUT <= 0;  //0 / 106 = 0
    16'b00000000_01101011 : OUT <= 0;  //0 / 107 = 0
    16'b00000000_01101100 : OUT <= 0;  //0 / 108 = 0
    16'b00000000_01101101 : OUT <= 0;  //0 / 109 = 0
    16'b00000000_01101110 : OUT <= 0;  //0 / 110 = 0
    16'b00000000_01101111 : OUT <= 0;  //0 / 111 = 0
    16'b00000000_01110000 : OUT <= 0;  //0 / 112 = 0
    16'b00000000_01110001 : OUT <= 0;  //0 / 113 = 0
    16'b00000000_01110010 : OUT <= 0;  //0 / 114 = 0
    16'b00000000_01110011 : OUT <= 0;  //0 / 115 = 0
    16'b00000000_01110100 : OUT <= 0;  //0 / 116 = 0
    16'b00000000_01110101 : OUT <= 0;  //0 / 117 = 0
    16'b00000000_01110110 : OUT <= 0;  //0 / 118 = 0
    16'b00000000_01110111 : OUT <= 0;  //0 / 119 = 0
    16'b00000000_01111000 : OUT <= 0;  //0 / 120 = 0
    16'b00000000_01111001 : OUT <= 0;  //0 / 121 = 0
    16'b00000000_01111010 : OUT <= 0;  //0 / 122 = 0
    16'b00000000_01111011 : OUT <= 0;  //0 / 123 = 0
    16'b00000000_01111100 : OUT <= 0;  //0 / 124 = 0
    16'b00000000_01111101 : OUT <= 0;  //0 / 125 = 0
    16'b00000000_01111110 : OUT <= 0;  //0 / 126 = 0
    16'b00000000_01111111 : OUT <= 0;  //0 / 127 = 0
    16'b00000000_10000000 : OUT <= 0;  //0 / 128 = 0
    16'b00000000_10000001 : OUT <= 0;  //0 / 129 = 0
    16'b00000000_10000010 : OUT <= 0;  //0 / 130 = 0
    16'b00000000_10000011 : OUT <= 0;  //0 / 131 = 0
    16'b00000000_10000100 : OUT <= 0;  //0 / 132 = 0
    16'b00000000_10000101 : OUT <= 0;  //0 / 133 = 0
    16'b00000000_10000110 : OUT <= 0;  //0 / 134 = 0
    16'b00000000_10000111 : OUT <= 0;  //0 / 135 = 0
    16'b00000000_10001000 : OUT <= 0;  //0 / 136 = 0
    16'b00000000_10001001 : OUT <= 0;  //0 / 137 = 0
    16'b00000000_10001010 : OUT <= 0;  //0 / 138 = 0
    16'b00000000_10001011 : OUT <= 0;  //0 / 139 = 0
    16'b00000000_10001100 : OUT <= 0;  //0 / 140 = 0
    16'b00000000_10001101 : OUT <= 0;  //0 / 141 = 0
    16'b00000000_10001110 : OUT <= 0;  //0 / 142 = 0
    16'b00000000_10001111 : OUT <= 0;  //0 / 143 = 0
    16'b00000000_10010000 : OUT <= 0;  //0 / 144 = 0
    16'b00000000_10010001 : OUT <= 0;  //0 / 145 = 0
    16'b00000000_10010010 : OUT <= 0;  //0 / 146 = 0
    16'b00000000_10010011 : OUT <= 0;  //0 / 147 = 0
    16'b00000000_10010100 : OUT <= 0;  //0 / 148 = 0
    16'b00000000_10010101 : OUT <= 0;  //0 / 149 = 0
    16'b00000000_10010110 : OUT <= 0;  //0 / 150 = 0
    16'b00000000_10010111 : OUT <= 0;  //0 / 151 = 0
    16'b00000000_10011000 : OUT <= 0;  //0 / 152 = 0
    16'b00000000_10011001 : OUT <= 0;  //0 / 153 = 0
    16'b00000000_10011010 : OUT <= 0;  //0 / 154 = 0
    16'b00000000_10011011 : OUT <= 0;  //0 / 155 = 0
    16'b00000000_10011100 : OUT <= 0;  //0 / 156 = 0
    16'b00000000_10011101 : OUT <= 0;  //0 / 157 = 0
    16'b00000000_10011110 : OUT <= 0;  //0 / 158 = 0
    16'b00000000_10011111 : OUT <= 0;  //0 / 159 = 0
    16'b00000000_10100000 : OUT <= 0;  //0 / 160 = 0
    16'b00000000_10100001 : OUT <= 0;  //0 / 161 = 0
    16'b00000000_10100010 : OUT <= 0;  //0 / 162 = 0
    16'b00000000_10100011 : OUT <= 0;  //0 / 163 = 0
    16'b00000000_10100100 : OUT <= 0;  //0 / 164 = 0
    16'b00000000_10100101 : OUT <= 0;  //0 / 165 = 0
    16'b00000000_10100110 : OUT <= 0;  //0 / 166 = 0
    16'b00000000_10100111 : OUT <= 0;  //0 / 167 = 0
    16'b00000000_10101000 : OUT <= 0;  //0 / 168 = 0
    16'b00000000_10101001 : OUT <= 0;  //0 / 169 = 0
    16'b00000000_10101010 : OUT <= 0;  //0 / 170 = 0
    16'b00000000_10101011 : OUT <= 0;  //0 / 171 = 0
    16'b00000000_10101100 : OUT <= 0;  //0 / 172 = 0
    16'b00000000_10101101 : OUT <= 0;  //0 / 173 = 0
    16'b00000000_10101110 : OUT <= 0;  //0 / 174 = 0
    16'b00000000_10101111 : OUT <= 0;  //0 / 175 = 0
    16'b00000000_10110000 : OUT <= 0;  //0 / 176 = 0
    16'b00000000_10110001 : OUT <= 0;  //0 / 177 = 0
    16'b00000000_10110010 : OUT <= 0;  //0 / 178 = 0
    16'b00000000_10110011 : OUT <= 0;  //0 / 179 = 0
    16'b00000000_10110100 : OUT <= 0;  //0 / 180 = 0
    16'b00000000_10110101 : OUT <= 0;  //0 / 181 = 0
    16'b00000000_10110110 : OUT <= 0;  //0 / 182 = 0
    16'b00000000_10110111 : OUT <= 0;  //0 / 183 = 0
    16'b00000000_10111000 : OUT <= 0;  //0 / 184 = 0
    16'b00000000_10111001 : OUT <= 0;  //0 / 185 = 0
    16'b00000000_10111010 : OUT <= 0;  //0 / 186 = 0
    16'b00000000_10111011 : OUT <= 0;  //0 / 187 = 0
    16'b00000000_10111100 : OUT <= 0;  //0 / 188 = 0
    16'b00000000_10111101 : OUT <= 0;  //0 / 189 = 0
    16'b00000000_10111110 : OUT <= 0;  //0 / 190 = 0
    16'b00000000_10111111 : OUT <= 0;  //0 / 191 = 0
    16'b00000000_11000000 : OUT <= 0;  //0 / 192 = 0
    16'b00000000_11000001 : OUT <= 0;  //0 / 193 = 0
    16'b00000000_11000010 : OUT <= 0;  //0 / 194 = 0
    16'b00000000_11000011 : OUT <= 0;  //0 / 195 = 0
    16'b00000000_11000100 : OUT <= 0;  //0 / 196 = 0
    16'b00000000_11000101 : OUT <= 0;  //0 / 197 = 0
    16'b00000000_11000110 : OUT <= 0;  //0 / 198 = 0
    16'b00000000_11000111 : OUT <= 0;  //0 / 199 = 0
    16'b00000000_11001000 : OUT <= 0;  //0 / 200 = 0
    16'b00000000_11001001 : OUT <= 0;  //0 / 201 = 0
    16'b00000000_11001010 : OUT <= 0;  //0 / 202 = 0
    16'b00000000_11001011 : OUT <= 0;  //0 / 203 = 0
    16'b00000000_11001100 : OUT <= 0;  //0 / 204 = 0
    16'b00000000_11001101 : OUT <= 0;  //0 / 205 = 0
    16'b00000000_11001110 : OUT <= 0;  //0 / 206 = 0
    16'b00000000_11001111 : OUT <= 0;  //0 / 207 = 0
    16'b00000000_11010000 : OUT <= 0;  //0 / 208 = 0
    16'b00000000_11010001 : OUT <= 0;  //0 / 209 = 0
    16'b00000000_11010010 : OUT <= 0;  //0 / 210 = 0
    16'b00000000_11010011 : OUT <= 0;  //0 / 211 = 0
    16'b00000000_11010100 : OUT <= 0;  //0 / 212 = 0
    16'b00000000_11010101 : OUT <= 0;  //0 / 213 = 0
    16'b00000000_11010110 : OUT <= 0;  //0 / 214 = 0
    16'b00000000_11010111 : OUT <= 0;  //0 / 215 = 0
    16'b00000000_11011000 : OUT <= 0;  //0 / 216 = 0
    16'b00000000_11011001 : OUT <= 0;  //0 / 217 = 0
    16'b00000000_11011010 : OUT <= 0;  //0 / 218 = 0
    16'b00000000_11011011 : OUT <= 0;  //0 / 219 = 0
    16'b00000000_11011100 : OUT <= 0;  //0 / 220 = 0
    16'b00000000_11011101 : OUT <= 0;  //0 / 221 = 0
    16'b00000000_11011110 : OUT <= 0;  //0 / 222 = 0
    16'b00000000_11011111 : OUT <= 0;  //0 / 223 = 0
    16'b00000000_11100000 : OUT <= 0;  //0 / 224 = 0
    16'b00000000_11100001 : OUT <= 0;  //0 / 225 = 0
    16'b00000000_11100010 : OUT <= 0;  //0 / 226 = 0
    16'b00000000_11100011 : OUT <= 0;  //0 / 227 = 0
    16'b00000000_11100100 : OUT <= 0;  //0 / 228 = 0
    16'b00000000_11100101 : OUT <= 0;  //0 / 229 = 0
    16'b00000000_11100110 : OUT <= 0;  //0 / 230 = 0
    16'b00000000_11100111 : OUT <= 0;  //0 / 231 = 0
    16'b00000000_11101000 : OUT <= 0;  //0 / 232 = 0
    16'b00000000_11101001 : OUT <= 0;  //0 / 233 = 0
    16'b00000000_11101010 : OUT <= 0;  //0 / 234 = 0
    16'b00000000_11101011 : OUT <= 0;  //0 / 235 = 0
    16'b00000000_11101100 : OUT <= 0;  //0 / 236 = 0
    16'b00000000_11101101 : OUT <= 0;  //0 / 237 = 0
    16'b00000000_11101110 : OUT <= 0;  //0 / 238 = 0
    16'b00000000_11101111 : OUT <= 0;  //0 / 239 = 0
    16'b00000000_11110000 : OUT <= 0;  //0 / 240 = 0
    16'b00000000_11110001 : OUT <= 0;  //0 / 241 = 0
    16'b00000000_11110010 : OUT <= 0;  //0 / 242 = 0
    16'b00000000_11110011 : OUT <= 0;  //0 / 243 = 0
    16'b00000000_11110100 : OUT <= 0;  //0 / 244 = 0
    16'b00000000_11110101 : OUT <= 0;  //0 / 245 = 0
    16'b00000000_11110110 : OUT <= 0;  //0 / 246 = 0
    16'b00000000_11110111 : OUT <= 0;  //0 / 247 = 0
    16'b00000000_11111000 : OUT <= 0;  //0 / 248 = 0
    16'b00000000_11111001 : OUT <= 0;  //0 / 249 = 0
    16'b00000000_11111010 : OUT <= 0;  //0 / 250 = 0
    16'b00000000_11111011 : OUT <= 0;  //0 / 251 = 0
    16'b00000000_11111100 : OUT <= 0;  //0 / 252 = 0
    16'b00000000_11111101 : OUT <= 0;  //0 / 253 = 0
    16'b00000000_11111110 : OUT <= 0;  //0 / 254 = 0
    16'b00000000_11111111 : OUT <= 0;  //0 / 255 = 0
    16'b00000001_00000000 : OUT <= 0;  //1 / 0 = 0
    16'b00000001_00000001 : OUT <= 1;  //1 / 1 = 1
    16'b00000001_00000010 : OUT <= 0;  //1 / 2 = 0
    16'b00000001_00000011 : OUT <= 0;  //1 / 3 = 0
    16'b00000001_00000100 : OUT <= 0;  //1 / 4 = 0
    16'b00000001_00000101 : OUT <= 0;  //1 / 5 = 0
    16'b00000001_00000110 : OUT <= 0;  //1 / 6 = 0
    16'b00000001_00000111 : OUT <= 0;  //1 / 7 = 0
    16'b00000001_00001000 : OUT <= 0;  //1 / 8 = 0
    16'b00000001_00001001 : OUT <= 0;  //1 / 9 = 0
    16'b00000001_00001010 : OUT <= 0;  //1 / 10 = 0
    16'b00000001_00001011 : OUT <= 0;  //1 / 11 = 0
    16'b00000001_00001100 : OUT <= 0;  //1 / 12 = 0
    16'b00000001_00001101 : OUT <= 0;  //1 / 13 = 0
    16'b00000001_00001110 : OUT <= 0;  //1 / 14 = 0
    16'b00000001_00001111 : OUT <= 0;  //1 / 15 = 0
    16'b00000001_00010000 : OUT <= 0;  //1 / 16 = 0
    16'b00000001_00010001 : OUT <= 0;  //1 / 17 = 0
    16'b00000001_00010010 : OUT <= 0;  //1 / 18 = 0
    16'b00000001_00010011 : OUT <= 0;  //1 / 19 = 0
    16'b00000001_00010100 : OUT <= 0;  //1 / 20 = 0
    16'b00000001_00010101 : OUT <= 0;  //1 / 21 = 0
    16'b00000001_00010110 : OUT <= 0;  //1 / 22 = 0
    16'b00000001_00010111 : OUT <= 0;  //1 / 23 = 0
    16'b00000001_00011000 : OUT <= 0;  //1 / 24 = 0
    16'b00000001_00011001 : OUT <= 0;  //1 / 25 = 0
    16'b00000001_00011010 : OUT <= 0;  //1 / 26 = 0
    16'b00000001_00011011 : OUT <= 0;  //1 / 27 = 0
    16'b00000001_00011100 : OUT <= 0;  //1 / 28 = 0
    16'b00000001_00011101 : OUT <= 0;  //1 / 29 = 0
    16'b00000001_00011110 : OUT <= 0;  //1 / 30 = 0
    16'b00000001_00011111 : OUT <= 0;  //1 / 31 = 0
    16'b00000001_00100000 : OUT <= 0;  //1 / 32 = 0
    16'b00000001_00100001 : OUT <= 0;  //1 / 33 = 0
    16'b00000001_00100010 : OUT <= 0;  //1 / 34 = 0
    16'b00000001_00100011 : OUT <= 0;  //1 / 35 = 0
    16'b00000001_00100100 : OUT <= 0;  //1 / 36 = 0
    16'b00000001_00100101 : OUT <= 0;  //1 / 37 = 0
    16'b00000001_00100110 : OUT <= 0;  //1 / 38 = 0
    16'b00000001_00100111 : OUT <= 0;  //1 / 39 = 0
    16'b00000001_00101000 : OUT <= 0;  //1 / 40 = 0
    16'b00000001_00101001 : OUT <= 0;  //1 / 41 = 0
    16'b00000001_00101010 : OUT <= 0;  //1 / 42 = 0
    16'b00000001_00101011 : OUT <= 0;  //1 / 43 = 0
    16'b00000001_00101100 : OUT <= 0;  //1 / 44 = 0
    16'b00000001_00101101 : OUT <= 0;  //1 / 45 = 0
    16'b00000001_00101110 : OUT <= 0;  //1 / 46 = 0
    16'b00000001_00101111 : OUT <= 0;  //1 / 47 = 0
    16'b00000001_00110000 : OUT <= 0;  //1 / 48 = 0
    16'b00000001_00110001 : OUT <= 0;  //1 / 49 = 0
    16'b00000001_00110010 : OUT <= 0;  //1 / 50 = 0
    16'b00000001_00110011 : OUT <= 0;  //1 / 51 = 0
    16'b00000001_00110100 : OUT <= 0;  //1 / 52 = 0
    16'b00000001_00110101 : OUT <= 0;  //1 / 53 = 0
    16'b00000001_00110110 : OUT <= 0;  //1 / 54 = 0
    16'b00000001_00110111 : OUT <= 0;  //1 / 55 = 0
    16'b00000001_00111000 : OUT <= 0;  //1 / 56 = 0
    16'b00000001_00111001 : OUT <= 0;  //1 / 57 = 0
    16'b00000001_00111010 : OUT <= 0;  //1 / 58 = 0
    16'b00000001_00111011 : OUT <= 0;  //1 / 59 = 0
    16'b00000001_00111100 : OUT <= 0;  //1 / 60 = 0
    16'b00000001_00111101 : OUT <= 0;  //1 / 61 = 0
    16'b00000001_00111110 : OUT <= 0;  //1 / 62 = 0
    16'b00000001_00111111 : OUT <= 0;  //1 / 63 = 0
    16'b00000001_01000000 : OUT <= 0;  //1 / 64 = 0
    16'b00000001_01000001 : OUT <= 0;  //1 / 65 = 0
    16'b00000001_01000010 : OUT <= 0;  //1 / 66 = 0
    16'b00000001_01000011 : OUT <= 0;  //1 / 67 = 0
    16'b00000001_01000100 : OUT <= 0;  //1 / 68 = 0
    16'b00000001_01000101 : OUT <= 0;  //1 / 69 = 0
    16'b00000001_01000110 : OUT <= 0;  //1 / 70 = 0
    16'b00000001_01000111 : OUT <= 0;  //1 / 71 = 0
    16'b00000001_01001000 : OUT <= 0;  //1 / 72 = 0
    16'b00000001_01001001 : OUT <= 0;  //1 / 73 = 0
    16'b00000001_01001010 : OUT <= 0;  //1 / 74 = 0
    16'b00000001_01001011 : OUT <= 0;  //1 / 75 = 0
    16'b00000001_01001100 : OUT <= 0;  //1 / 76 = 0
    16'b00000001_01001101 : OUT <= 0;  //1 / 77 = 0
    16'b00000001_01001110 : OUT <= 0;  //1 / 78 = 0
    16'b00000001_01001111 : OUT <= 0;  //1 / 79 = 0
    16'b00000001_01010000 : OUT <= 0;  //1 / 80 = 0
    16'b00000001_01010001 : OUT <= 0;  //1 / 81 = 0
    16'b00000001_01010010 : OUT <= 0;  //1 / 82 = 0
    16'b00000001_01010011 : OUT <= 0;  //1 / 83 = 0
    16'b00000001_01010100 : OUT <= 0;  //1 / 84 = 0
    16'b00000001_01010101 : OUT <= 0;  //1 / 85 = 0
    16'b00000001_01010110 : OUT <= 0;  //1 / 86 = 0
    16'b00000001_01010111 : OUT <= 0;  //1 / 87 = 0
    16'b00000001_01011000 : OUT <= 0;  //1 / 88 = 0
    16'b00000001_01011001 : OUT <= 0;  //1 / 89 = 0
    16'b00000001_01011010 : OUT <= 0;  //1 / 90 = 0
    16'b00000001_01011011 : OUT <= 0;  //1 / 91 = 0
    16'b00000001_01011100 : OUT <= 0;  //1 / 92 = 0
    16'b00000001_01011101 : OUT <= 0;  //1 / 93 = 0
    16'b00000001_01011110 : OUT <= 0;  //1 / 94 = 0
    16'b00000001_01011111 : OUT <= 0;  //1 / 95 = 0
    16'b00000001_01100000 : OUT <= 0;  //1 / 96 = 0
    16'b00000001_01100001 : OUT <= 0;  //1 / 97 = 0
    16'b00000001_01100010 : OUT <= 0;  //1 / 98 = 0
    16'b00000001_01100011 : OUT <= 0;  //1 / 99 = 0
    16'b00000001_01100100 : OUT <= 0;  //1 / 100 = 0
    16'b00000001_01100101 : OUT <= 0;  //1 / 101 = 0
    16'b00000001_01100110 : OUT <= 0;  //1 / 102 = 0
    16'b00000001_01100111 : OUT <= 0;  //1 / 103 = 0
    16'b00000001_01101000 : OUT <= 0;  //1 / 104 = 0
    16'b00000001_01101001 : OUT <= 0;  //1 / 105 = 0
    16'b00000001_01101010 : OUT <= 0;  //1 / 106 = 0
    16'b00000001_01101011 : OUT <= 0;  //1 / 107 = 0
    16'b00000001_01101100 : OUT <= 0;  //1 / 108 = 0
    16'b00000001_01101101 : OUT <= 0;  //1 / 109 = 0
    16'b00000001_01101110 : OUT <= 0;  //1 / 110 = 0
    16'b00000001_01101111 : OUT <= 0;  //1 / 111 = 0
    16'b00000001_01110000 : OUT <= 0;  //1 / 112 = 0
    16'b00000001_01110001 : OUT <= 0;  //1 / 113 = 0
    16'b00000001_01110010 : OUT <= 0;  //1 / 114 = 0
    16'b00000001_01110011 : OUT <= 0;  //1 / 115 = 0
    16'b00000001_01110100 : OUT <= 0;  //1 / 116 = 0
    16'b00000001_01110101 : OUT <= 0;  //1 / 117 = 0
    16'b00000001_01110110 : OUT <= 0;  //1 / 118 = 0
    16'b00000001_01110111 : OUT <= 0;  //1 / 119 = 0
    16'b00000001_01111000 : OUT <= 0;  //1 / 120 = 0
    16'b00000001_01111001 : OUT <= 0;  //1 / 121 = 0
    16'b00000001_01111010 : OUT <= 0;  //1 / 122 = 0
    16'b00000001_01111011 : OUT <= 0;  //1 / 123 = 0
    16'b00000001_01111100 : OUT <= 0;  //1 / 124 = 0
    16'b00000001_01111101 : OUT <= 0;  //1 / 125 = 0
    16'b00000001_01111110 : OUT <= 0;  //1 / 126 = 0
    16'b00000001_01111111 : OUT <= 0;  //1 / 127 = 0
    16'b00000001_10000000 : OUT <= 0;  //1 / 128 = 0
    16'b00000001_10000001 : OUT <= 0;  //1 / 129 = 0
    16'b00000001_10000010 : OUT <= 0;  //1 / 130 = 0
    16'b00000001_10000011 : OUT <= 0;  //1 / 131 = 0
    16'b00000001_10000100 : OUT <= 0;  //1 / 132 = 0
    16'b00000001_10000101 : OUT <= 0;  //1 / 133 = 0
    16'b00000001_10000110 : OUT <= 0;  //1 / 134 = 0
    16'b00000001_10000111 : OUT <= 0;  //1 / 135 = 0
    16'b00000001_10001000 : OUT <= 0;  //1 / 136 = 0
    16'b00000001_10001001 : OUT <= 0;  //1 / 137 = 0
    16'b00000001_10001010 : OUT <= 0;  //1 / 138 = 0
    16'b00000001_10001011 : OUT <= 0;  //1 / 139 = 0
    16'b00000001_10001100 : OUT <= 0;  //1 / 140 = 0
    16'b00000001_10001101 : OUT <= 0;  //1 / 141 = 0
    16'b00000001_10001110 : OUT <= 0;  //1 / 142 = 0
    16'b00000001_10001111 : OUT <= 0;  //1 / 143 = 0
    16'b00000001_10010000 : OUT <= 0;  //1 / 144 = 0
    16'b00000001_10010001 : OUT <= 0;  //1 / 145 = 0
    16'b00000001_10010010 : OUT <= 0;  //1 / 146 = 0
    16'b00000001_10010011 : OUT <= 0;  //1 / 147 = 0
    16'b00000001_10010100 : OUT <= 0;  //1 / 148 = 0
    16'b00000001_10010101 : OUT <= 0;  //1 / 149 = 0
    16'b00000001_10010110 : OUT <= 0;  //1 / 150 = 0
    16'b00000001_10010111 : OUT <= 0;  //1 / 151 = 0
    16'b00000001_10011000 : OUT <= 0;  //1 / 152 = 0
    16'b00000001_10011001 : OUT <= 0;  //1 / 153 = 0
    16'b00000001_10011010 : OUT <= 0;  //1 / 154 = 0
    16'b00000001_10011011 : OUT <= 0;  //1 / 155 = 0
    16'b00000001_10011100 : OUT <= 0;  //1 / 156 = 0
    16'b00000001_10011101 : OUT <= 0;  //1 / 157 = 0
    16'b00000001_10011110 : OUT <= 0;  //1 / 158 = 0
    16'b00000001_10011111 : OUT <= 0;  //1 / 159 = 0
    16'b00000001_10100000 : OUT <= 0;  //1 / 160 = 0
    16'b00000001_10100001 : OUT <= 0;  //1 / 161 = 0
    16'b00000001_10100010 : OUT <= 0;  //1 / 162 = 0
    16'b00000001_10100011 : OUT <= 0;  //1 / 163 = 0
    16'b00000001_10100100 : OUT <= 0;  //1 / 164 = 0
    16'b00000001_10100101 : OUT <= 0;  //1 / 165 = 0
    16'b00000001_10100110 : OUT <= 0;  //1 / 166 = 0
    16'b00000001_10100111 : OUT <= 0;  //1 / 167 = 0
    16'b00000001_10101000 : OUT <= 0;  //1 / 168 = 0
    16'b00000001_10101001 : OUT <= 0;  //1 / 169 = 0
    16'b00000001_10101010 : OUT <= 0;  //1 / 170 = 0
    16'b00000001_10101011 : OUT <= 0;  //1 / 171 = 0
    16'b00000001_10101100 : OUT <= 0;  //1 / 172 = 0
    16'b00000001_10101101 : OUT <= 0;  //1 / 173 = 0
    16'b00000001_10101110 : OUT <= 0;  //1 / 174 = 0
    16'b00000001_10101111 : OUT <= 0;  //1 / 175 = 0
    16'b00000001_10110000 : OUT <= 0;  //1 / 176 = 0
    16'b00000001_10110001 : OUT <= 0;  //1 / 177 = 0
    16'b00000001_10110010 : OUT <= 0;  //1 / 178 = 0
    16'b00000001_10110011 : OUT <= 0;  //1 / 179 = 0
    16'b00000001_10110100 : OUT <= 0;  //1 / 180 = 0
    16'b00000001_10110101 : OUT <= 0;  //1 / 181 = 0
    16'b00000001_10110110 : OUT <= 0;  //1 / 182 = 0
    16'b00000001_10110111 : OUT <= 0;  //1 / 183 = 0
    16'b00000001_10111000 : OUT <= 0;  //1 / 184 = 0
    16'b00000001_10111001 : OUT <= 0;  //1 / 185 = 0
    16'b00000001_10111010 : OUT <= 0;  //1 / 186 = 0
    16'b00000001_10111011 : OUT <= 0;  //1 / 187 = 0
    16'b00000001_10111100 : OUT <= 0;  //1 / 188 = 0
    16'b00000001_10111101 : OUT <= 0;  //1 / 189 = 0
    16'b00000001_10111110 : OUT <= 0;  //1 / 190 = 0
    16'b00000001_10111111 : OUT <= 0;  //1 / 191 = 0
    16'b00000001_11000000 : OUT <= 0;  //1 / 192 = 0
    16'b00000001_11000001 : OUT <= 0;  //1 / 193 = 0
    16'b00000001_11000010 : OUT <= 0;  //1 / 194 = 0
    16'b00000001_11000011 : OUT <= 0;  //1 / 195 = 0
    16'b00000001_11000100 : OUT <= 0;  //1 / 196 = 0
    16'b00000001_11000101 : OUT <= 0;  //1 / 197 = 0
    16'b00000001_11000110 : OUT <= 0;  //1 / 198 = 0
    16'b00000001_11000111 : OUT <= 0;  //1 / 199 = 0
    16'b00000001_11001000 : OUT <= 0;  //1 / 200 = 0
    16'b00000001_11001001 : OUT <= 0;  //1 / 201 = 0
    16'b00000001_11001010 : OUT <= 0;  //1 / 202 = 0
    16'b00000001_11001011 : OUT <= 0;  //1 / 203 = 0
    16'b00000001_11001100 : OUT <= 0;  //1 / 204 = 0
    16'b00000001_11001101 : OUT <= 0;  //1 / 205 = 0
    16'b00000001_11001110 : OUT <= 0;  //1 / 206 = 0
    16'b00000001_11001111 : OUT <= 0;  //1 / 207 = 0
    16'b00000001_11010000 : OUT <= 0;  //1 / 208 = 0
    16'b00000001_11010001 : OUT <= 0;  //1 / 209 = 0
    16'b00000001_11010010 : OUT <= 0;  //1 / 210 = 0
    16'b00000001_11010011 : OUT <= 0;  //1 / 211 = 0
    16'b00000001_11010100 : OUT <= 0;  //1 / 212 = 0
    16'b00000001_11010101 : OUT <= 0;  //1 / 213 = 0
    16'b00000001_11010110 : OUT <= 0;  //1 / 214 = 0
    16'b00000001_11010111 : OUT <= 0;  //1 / 215 = 0
    16'b00000001_11011000 : OUT <= 0;  //1 / 216 = 0
    16'b00000001_11011001 : OUT <= 0;  //1 / 217 = 0
    16'b00000001_11011010 : OUT <= 0;  //1 / 218 = 0
    16'b00000001_11011011 : OUT <= 0;  //1 / 219 = 0
    16'b00000001_11011100 : OUT <= 0;  //1 / 220 = 0
    16'b00000001_11011101 : OUT <= 0;  //1 / 221 = 0
    16'b00000001_11011110 : OUT <= 0;  //1 / 222 = 0
    16'b00000001_11011111 : OUT <= 0;  //1 / 223 = 0
    16'b00000001_11100000 : OUT <= 0;  //1 / 224 = 0
    16'b00000001_11100001 : OUT <= 0;  //1 / 225 = 0
    16'b00000001_11100010 : OUT <= 0;  //1 / 226 = 0
    16'b00000001_11100011 : OUT <= 0;  //1 / 227 = 0
    16'b00000001_11100100 : OUT <= 0;  //1 / 228 = 0
    16'b00000001_11100101 : OUT <= 0;  //1 / 229 = 0
    16'b00000001_11100110 : OUT <= 0;  //1 / 230 = 0
    16'b00000001_11100111 : OUT <= 0;  //1 / 231 = 0
    16'b00000001_11101000 : OUT <= 0;  //1 / 232 = 0
    16'b00000001_11101001 : OUT <= 0;  //1 / 233 = 0
    16'b00000001_11101010 : OUT <= 0;  //1 / 234 = 0
    16'b00000001_11101011 : OUT <= 0;  //1 / 235 = 0
    16'b00000001_11101100 : OUT <= 0;  //1 / 236 = 0
    16'b00000001_11101101 : OUT <= 0;  //1 / 237 = 0
    16'b00000001_11101110 : OUT <= 0;  //1 / 238 = 0
    16'b00000001_11101111 : OUT <= 0;  //1 / 239 = 0
    16'b00000001_11110000 : OUT <= 0;  //1 / 240 = 0
    16'b00000001_11110001 : OUT <= 0;  //1 / 241 = 0
    16'b00000001_11110010 : OUT <= 0;  //1 / 242 = 0
    16'b00000001_11110011 : OUT <= 0;  //1 / 243 = 0
    16'b00000001_11110100 : OUT <= 0;  //1 / 244 = 0
    16'b00000001_11110101 : OUT <= 0;  //1 / 245 = 0
    16'b00000001_11110110 : OUT <= 0;  //1 / 246 = 0
    16'b00000001_11110111 : OUT <= 0;  //1 / 247 = 0
    16'b00000001_11111000 : OUT <= 0;  //1 / 248 = 0
    16'b00000001_11111001 : OUT <= 0;  //1 / 249 = 0
    16'b00000001_11111010 : OUT <= 0;  //1 / 250 = 0
    16'b00000001_11111011 : OUT <= 0;  //1 / 251 = 0
    16'b00000001_11111100 : OUT <= 0;  //1 / 252 = 0
    16'b00000001_11111101 : OUT <= 0;  //1 / 253 = 0
    16'b00000001_11111110 : OUT <= 0;  //1 / 254 = 0
    16'b00000001_11111111 : OUT <= 0;  //1 / 255 = 0
    16'b00000010_00000000 : OUT <= 0;  //2 / 0 = 0
    16'b00000010_00000001 : OUT <= 2;  //2 / 1 = 2
    16'b00000010_00000010 : OUT <= 1;  //2 / 2 = 1
    16'b00000010_00000011 : OUT <= 0;  //2 / 3 = 0
    16'b00000010_00000100 : OUT <= 0;  //2 / 4 = 0
    16'b00000010_00000101 : OUT <= 0;  //2 / 5 = 0
    16'b00000010_00000110 : OUT <= 0;  //2 / 6 = 0
    16'b00000010_00000111 : OUT <= 0;  //2 / 7 = 0
    16'b00000010_00001000 : OUT <= 0;  //2 / 8 = 0
    16'b00000010_00001001 : OUT <= 0;  //2 / 9 = 0
    16'b00000010_00001010 : OUT <= 0;  //2 / 10 = 0
    16'b00000010_00001011 : OUT <= 0;  //2 / 11 = 0
    16'b00000010_00001100 : OUT <= 0;  //2 / 12 = 0
    16'b00000010_00001101 : OUT <= 0;  //2 / 13 = 0
    16'b00000010_00001110 : OUT <= 0;  //2 / 14 = 0
    16'b00000010_00001111 : OUT <= 0;  //2 / 15 = 0
    16'b00000010_00010000 : OUT <= 0;  //2 / 16 = 0
    16'b00000010_00010001 : OUT <= 0;  //2 / 17 = 0
    16'b00000010_00010010 : OUT <= 0;  //2 / 18 = 0
    16'b00000010_00010011 : OUT <= 0;  //2 / 19 = 0
    16'b00000010_00010100 : OUT <= 0;  //2 / 20 = 0
    16'b00000010_00010101 : OUT <= 0;  //2 / 21 = 0
    16'b00000010_00010110 : OUT <= 0;  //2 / 22 = 0
    16'b00000010_00010111 : OUT <= 0;  //2 / 23 = 0
    16'b00000010_00011000 : OUT <= 0;  //2 / 24 = 0
    16'b00000010_00011001 : OUT <= 0;  //2 / 25 = 0
    16'b00000010_00011010 : OUT <= 0;  //2 / 26 = 0
    16'b00000010_00011011 : OUT <= 0;  //2 / 27 = 0
    16'b00000010_00011100 : OUT <= 0;  //2 / 28 = 0
    16'b00000010_00011101 : OUT <= 0;  //2 / 29 = 0
    16'b00000010_00011110 : OUT <= 0;  //2 / 30 = 0
    16'b00000010_00011111 : OUT <= 0;  //2 / 31 = 0
    16'b00000010_00100000 : OUT <= 0;  //2 / 32 = 0
    16'b00000010_00100001 : OUT <= 0;  //2 / 33 = 0
    16'b00000010_00100010 : OUT <= 0;  //2 / 34 = 0
    16'b00000010_00100011 : OUT <= 0;  //2 / 35 = 0
    16'b00000010_00100100 : OUT <= 0;  //2 / 36 = 0
    16'b00000010_00100101 : OUT <= 0;  //2 / 37 = 0
    16'b00000010_00100110 : OUT <= 0;  //2 / 38 = 0
    16'b00000010_00100111 : OUT <= 0;  //2 / 39 = 0
    16'b00000010_00101000 : OUT <= 0;  //2 / 40 = 0
    16'b00000010_00101001 : OUT <= 0;  //2 / 41 = 0
    16'b00000010_00101010 : OUT <= 0;  //2 / 42 = 0
    16'b00000010_00101011 : OUT <= 0;  //2 / 43 = 0
    16'b00000010_00101100 : OUT <= 0;  //2 / 44 = 0
    16'b00000010_00101101 : OUT <= 0;  //2 / 45 = 0
    16'b00000010_00101110 : OUT <= 0;  //2 / 46 = 0
    16'b00000010_00101111 : OUT <= 0;  //2 / 47 = 0
    16'b00000010_00110000 : OUT <= 0;  //2 / 48 = 0
    16'b00000010_00110001 : OUT <= 0;  //2 / 49 = 0
    16'b00000010_00110010 : OUT <= 0;  //2 / 50 = 0
    16'b00000010_00110011 : OUT <= 0;  //2 / 51 = 0
    16'b00000010_00110100 : OUT <= 0;  //2 / 52 = 0
    16'b00000010_00110101 : OUT <= 0;  //2 / 53 = 0
    16'b00000010_00110110 : OUT <= 0;  //2 / 54 = 0
    16'b00000010_00110111 : OUT <= 0;  //2 / 55 = 0
    16'b00000010_00111000 : OUT <= 0;  //2 / 56 = 0
    16'b00000010_00111001 : OUT <= 0;  //2 / 57 = 0
    16'b00000010_00111010 : OUT <= 0;  //2 / 58 = 0
    16'b00000010_00111011 : OUT <= 0;  //2 / 59 = 0
    16'b00000010_00111100 : OUT <= 0;  //2 / 60 = 0
    16'b00000010_00111101 : OUT <= 0;  //2 / 61 = 0
    16'b00000010_00111110 : OUT <= 0;  //2 / 62 = 0
    16'b00000010_00111111 : OUT <= 0;  //2 / 63 = 0
    16'b00000010_01000000 : OUT <= 0;  //2 / 64 = 0
    16'b00000010_01000001 : OUT <= 0;  //2 / 65 = 0
    16'b00000010_01000010 : OUT <= 0;  //2 / 66 = 0
    16'b00000010_01000011 : OUT <= 0;  //2 / 67 = 0
    16'b00000010_01000100 : OUT <= 0;  //2 / 68 = 0
    16'b00000010_01000101 : OUT <= 0;  //2 / 69 = 0
    16'b00000010_01000110 : OUT <= 0;  //2 / 70 = 0
    16'b00000010_01000111 : OUT <= 0;  //2 / 71 = 0
    16'b00000010_01001000 : OUT <= 0;  //2 / 72 = 0
    16'b00000010_01001001 : OUT <= 0;  //2 / 73 = 0
    16'b00000010_01001010 : OUT <= 0;  //2 / 74 = 0
    16'b00000010_01001011 : OUT <= 0;  //2 / 75 = 0
    16'b00000010_01001100 : OUT <= 0;  //2 / 76 = 0
    16'b00000010_01001101 : OUT <= 0;  //2 / 77 = 0
    16'b00000010_01001110 : OUT <= 0;  //2 / 78 = 0
    16'b00000010_01001111 : OUT <= 0;  //2 / 79 = 0
    16'b00000010_01010000 : OUT <= 0;  //2 / 80 = 0
    16'b00000010_01010001 : OUT <= 0;  //2 / 81 = 0
    16'b00000010_01010010 : OUT <= 0;  //2 / 82 = 0
    16'b00000010_01010011 : OUT <= 0;  //2 / 83 = 0
    16'b00000010_01010100 : OUT <= 0;  //2 / 84 = 0
    16'b00000010_01010101 : OUT <= 0;  //2 / 85 = 0
    16'b00000010_01010110 : OUT <= 0;  //2 / 86 = 0
    16'b00000010_01010111 : OUT <= 0;  //2 / 87 = 0
    16'b00000010_01011000 : OUT <= 0;  //2 / 88 = 0
    16'b00000010_01011001 : OUT <= 0;  //2 / 89 = 0
    16'b00000010_01011010 : OUT <= 0;  //2 / 90 = 0
    16'b00000010_01011011 : OUT <= 0;  //2 / 91 = 0
    16'b00000010_01011100 : OUT <= 0;  //2 / 92 = 0
    16'b00000010_01011101 : OUT <= 0;  //2 / 93 = 0
    16'b00000010_01011110 : OUT <= 0;  //2 / 94 = 0
    16'b00000010_01011111 : OUT <= 0;  //2 / 95 = 0
    16'b00000010_01100000 : OUT <= 0;  //2 / 96 = 0
    16'b00000010_01100001 : OUT <= 0;  //2 / 97 = 0
    16'b00000010_01100010 : OUT <= 0;  //2 / 98 = 0
    16'b00000010_01100011 : OUT <= 0;  //2 / 99 = 0
    16'b00000010_01100100 : OUT <= 0;  //2 / 100 = 0
    16'b00000010_01100101 : OUT <= 0;  //2 / 101 = 0
    16'b00000010_01100110 : OUT <= 0;  //2 / 102 = 0
    16'b00000010_01100111 : OUT <= 0;  //2 / 103 = 0
    16'b00000010_01101000 : OUT <= 0;  //2 / 104 = 0
    16'b00000010_01101001 : OUT <= 0;  //2 / 105 = 0
    16'b00000010_01101010 : OUT <= 0;  //2 / 106 = 0
    16'b00000010_01101011 : OUT <= 0;  //2 / 107 = 0
    16'b00000010_01101100 : OUT <= 0;  //2 / 108 = 0
    16'b00000010_01101101 : OUT <= 0;  //2 / 109 = 0
    16'b00000010_01101110 : OUT <= 0;  //2 / 110 = 0
    16'b00000010_01101111 : OUT <= 0;  //2 / 111 = 0
    16'b00000010_01110000 : OUT <= 0;  //2 / 112 = 0
    16'b00000010_01110001 : OUT <= 0;  //2 / 113 = 0
    16'b00000010_01110010 : OUT <= 0;  //2 / 114 = 0
    16'b00000010_01110011 : OUT <= 0;  //2 / 115 = 0
    16'b00000010_01110100 : OUT <= 0;  //2 / 116 = 0
    16'b00000010_01110101 : OUT <= 0;  //2 / 117 = 0
    16'b00000010_01110110 : OUT <= 0;  //2 / 118 = 0
    16'b00000010_01110111 : OUT <= 0;  //2 / 119 = 0
    16'b00000010_01111000 : OUT <= 0;  //2 / 120 = 0
    16'b00000010_01111001 : OUT <= 0;  //2 / 121 = 0
    16'b00000010_01111010 : OUT <= 0;  //2 / 122 = 0
    16'b00000010_01111011 : OUT <= 0;  //2 / 123 = 0
    16'b00000010_01111100 : OUT <= 0;  //2 / 124 = 0
    16'b00000010_01111101 : OUT <= 0;  //2 / 125 = 0
    16'b00000010_01111110 : OUT <= 0;  //2 / 126 = 0
    16'b00000010_01111111 : OUT <= 0;  //2 / 127 = 0
    16'b00000010_10000000 : OUT <= 0;  //2 / 128 = 0
    16'b00000010_10000001 : OUT <= 0;  //2 / 129 = 0
    16'b00000010_10000010 : OUT <= 0;  //2 / 130 = 0
    16'b00000010_10000011 : OUT <= 0;  //2 / 131 = 0
    16'b00000010_10000100 : OUT <= 0;  //2 / 132 = 0
    16'b00000010_10000101 : OUT <= 0;  //2 / 133 = 0
    16'b00000010_10000110 : OUT <= 0;  //2 / 134 = 0
    16'b00000010_10000111 : OUT <= 0;  //2 / 135 = 0
    16'b00000010_10001000 : OUT <= 0;  //2 / 136 = 0
    16'b00000010_10001001 : OUT <= 0;  //2 / 137 = 0
    16'b00000010_10001010 : OUT <= 0;  //2 / 138 = 0
    16'b00000010_10001011 : OUT <= 0;  //2 / 139 = 0
    16'b00000010_10001100 : OUT <= 0;  //2 / 140 = 0
    16'b00000010_10001101 : OUT <= 0;  //2 / 141 = 0
    16'b00000010_10001110 : OUT <= 0;  //2 / 142 = 0
    16'b00000010_10001111 : OUT <= 0;  //2 / 143 = 0
    16'b00000010_10010000 : OUT <= 0;  //2 / 144 = 0
    16'b00000010_10010001 : OUT <= 0;  //2 / 145 = 0
    16'b00000010_10010010 : OUT <= 0;  //2 / 146 = 0
    16'b00000010_10010011 : OUT <= 0;  //2 / 147 = 0
    16'b00000010_10010100 : OUT <= 0;  //2 / 148 = 0
    16'b00000010_10010101 : OUT <= 0;  //2 / 149 = 0
    16'b00000010_10010110 : OUT <= 0;  //2 / 150 = 0
    16'b00000010_10010111 : OUT <= 0;  //2 / 151 = 0
    16'b00000010_10011000 : OUT <= 0;  //2 / 152 = 0
    16'b00000010_10011001 : OUT <= 0;  //2 / 153 = 0
    16'b00000010_10011010 : OUT <= 0;  //2 / 154 = 0
    16'b00000010_10011011 : OUT <= 0;  //2 / 155 = 0
    16'b00000010_10011100 : OUT <= 0;  //2 / 156 = 0
    16'b00000010_10011101 : OUT <= 0;  //2 / 157 = 0
    16'b00000010_10011110 : OUT <= 0;  //2 / 158 = 0
    16'b00000010_10011111 : OUT <= 0;  //2 / 159 = 0
    16'b00000010_10100000 : OUT <= 0;  //2 / 160 = 0
    16'b00000010_10100001 : OUT <= 0;  //2 / 161 = 0
    16'b00000010_10100010 : OUT <= 0;  //2 / 162 = 0
    16'b00000010_10100011 : OUT <= 0;  //2 / 163 = 0
    16'b00000010_10100100 : OUT <= 0;  //2 / 164 = 0
    16'b00000010_10100101 : OUT <= 0;  //2 / 165 = 0
    16'b00000010_10100110 : OUT <= 0;  //2 / 166 = 0
    16'b00000010_10100111 : OUT <= 0;  //2 / 167 = 0
    16'b00000010_10101000 : OUT <= 0;  //2 / 168 = 0
    16'b00000010_10101001 : OUT <= 0;  //2 / 169 = 0
    16'b00000010_10101010 : OUT <= 0;  //2 / 170 = 0
    16'b00000010_10101011 : OUT <= 0;  //2 / 171 = 0
    16'b00000010_10101100 : OUT <= 0;  //2 / 172 = 0
    16'b00000010_10101101 : OUT <= 0;  //2 / 173 = 0
    16'b00000010_10101110 : OUT <= 0;  //2 / 174 = 0
    16'b00000010_10101111 : OUT <= 0;  //2 / 175 = 0
    16'b00000010_10110000 : OUT <= 0;  //2 / 176 = 0
    16'b00000010_10110001 : OUT <= 0;  //2 / 177 = 0
    16'b00000010_10110010 : OUT <= 0;  //2 / 178 = 0
    16'b00000010_10110011 : OUT <= 0;  //2 / 179 = 0
    16'b00000010_10110100 : OUT <= 0;  //2 / 180 = 0
    16'b00000010_10110101 : OUT <= 0;  //2 / 181 = 0
    16'b00000010_10110110 : OUT <= 0;  //2 / 182 = 0
    16'b00000010_10110111 : OUT <= 0;  //2 / 183 = 0
    16'b00000010_10111000 : OUT <= 0;  //2 / 184 = 0
    16'b00000010_10111001 : OUT <= 0;  //2 / 185 = 0
    16'b00000010_10111010 : OUT <= 0;  //2 / 186 = 0
    16'b00000010_10111011 : OUT <= 0;  //2 / 187 = 0
    16'b00000010_10111100 : OUT <= 0;  //2 / 188 = 0
    16'b00000010_10111101 : OUT <= 0;  //2 / 189 = 0
    16'b00000010_10111110 : OUT <= 0;  //2 / 190 = 0
    16'b00000010_10111111 : OUT <= 0;  //2 / 191 = 0
    16'b00000010_11000000 : OUT <= 0;  //2 / 192 = 0
    16'b00000010_11000001 : OUT <= 0;  //2 / 193 = 0
    16'b00000010_11000010 : OUT <= 0;  //2 / 194 = 0
    16'b00000010_11000011 : OUT <= 0;  //2 / 195 = 0
    16'b00000010_11000100 : OUT <= 0;  //2 / 196 = 0
    16'b00000010_11000101 : OUT <= 0;  //2 / 197 = 0
    16'b00000010_11000110 : OUT <= 0;  //2 / 198 = 0
    16'b00000010_11000111 : OUT <= 0;  //2 / 199 = 0
    16'b00000010_11001000 : OUT <= 0;  //2 / 200 = 0
    16'b00000010_11001001 : OUT <= 0;  //2 / 201 = 0
    16'b00000010_11001010 : OUT <= 0;  //2 / 202 = 0
    16'b00000010_11001011 : OUT <= 0;  //2 / 203 = 0
    16'b00000010_11001100 : OUT <= 0;  //2 / 204 = 0
    16'b00000010_11001101 : OUT <= 0;  //2 / 205 = 0
    16'b00000010_11001110 : OUT <= 0;  //2 / 206 = 0
    16'b00000010_11001111 : OUT <= 0;  //2 / 207 = 0
    16'b00000010_11010000 : OUT <= 0;  //2 / 208 = 0
    16'b00000010_11010001 : OUT <= 0;  //2 / 209 = 0
    16'b00000010_11010010 : OUT <= 0;  //2 / 210 = 0
    16'b00000010_11010011 : OUT <= 0;  //2 / 211 = 0
    16'b00000010_11010100 : OUT <= 0;  //2 / 212 = 0
    16'b00000010_11010101 : OUT <= 0;  //2 / 213 = 0
    16'b00000010_11010110 : OUT <= 0;  //2 / 214 = 0
    16'b00000010_11010111 : OUT <= 0;  //2 / 215 = 0
    16'b00000010_11011000 : OUT <= 0;  //2 / 216 = 0
    16'b00000010_11011001 : OUT <= 0;  //2 / 217 = 0
    16'b00000010_11011010 : OUT <= 0;  //2 / 218 = 0
    16'b00000010_11011011 : OUT <= 0;  //2 / 219 = 0
    16'b00000010_11011100 : OUT <= 0;  //2 / 220 = 0
    16'b00000010_11011101 : OUT <= 0;  //2 / 221 = 0
    16'b00000010_11011110 : OUT <= 0;  //2 / 222 = 0
    16'b00000010_11011111 : OUT <= 0;  //2 / 223 = 0
    16'b00000010_11100000 : OUT <= 0;  //2 / 224 = 0
    16'b00000010_11100001 : OUT <= 0;  //2 / 225 = 0
    16'b00000010_11100010 : OUT <= 0;  //2 / 226 = 0
    16'b00000010_11100011 : OUT <= 0;  //2 / 227 = 0
    16'b00000010_11100100 : OUT <= 0;  //2 / 228 = 0
    16'b00000010_11100101 : OUT <= 0;  //2 / 229 = 0
    16'b00000010_11100110 : OUT <= 0;  //2 / 230 = 0
    16'b00000010_11100111 : OUT <= 0;  //2 / 231 = 0
    16'b00000010_11101000 : OUT <= 0;  //2 / 232 = 0
    16'b00000010_11101001 : OUT <= 0;  //2 / 233 = 0
    16'b00000010_11101010 : OUT <= 0;  //2 / 234 = 0
    16'b00000010_11101011 : OUT <= 0;  //2 / 235 = 0
    16'b00000010_11101100 : OUT <= 0;  //2 / 236 = 0
    16'b00000010_11101101 : OUT <= 0;  //2 / 237 = 0
    16'b00000010_11101110 : OUT <= 0;  //2 / 238 = 0
    16'b00000010_11101111 : OUT <= 0;  //2 / 239 = 0
    16'b00000010_11110000 : OUT <= 0;  //2 / 240 = 0
    16'b00000010_11110001 : OUT <= 0;  //2 / 241 = 0
    16'b00000010_11110010 : OUT <= 0;  //2 / 242 = 0
    16'b00000010_11110011 : OUT <= 0;  //2 / 243 = 0
    16'b00000010_11110100 : OUT <= 0;  //2 / 244 = 0
    16'b00000010_11110101 : OUT <= 0;  //2 / 245 = 0
    16'b00000010_11110110 : OUT <= 0;  //2 / 246 = 0
    16'b00000010_11110111 : OUT <= 0;  //2 / 247 = 0
    16'b00000010_11111000 : OUT <= 0;  //2 / 248 = 0
    16'b00000010_11111001 : OUT <= 0;  //2 / 249 = 0
    16'b00000010_11111010 : OUT <= 0;  //2 / 250 = 0
    16'b00000010_11111011 : OUT <= 0;  //2 / 251 = 0
    16'b00000010_11111100 : OUT <= 0;  //2 / 252 = 0
    16'b00000010_11111101 : OUT <= 0;  //2 / 253 = 0
    16'b00000010_11111110 : OUT <= 0;  //2 / 254 = 0
    16'b00000010_11111111 : OUT <= 0;  //2 / 255 = 0
    16'b00000011_00000000 : OUT <= 0;  //3 / 0 = 0
    16'b00000011_00000001 : OUT <= 3;  //3 / 1 = 3
    16'b00000011_00000010 : OUT <= 1;  //3 / 2 = 1
    16'b00000011_00000011 : OUT <= 1;  //3 / 3 = 1
    16'b00000011_00000100 : OUT <= 0;  //3 / 4 = 0
    16'b00000011_00000101 : OUT <= 0;  //3 / 5 = 0
    16'b00000011_00000110 : OUT <= 0;  //3 / 6 = 0
    16'b00000011_00000111 : OUT <= 0;  //3 / 7 = 0
    16'b00000011_00001000 : OUT <= 0;  //3 / 8 = 0
    16'b00000011_00001001 : OUT <= 0;  //3 / 9 = 0
    16'b00000011_00001010 : OUT <= 0;  //3 / 10 = 0
    16'b00000011_00001011 : OUT <= 0;  //3 / 11 = 0
    16'b00000011_00001100 : OUT <= 0;  //3 / 12 = 0
    16'b00000011_00001101 : OUT <= 0;  //3 / 13 = 0
    16'b00000011_00001110 : OUT <= 0;  //3 / 14 = 0
    16'b00000011_00001111 : OUT <= 0;  //3 / 15 = 0
    16'b00000011_00010000 : OUT <= 0;  //3 / 16 = 0
    16'b00000011_00010001 : OUT <= 0;  //3 / 17 = 0
    16'b00000011_00010010 : OUT <= 0;  //3 / 18 = 0
    16'b00000011_00010011 : OUT <= 0;  //3 / 19 = 0
    16'b00000011_00010100 : OUT <= 0;  //3 / 20 = 0
    16'b00000011_00010101 : OUT <= 0;  //3 / 21 = 0
    16'b00000011_00010110 : OUT <= 0;  //3 / 22 = 0
    16'b00000011_00010111 : OUT <= 0;  //3 / 23 = 0
    16'b00000011_00011000 : OUT <= 0;  //3 / 24 = 0
    16'b00000011_00011001 : OUT <= 0;  //3 / 25 = 0
    16'b00000011_00011010 : OUT <= 0;  //3 / 26 = 0
    16'b00000011_00011011 : OUT <= 0;  //3 / 27 = 0
    16'b00000011_00011100 : OUT <= 0;  //3 / 28 = 0
    16'b00000011_00011101 : OUT <= 0;  //3 / 29 = 0
    16'b00000011_00011110 : OUT <= 0;  //3 / 30 = 0
    16'b00000011_00011111 : OUT <= 0;  //3 / 31 = 0
    16'b00000011_00100000 : OUT <= 0;  //3 / 32 = 0
    16'b00000011_00100001 : OUT <= 0;  //3 / 33 = 0
    16'b00000011_00100010 : OUT <= 0;  //3 / 34 = 0
    16'b00000011_00100011 : OUT <= 0;  //3 / 35 = 0
    16'b00000011_00100100 : OUT <= 0;  //3 / 36 = 0
    16'b00000011_00100101 : OUT <= 0;  //3 / 37 = 0
    16'b00000011_00100110 : OUT <= 0;  //3 / 38 = 0
    16'b00000011_00100111 : OUT <= 0;  //3 / 39 = 0
    16'b00000011_00101000 : OUT <= 0;  //3 / 40 = 0
    16'b00000011_00101001 : OUT <= 0;  //3 / 41 = 0
    16'b00000011_00101010 : OUT <= 0;  //3 / 42 = 0
    16'b00000011_00101011 : OUT <= 0;  //3 / 43 = 0
    16'b00000011_00101100 : OUT <= 0;  //3 / 44 = 0
    16'b00000011_00101101 : OUT <= 0;  //3 / 45 = 0
    16'b00000011_00101110 : OUT <= 0;  //3 / 46 = 0
    16'b00000011_00101111 : OUT <= 0;  //3 / 47 = 0
    16'b00000011_00110000 : OUT <= 0;  //3 / 48 = 0
    16'b00000011_00110001 : OUT <= 0;  //3 / 49 = 0
    16'b00000011_00110010 : OUT <= 0;  //3 / 50 = 0
    16'b00000011_00110011 : OUT <= 0;  //3 / 51 = 0
    16'b00000011_00110100 : OUT <= 0;  //3 / 52 = 0
    16'b00000011_00110101 : OUT <= 0;  //3 / 53 = 0
    16'b00000011_00110110 : OUT <= 0;  //3 / 54 = 0
    16'b00000011_00110111 : OUT <= 0;  //3 / 55 = 0
    16'b00000011_00111000 : OUT <= 0;  //3 / 56 = 0
    16'b00000011_00111001 : OUT <= 0;  //3 / 57 = 0
    16'b00000011_00111010 : OUT <= 0;  //3 / 58 = 0
    16'b00000011_00111011 : OUT <= 0;  //3 / 59 = 0
    16'b00000011_00111100 : OUT <= 0;  //3 / 60 = 0
    16'b00000011_00111101 : OUT <= 0;  //3 / 61 = 0
    16'b00000011_00111110 : OUT <= 0;  //3 / 62 = 0
    16'b00000011_00111111 : OUT <= 0;  //3 / 63 = 0
    16'b00000011_01000000 : OUT <= 0;  //3 / 64 = 0
    16'b00000011_01000001 : OUT <= 0;  //3 / 65 = 0
    16'b00000011_01000010 : OUT <= 0;  //3 / 66 = 0
    16'b00000011_01000011 : OUT <= 0;  //3 / 67 = 0
    16'b00000011_01000100 : OUT <= 0;  //3 / 68 = 0
    16'b00000011_01000101 : OUT <= 0;  //3 / 69 = 0
    16'b00000011_01000110 : OUT <= 0;  //3 / 70 = 0
    16'b00000011_01000111 : OUT <= 0;  //3 / 71 = 0
    16'b00000011_01001000 : OUT <= 0;  //3 / 72 = 0
    16'b00000011_01001001 : OUT <= 0;  //3 / 73 = 0
    16'b00000011_01001010 : OUT <= 0;  //3 / 74 = 0
    16'b00000011_01001011 : OUT <= 0;  //3 / 75 = 0
    16'b00000011_01001100 : OUT <= 0;  //3 / 76 = 0
    16'b00000011_01001101 : OUT <= 0;  //3 / 77 = 0
    16'b00000011_01001110 : OUT <= 0;  //3 / 78 = 0
    16'b00000011_01001111 : OUT <= 0;  //3 / 79 = 0
    16'b00000011_01010000 : OUT <= 0;  //3 / 80 = 0
    16'b00000011_01010001 : OUT <= 0;  //3 / 81 = 0
    16'b00000011_01010010 : OUT <= 0;  //3 / 82 = 0
    16'b00000011_01010011 : OUT <= 0;  //3 / 83 = 0
    16'b00000011_01010100 : OUT <= 0;  //3 / 84 = 0
    16'b00000011_01010101 : OUT <= 0;  //3 / 85 = 0
    16'b00000011_01010110 : OUT <= 0;  //3 / 86 = 0
    16'b00000011_01010111 : OUT <= 0;  //3 / 87 = 0
    16'b00000011_01011000 : OUT <= 0;  //3 / 88 = 0
    16'b00000011_01011001 : OUT <= 0;  //3 / 89 = 0
    16'b00000011_01011010 : OUT <= 0;  //3 / 90 = 0
    16'b00000011_01011011 : OUT <= 0;  //3 / 91 = 0
    16'b00000011_01011100 : OUT <= 0;  //3 / 92 = 0
    16'b00000011_01011101 : OUT <= 0;  //3 / 93 = 0
    16'b00000011_01011110 : OUT <= 0;  //3 / 94 = 0
    16'b00000011_01011111 : OUT <= 0;  //3 / 95 = 0
    16'b00000011_01100000 : OUT <= 0;  //3 / 96 = 0
    16'b00000011_01100001 : OUT <= 0;  //3 / 97 = 0
    16'b00000011_01100010 : OUT <= 0;  //3 / 98 = 0
    16'b00000011_01100011 : OUT <= 0;  //3 / 99 = 0
    16'b00000011_01100100 : OUT <= 0;  //3 / 100 = 0
    16'b00000011_01100101 : OUT <= 0;  //3 / 101 = 0
    16'b00000011_01100110 : OUT <= 0;  //3 / 102 = 0
    16'b00000011_01100111 : OUT <= 0;  //3 / 103 = 0
    16'b00000011_01101000 : OUT <= 0;  //3 / 104 = 0
    16'b00000011_01101001 : OUT <= 0;  //3 / 105 = 0
    16'b00000011_01101010 : OUT <= 0;  //3 / 106 = 0
    16'b00000011_01101011 : OUT <= 0;  //3 / 107 = 0
    16'b00000011_01101100 : OUT <= 0;  //3 / 108 = 0
    16'b00000011_01101101 : OUT <= 0;  //3 / 109 = 0
    16'b00000011_01101110 : OUT <= 0;  //3 / 110 = 0
    16'b00000011_01101111 : OUT <= 0;  //3 / 111 = 0
    16'b00000011_01110000 : OUT <= 0;  //3 / 112 = 0
    16'b00000011_01110001 : OUT <= 0;  //3 / 113 = 0
    16'b00000011_01110010 : OUT <= 0;  //3 / 114 = 0
    16'b00000011_01110011 : OUT <= 0;  //3 / 115 = 0
    16'b00000011_01110100 : OUT <= 0;  //3 / 116 = 0
    16'b00000011_01110101 : OUT <= 0;  //3 / 117 = 0
    16'b00000011_01110110 : OUT <= 0;  //3 / 118 = 0
    16'b00000011_01110111 : OUT <= 0;  //3 / 119 = 0
    16'b00000011_01111000 : OUT <= 0;  //3 / 120 = 0
    16'b00000011_01111001 : OUT <= 0;  //3 / 121 = 0
    16'b00000011_01111010 : OUT <= 0;  //3 / 122 = 0
    16'b00000011_01111011 : OUT <= 0;  //3 / 123 = 0
    16'b00000011_01111100 : OUT <= 0;  //3 / 124 = 0
    16'b00000011_01111101 : OUT <= 0;  //3 / 125 = 0
    16'b00000011_01111110 : OUT <= 0;  //3 / 126 = 0
    16'b00000011_01111111 : OUT <= 0;  //3 / 127 = 0
    16'b00000011_10000000 : OUT <= 0;  //3 / 128 = 0
    16'b00000011_10000001 : OUT <= 0;  //3 / 129 = 0
    16'b00000011_10000010 : OUT <= 0;  //3 / 130 = 0
    16'b00000011_10000011 : OUT <= 0;  //3 / 131 = 0
    16'b00000011_10000100 : OUT <= 0;  //3 / 132 = 0
    16'b00000011_10000101 : OUT <= 0;  //3 / 133 = 0
    16'b00000011_10000110 : OUT <= 0;  //3 / 134 = 0
    16'b00000011_10000111 : OUT <= 0;  //3 / 135 = 0
    16'b00000011_10001000 : OUT <= 0;  //3 / 136 = 0
    16'b00000011_10001001 : OUT <= 0;  //3 / 137 = 0
    16'b00000011_10001010 : OUT <= 0;  //3 / 138 = 0
    16'b00000011_10001011 : OUT <= 0;  //3 / 139 = 0
    16'b00000011_10001100 : OUT <= 0;  //3 / 140 = 0
    16'b00000011_10001101 : OUT <= 0;  //3 / 141 = 0
    16'b00000011_10001110 : OUT <= 0;  //3 / 142 = 0
    16'b00000011_10001111 : OUT <= 0;  //3 / 143 = 0
    16'b00000011_10010000 : OUT <= 0;  //3 / 144 = 0
    16'b00000011_10010001 : OUT <= 0;  //3 / 145 = 0
    16'b00000011_10010010 : OUT <= 0;  //3 / 146 = 0
    16'b00000011_10010011 : OUT <= 0;  //3 / 147 = 0
    16'b00000011_10010100 : OUT <= 0;  //3 / 148 = 0
    16'b00000011_10010101 : OUT <= 0;  //3 / 149 = 0
    16'b00000011_10010110 : OUT <= 0;  //3 / 150 = 0
    16'b00000011_10010111 : OUT <= 0;  //3 / 151 = 0
    16'b00000011_10011000 : OUT <= 0;  //3 / 152 = 0
    16'b00000011_10011001 : OUT <= 0;  //3 / 153 = 0
    16'b00000011_10011010 : OUT <= 0;  //3 / 154 = 0
    16'b00000011_10011011 : OUT <= 0;  //3 / 155 = 0
    16'b00000011_10011100 : OUT <= 0;  //3 / 156 = 0
    16'b00000011_10011101 : OUT <= 0;  //3 / 157 = 0
    16'b00000011_10011110 : OUT <= 0;  //3 / 158 = 0
    16'b00000011_10011111 : OUT <= 0;  //3 / 159 = 0
    16'b00000011_10100000 : OUT <= 0;  //3 / 160 = 0
    16'b00000011_10100001 : OUT <= 0;  //3 / 161 = 0
    16'b00000011_10100010 : OUT <= 0;  //3 / 162 = 0
    16'b00000011_10100011 : OUT <= 0;  //3 / 163 = 0
    16'b00000011_10100100 : OUT <= 0;  //3 / 164 = 0
    16'b00000011_10100101 : OUT <= 0;  //3 / 165 = 0
    16'b00000011_10100110 : OUT <= 0;  //3 / 166 = 0
    16'b00000011_10100111 : OUT <= 0;  //3 / 167 = 0
    16'b00000011_10101000 : OUT <= 0;  //3 / 168 = 0
    16'b00000011_10101001 : OUT <= 0;  //3 / 169 = 0
    16'b00000011_10101010 : OUT <= 0;  //3 / 170 = 0
    16'b00000011_10101011 : OUT <= 0;  //3 / 171 = 0
    16'b00000011_10101100 : OUT <= 0;  //3 / 172 = 0
    16'b00000011_10101101 : OUT <= 0;  //3 / 173 = 0
    16'b00000011_10101110 : OUT <= 0;  //3 / 174 = 0
    16'b00000011_10101111 : OUT <= 0;  //3 / 175 = 0
    16'b00000011_10110000 : OUT <= 0;  //3 / 176 = 0
    16'b00000011_10110001 : OUT <= 0;  //3 / 177 = 0
    16'b00000011_10110010 : OUT <= 0;  //3 / 178 = 0
    16'b00000011_10110011 : OUT <= 0;  //3 / 179 = 0
    16'b00000011_10110100 : OUT <= 0;  //3 / 180 = 0
    16'b00000011_10110101 : OUT <= 0;  //3 / 181 = 0
    16'b00000011_10110110 : OUT <= 0;  //3 / 182 = 0
    16'b00000011_10110111 : OUT <= 0;  //3 / 183 = 0
    16'b00000011_10111000 : OUT <= 0;  //3 / 184 = 0
    16'b00000011_10111001 : OUT <= 0;  //3 / 185 = 0
    16'b00000011_10111010 : OUT <= 0;  //3 / 186 = 0
    16'b00000011_10111011 : OUT <= 0;  //3 / 187 = 0
    16'b00000011_10111100 : OUT <= 0;  //3 / 188 = 0
    16'b00000011_10111101 : OUT <= 0;  //3 / 189 = 0
    16'b00000011_10111110 : OUT <= 0;  //3 / 190 = 0
    16'b00000011_10111111 : OUT <= 0;  //3 / 191 = 0
    16'b00000011_11000000 : OUT <= 0;  //3 / 192 = 0
    16'b00000011_11000001 : OUT <= 0;  //3 / 193 = 0
    16'b00000011_11000010 : OUT <= 0;  //3 / 194 = 0
    16'b00000011_11000011 : OUT <= 0;  //3 / 195 = 0
    16'b00000011_11000100 : OUT <= 0;  //3 / 196 = 0
    16'b00000011_11000101 : OUT <= 0;  //3 / 197 = 0
    16'b00000011_11000110 : OUT <= 0;  //3 / 198 = 0
    16'b00000011_11000111 : OUT <= 0;  //3 / 199 = 0
    16'b00000011_11001000 : OUT <= 0;  //3 / 200 = 0
    16'b00000011_11001001 : OUT <= 0;  //3 / 201 = 0
    16'b00000011_11001010 : OUT <= 0;  //3 / 202 = 0
    16'b00000011_11001011 : OUT <= 0;  //3 / 203 = 0
    16'b00000011_11001100 : OUT <= 0;  //3 / 204 = 0
    16'b00000011_11001101 : OUT <= 0;  //3 / 205 = 0
    16'b00000011_11001110 : OUT <= 0;  //3 / 206 = 0
    16'b00000011_11001111 : OUT <= 0;  //3 / 207 = 0
    16'b00000011_11010000 : OUT <= 0;  //3 / 208 = 0
    16'b00000011_11010001 : OUT <= 0;  //3 / 209 = 0
    16'b00000011_11010010 : OUT <= 0;  //3 / 210 = 0
    16'b00000011_11010011 : OUT <= 0;  //3 / 211 = 0
    16'b00000011_11010100 : OUT <= 0;  //3 / 212 = 0
    16'b00000011_11010101 : OUT <= 0;  //3 / 213 = 0
    16'b00000011_11010110 : OUT <= 0;  //3 / 214 = 0
    16'b00000011_11010111 : OUT <= 0;  //3 / 215 = 0
    16'b00000011_11011000 : OUT <= 0;  //3 / 216 = 0
    16'b00000011_11011001 : OUT <= 0;  //3 / 217 = 0
    16'b00000011_11011010 : OUT <= 0;  //3 / 218 = 0
    16'b00000011_11011011 : OUT <= 0;  //3 / 219 = 0
    16'b00000011_11011100 : OUT <= 0;  //3 / 220 = 0
    16'b00000011_11011101 : OUT <= 0;  //3 / 221 = 0
    16'b00000011_11011110 : OUT <= 0;  //3 / 222 = 0
    16'b00000011_11011111 : OUT <= 0;  //3 / 223 = 0
    16'b00000011_11100000 : OUT <= 0;  //3 / 224 = 0
    16'b00000011_11100001 : OUT <= 0;  //3 / 225 = 0
    16'b00000011_11100010 : OUT <= 0;  //3 / 226 = 0
    16'b00000011_11100011 : OUT <= 0;  //3 / 227 = 0
    16'b00000011_11100100 : OUT <= 0;  //3 / 228 = 0
    16'b00000011_11100101 : OUT <= 0;  //3 / 229 = 0
    16'b00000011_11100110 : OUT <= 0;  //3 / 230 = 0
    16'b00000011_11100111 : OUT <= 0;  //3 / 231 = 0
    16'b00000011_11101000 : OUT <= 0;  //3 / 232 = 0
    16'b00000011_11101001 : OUT <= 0;  //3 / 233 = 0
    16'b00000011_11101010 : OUT <= 0;  //3 / 234 = 0
    16'b00000011_11101011 : OUT <= 0;  //3 / 235 = 0
    16'b00000011_11101100 : OUT <= 0;  //3 / 236 = 0
    16'b00000011_11101101 : OUT <= 0;  //3 / 237 = 0
    16'b00000011_11101110 : OUT <= 0;  //3 / 238 = 0
    16'b00000011_11101111 : OUT <= 0;  //3 / 239 = 0
    16'b00000011_11110000 : OUT <= 0;  //3 / 240 = 0
    16'b00000011_11110001 : OUT <= 0;  //3 / 241 = 0
    16'b00000011_11110010 : OUT <= 0;  //3 / 242 = 0
    16'b00000011_11110011 : OUT <= 0;  //3 / 243 = 0
    16'b00000011_11110100 : OUT <= 0;  //3 / 244 = 0
    16'b00000011_11110101 : OUT <= 0;  //3 / 245 = 0
    16'b00000011_11110110 : OUT <= 0;  //3 / 246 = 0
    16'b00000011_11110111 : OUT <= 0;  //3 / 247 = 0
    16'b00000011_11111000 : OUT <= 0;  //3 / 248 = 0
    16'b00000011_11111001 : OUT <= 0;  //3 / 249 = 0
    16'b00000011_11111010 : OUT <= 0;  //3 / 250 = 0
    16'b00000011_11111011 : OUT <= 0;  //3 / 251 = 0
    16'b00000011_11111100 : OUT <= 0;  //3 / 252 = 0
    16'b00000011_11111101 : OUT <= 0;  //3 / 253 = 0
    16'b00000011_11111110 : OUT <= 0;  //3 / 254 = 0
    16'b00000011_11111111 : OUT <= 0;  //3 / 255 = 0
    16'b00000100_00000000 : OUT <= 0;  //4 / 0 = 0
    16'b00000100_00000001 : OUT <= 4;  //4 / 1 = 4
    16'b00000100_00000010 : OUT <= 2;  //4 / 2 = 2
    16'b00000100_00000011 : OUT <= 1;  //4 / 3 = 1
    16'b00000100_00000100 : OUT <= 1;  //4 / 4 = 1
    16'b00000100_00000101 : OUT <= 0;  //4 / 5 = 0
    16'b00000100_00000110 : OUT <= 0;  //4 / 6 = 0
    16'b00000100_00000111 : OUT <= 0;  //4 / 7 = 0
    16'b00000100_00001000 : OUT <= 0;  //4 / 8 = 0
    16'b00000100_00001001 : OUT <= 0;  //4 / 9 = 0
    16'b00000100_00001010 : OUT <= 0;  //4 / 10 = 0
    16'b00000100_00001011 : OUT <= 0;  //4 / 11 = 0
    16'b00000100_00001100 : OUT <= 0;  //4 / 12 = 0
    16'b00000100_00001101 : OUT <= 0;  //4 / 13 = 0
    16'b00000100_00001110 : OUT <= 0;  //4 / 14 = 0
    16'b00000100_00001111 : OUT <= 0;  //4 / 15 = 0
    16'b00000100_00010000 : OUT <= 0;  //4 / 16 = 0
    16'b00000100_00010001 : OUT <= 0;  //4 / 17 = 0
    16'b00000100_00010010 : OUT <= 0;  //4 / 18 = 0
    16'b00000100_00010011 : OUT <= 0;  //4 / 19 = 0
    16'b00000100_00010100 : OUT <= 0;  //4 / 20 = 0
    16'b00000100_00010101 : OUT <= 0;  //4 / 21 = 0
    16'b00000100_00010110 : OUT <= 0;  //4 / 22 = 0
    16'b00000100_00010111 : OUT <= 0;  //4 / 23 = 0
    16'b00000100_00011000 : OUT <= 0;  //4 / 24 = 0
    16'b00000100_00011001 : OUT <= 0;  //4 / 25 = 0
    16'b00000100_00011010 : OUT <= 0;  //4 / 26 = 0
    16'b00000100_00011011 : OUT <= 0;  //4 / 27 = 0
    16'b00000100_00011100 : OUT <= 0;  //4 / 28 = 0
    16'b00000100_00011101 : OUT <= 0;  //4 / 29 = 0
    16'b00000100_00011110 : OUT <= 0;  //4 / 30 = 0
    16'b00000100_00011111 : OUT <= 0;  //4 / 31 = 0
    16'b00000100_00100000 : OUT <= 0;  //4 / 32 = 0
    16'b00000100_00100001 : OUT <= 0;  //4 / 33 = 0
    16'b00000100_00100010 : OUT <= 0;  //4 / 34 = 0
    16'b00000100_00100011 : OUT <= 0;  //4 / 35 = 0
    16'b00000100_00100100 : OUT <= 0;  //4 / 36 = 0
    16'b00000100_00100101 : OUT <= 0;  //4 / 37 = 0
    16'b00000100_00100110 : OUT <= 0;  //4 / 38 = 0
    16'b00000100_00100111 : OUT <= 0;  //4 / 39 = 0
    16'b00000100_00101000 : OUT <= 0;  //4 / 40 = 0
    16'b00000100_00101001 : OUT <= 0;  //4 / 41 = 0
    16'b00000100_00101010 : OUT <= 0;  //4 / 42 = 0
    16'b00000100_00101011 : OUT <= 0;  //4 / 43 = 0
    16'b00000100_00101100 : OUT <= 0;  //4 / 44 = 0
    16'b00000100_00101101 : OUT <= 0;  //4 / 45 = 0
    16'b00000100_00101110 : OUT <= 0;  //4 / 46 = 0
    16'b00000100_00101111 : OUT <= 0;  //4 / 47 = 0
    16'b00000100_00110000 : OUT <= 0;  //4 / 48 = 0
    16'b00000100_00110001 : OUT <= 0;  //4 / 49 = 0
    16'b00000100_00110010 : OUT <= 0;  //4 / 50 = 0
    16'b00000100_00110011 : OUT <= 0;  //4 / 51 = 0
    16'b00000100_00110100 : OUT <= 0;  //4 / 52 = 0
    16'b00000100_00110101 : OUT <= 0;  //4 / 53 = 0
    16'b00000100_00110110 : OUT <= 0;  //4 / 54 = 0
    16'b00000100_00110111 : OUT <= 0;  //4 / 55 = 0
    16'b00000100_00111000 : OUT <= 0;  //4 / 56 = 0
    16'b00000100_00111001 : OUT <= 0;  //4 / 57 = 0
    16'b00000100_00111010 : OUT <= 0;  //4 / 58 = 0
    16'b00000100_00111011 : OUT <= 0;  //4 / 59 = 0
    16'b00000100_00111100 : OUT <= 0;  //4 / 60 = 0
    16'b00000100_00111101 : OUT <= 0;  //4 / 61 = 0
    16'b00000100_00111110 : OUT <= 0;  //4 / 62 = 0
    16'b00000100_00111111 : OUT <= 0;  //4 / 63 = 0
    16'b00000100_01000000 : OUT <= 0;  //4 / 64 = 0
    16'b00000100_01000001 : OUT <= 0;  //4 / 65 = 0
    16'b00000100_01000010 : OUT <= 0;  //4 / 66 = 0
    16'b00000100_01000011 : OUT <= 0;  //4 / 67 = 0
    16'b00000100_01000100 : OUT <= 0;  //4 / 68 = 0
    16'b00000100_01000101 : OUT <= 0;  //4 / 69 = 0
    16'b00000100_01000110 : OUT <= 0;  //4 / 70 = 0
    16'b00000100_01000111 : OUT <= 0;  //4 / 71 = 0
    16'b00000100_01001000 : OUT <= 0;  //4 / 72 = 0
    16'b00000100_01001001 : OUT <= 0;  //4 / 73 = 0
    16'b00000100_01001010 : OUT <= 0;  //4 / 74 = 0
    16'b00000100_01001011 : OUT <= 0;  //4 / 75 = 0
    16'b00000100_01001100 : OUT <= 0;  //4 / 76 = 0
    16'b00000100_01001101 : OUT <= 0;  //4 / 77 = 0
    16'b00000100_01001110 : OUT <= 0;  //4 / 78 = 0
    16'b00000100_01001111 : OUT <= 0;  //4 / 79 = 0
    16'b00000100_01010000 : OUT <= 0;  //4 / 80 = 0
    16'b00000100_01010001 : OUT <= 0;  //4 / 81 = 0
    16'b00000100_01010010 : OUT <= 0;  //4 / 82 = 0
    16'b00000100_01010011 : OUT <= 0;  //4 / 83 = 0
    16'b00000100_01010100 : OUT <= 0;  //4 / 84 = 0
    16'b00000100_01010101 : OUT <= 0;  //4 / 85 = 0
    16'b00000100_01010110 : OUT <= 0;  //4 / 86 = 0
    16'b00000100_01010111 : OUT <= 0;  //4 / 87 = 0
    16'b00000100_01011000 : OUT <= 0;  //4 / 88 = 0
    16'b00000100_01011001 : OUT <= 0;  //4 / 89 = 0
    16'b00000100_01011010 : OUT <= 0;  //4 / 90 = 0
    16'b00000100_01011011 : OUT <= 0;  //4 / 91 = 0
    16'b00000100_01011100 : OUT <= 0;  //4 / 92 = 0
    16'b00000100_01011101 : OUT <= 0;  //4 / 93 = 0
    16'b00000100_01011110 : OUT <= 0;  //4 / 94 = 0
    16'b00000100_01011111 : OUT <= 0;  //4 / 95 = 0
    16'b00000100_01100000 : OUT <= 0;  //4 / 96 = 0
    16'b00000100_01100001 : OUT <= 0;  //4 / 97 = 0
    16'b00000100_01100010 : OUT <= 0;  //4 / 98 = 0
    16'b00000100_01100011 : OUT <= 0;  //4 / 99 = 0
    16'b00000100_01100100 : OUT <= 0;  //4 / 100 = 0
    16'b00000100_01100101 : OUT <= 0;  //4 / 101 = 0
    16'b00000100_01100110 : OUT <= 0;  //4 / 102 = 0
    16'b00000100_01100111 : OUT <= 0;  //4 / 103 = 0
    16'b00000100_01101000 : OUT <= 0;  //4 / 104 = 0
    16'b00000100_01101001 : OUT <= 0;  //4 / 105 = 0
    16'b00000100_01101010 : OUT <= 0;  //4 / 106 = 0
    16'b00000100_01101011 : OUT <= 0;  //4 / 107 = 0
    16'b00000100_01101100 : OUT <= 0;  //4 / 108 = 0
    16'b00000100_01101101 : OUT <= 0;  //4 / 109 = 0
    16'b00000100_01101110 : OUT <= 0;  //4 / 110 = 0
    16'b00000100_01101111 : OUT <= 0;  //4 / 111 = 0
    16'b00000100_01110000 : OUT <= 0;  //4 / 112 = 0
    16'b00000100_01110001 : OUT <= 0;  //4 / 113 = 0
    16'b00000100_01110010 : OUT <= 0;  //4 / 114 = 0
    16'b00000100_01110011 : OUT <= 0;  //4 / 115 = 0
    16'b00000100_01110100 : OUT <= 0;  //4 / 116 = 0
    16'b00000100_01110101 : OUT <= 0;  //4 / 117 = 0
    16'b00000100_01110110 : OUT <= 0;  //4 / 118 = 0
    16'b00000100_01110111 : OUT <= 0;  //4 / 119 = 0
    16'b00000100_01111000 : OUT <= 0;  //4 / 120 = 0
    16'b00000100_01111001 : OUT <= 0;  //4 / 121 = 0
    16'b00000100_01111010 : OUT <= 0;  //4 / 122 = 0
    16'b00000100_01111011 : OUT <= 0;  //4 / 123 = 0
    16'b00000100_01111100 : OUT <= 0;  //4 / 124 = 0
    16'b00000100_01111101 : OUT <= 0;  //4 / 125 = 0
    16'b00000100_01111110 : OUT <= 0;  //4 / 126 = 0
    16'b00000100_01111111 : OUT <= 0;  //4 / 127 = 0
    16'b00000100_10000000 : OUT <= 0;  //4 / 128 = 0
    16'b00000100_10000001 : OUT <= 0;  //4 / 129 = 0
    16'b00000100_10000010 : OUT <= 0;  //4 / 130 = 0
    16'b00000100_10000011 : OUT <= 0;  //4 / 131 = 0
    16'b00000100_10000100 : OUT <= 0;  //4 / 132 = 0
    16'b00000100_10000101 : OUT <= 0;  //4 / 133 = 0
    16'b00000100_10000110 : OUT <= 0;  //4 / 134 = 0
    16'b00000100_10000111 : OUT <= 0;  //4 / 135 = 0
    16'b00000100_10001000 : OUT <= 0;  //4 / 136 = 0
    16'b00000100_10001001 : OUT <= 0;  //4 / 137 = 0
    16'b00000100_10001010 : OUT <= 0;  //4 / 138 = 0
    16'b00000100_10001011 : OUT <= 0;  //4 / 139 = 0
    16'b00000100_10001100 : OUT <= 0;  //4 / 140 = 0
    16'b00000100_10001101 : OUT <= 0;  //4 / 141 = 0
    16'b00000100_10001110 : OUT <= 0;  //4 / 142 = 0
    16'b00000100_10001111 : OUT <= 0;  //4 / 143 = 0
    16'b00000100_10010000 : OUT <= 0;  //4 / 144 = 0
    16'b00000100_10010001 : OUT <= 0;  //4 / 145 = 0
    16'b00000100_10010010 : OUT <= 0;  //4 / 146 = 0
    16'b00000100_10010011 : OUT <= 0;  //4 / 147 = 0
    16'b00000100_10010100 : OUT <= 0;  //4 / 148 = 0
    16'b00000100_10010101 : OUT <= 0;  //4 / 149 = 0
    16'b00000100_10010110 : OUT <= 0;  //4 / 150 = 0
    16'b00000100_10010111 : OUT <= 0;  //4 / 151 = 0
    16'b00000100_10011000 : OUT <= 0;  //4 / 152 = 0
    16'b00000100_10011001 : OUT <= 0;  //4 / 153 = 0
    16'b00000100_10011010 : OUT <= 0;  //4 / 154 = 0
    16'b00000100_10011011 : OUT <= 0;  //4 / 155 = 0
    16'b00000100_10011100 : OUT <= 0;  //4 / 156 = 0
    16'b00000100_10011101 : OUT <= 0;  //4 / 157 = 0
    16'b00000100_10011110 : OUT <= 0;  //4 / 158 = 0
    16'b00000100_10011111 : OUT <= 0;  //4 / 159 = 0
    16'b00000100_10100000 : OUT <= 0;  //4 / 160 = 0
    16'b00000100_10100001 : OUT <= 0;  //4 / 161 = 0
    16'b00000100_10100010 : OUT <= 0;  //4 / 162 = 0
    16'b00000100_10100011 : OUT <= 0;  //4 / 163 = 0
    16'b00000100_10100100 : OUT <= 0;  //4 / 164 = 0
    16'b00000100_10100101 : OUT <= 0;  //4 / 165 = 0
    16'b00000100_10100110 : OUT <= 0;  //4 / 166 = 0
    16'b00000100_10100111 : OUT <= 0;  //4 / 167 = 0
    16'b00000100_10101000 : OUT <= 0;  //4 / 168 = 0
    16'b00000100_10101001 : OUT <= 0;  //4 / 169 = 0
    16'b00000100_10101010 : OUT <= 0;  //4 / 170 = 0
    16'b00000100_10101011 : OUT <= 0;  //4 / 171 = 0
    16'b00000100_10101100 : OUT <= 0;  //4 / 172 = 0
    16'b00000100_10101101 : OUT <= 0;  //4 / 173 = 0
    16'b00000100_10101110 : OUT <= 0;  //4 / 174 = 0
    16'b00000100_10101111 : OUT <= 0;  //4 / 175 = 0
    16'b00000100_10110000 : OUT <= 0;  //4 / 176 = 0
    16'b00000100_10110001 : OUT <= 0;  //4 / 177 = 0
    16'b00000100_10110010 : OUT <= 0;  //4 / 178 = 0
    16'b00000100_10110011 : OUT <= 0;  //4 / 179 = 0
    16'b00000100_10110100 : OUT <= 0;  //4 / 180 = 0
    16'b00000100_10110101 : OUT <= 0;  //4 / 181 = 0
    16'b00000100_10110110 : OUT <= 0;  //4 / 182 = 0
    16'b00000100_10110111 : OUT <= 0;  //4 / 183 = 0
    16'b00000100_10111000 : OUT <= 0;  //4 / 184 = 0
    16'b00000100_10111001 : OUT <= 0;  //4 / 185 = 0
    16'b00000100_10111010 : OUT <= 0;  //4 / 186 = 0
    16'b00000100_10111011 : OUT <= 0;  //4 / 187 = 0
    16'b00000100_10111100 : OUT <= 0;  //4 / 188 = 0
    16'b00000100_10111101 : OUT <= 0;  //4 / 189 = 0
    16'b00000100_10111110 : OUT <= 0;  //4 / 190 = 0
    16'b00000100_10111111 : OUT <= 0;  //4 / 191 = 0
    16'b00000100_11000000 : OUT <= 0;  //4 / 192 = 0
    16'b00000100_11000001 : OUT <= 0;  //4 / 193 = 0
    16'b00000100_11000010 : OUT <= 0;  //4 / 194 = 0
    16'b00000100_11000011 : OUT <= 0;  //4 / 195 = 0
    16'b00000100_11000100 : OUT <= 0;  //4 / 196 = 0
    16'b00000100_11000101 : OUT <= 0;  //4 / 197 = 0
    16'b00000100_11000110 : OUT <= 0;  //4 / 198 = 0
    16'b00000100_11000111 : OUT <= 0;  //4 / 199 = 0
    16'b00000100_11001000 : OUT <= 0;  //4 / 200 = 0
    16'b00000100_11001001 : OUT <= 0;  //4 / 201 = 0
    16'b00000100_11001010 : OUT <= 0;  //4 / 202 = 0
    16'b00000100_11001011 : OUT <= 0;  //4 / 203 = 0
    16'b00000100_11001100 : OUT <= 0;  //4 / 204 = 0
    16'b00000100_11001101 : OUT <= 0;  //4 / 205 = 0
    16'b00000100_11001110 : OUT <= 0;  //4 / 206 = 0
    16'b00000100_11001111 : OUT <= 0;  //4 / 207 = 0
    16'b00000100_11010000 : OUT <= 0;  //4 / 208 = 0
    16'b00000100_11010001 : OUT <= 0;  //4 / 209 = 0
    16'b00000100_11010010 : OUT <= 0;  //4 / 210 = 0
    16'b00000100_11010011 : OUT <= 0;  //4 / 211 = 0
    16'b00000100_11010100 : OUT <= 0;  //4 / 212 = 0
    16'b00000100_11010101 : OUT <= 0;  //4 / 213 = 0
    16'b00000100_11010110 : OUT <= 0;  //4 / 214 = 0
    16'b00000100_11010111 : OUT <= 0;  //4 / 215 = 0
    16'b00000100_11011000 : OUT <= 0;  //4 / 216 = 0
    16'b00000100_11011001 : OUT <= 0;  //4 / 217 = 0
    16'b00000100_11011010 : OUT <= 0;  //4 / 218 = 0
    16'b00000100_11011011 : OUT <= 0;  //4 / 219 = 0
    16'b00000100_11011100 : OUT <= 0;  //4 / 220 = 0
    16'b00000100_11011101 : OUT <= 0;  //4 / 221 = 0
    16'b00000100_11011110 : OUT <= 0;  //4 / 222 = 0
    16'b00000100_11011111 : OUT <= 0;  //4 / 223 = 0
    16'b00000100_11100000 : OUT <= 0;  //4 / 224 = 0
    16'b00000100_11100001 : OUT <= 0;  //4 / 225 = 0
    16'b00000100_11100010 : OUT <= 0;  //4 / 226 = 0
    16'b00000100_11100011 : OUT <= 0;  //4 / 227 = 0
    16'b00000100_11100100 : OUT <= 0;  //4 / 228 = 0
    16'b00000100_11100101 : OUT <= 0;  //4 / 229 = 0
    16'b00000100_11100110 : OUT <= 0;  //4 / 230 = 0
    16'b00000100_11100111 : OUT <= 0;  //4 / 231 = 0
    16'b00000100_11101000 : OUT <= 0;  //4 / 232 = 0
    16'b00000100_11101001 : OUT <= 0;  //4 / 233 = 0
    16'b00000100_11101010 : OUT <= 0;  //4 / 234 = 0
    16'b00000100_11101011 : OUT <= 0;  //4 / 235 = 0
    16'b00000100_11101100 : OUT <= 0;  //4 / 236 = 0
    16'b00000100_11101101 : OUT <= 0;  //4 / 237 = 0
    16'b00000100_11101110 : OUT <= 0;  //4 / 238 = 0
    16'b00000100_11101111 : OUT <= 0;  //4 / 239 = 0
    16'b00000100_11110000 : OUT <= 0;  //4 / 240 = 0
    16'b00000100_11110001 : OUT <= 0;  //4 / 241 = 0
    16'b00000100_11110010 : OUT <= 0;  //4 / 242 = 0
    16'b00000100_11110011 : OUT <= 0;  //4 / 243 = 0
    16'b00000100_11110100 : OUT <= 0;  //4 / 244 = 0
    16'b00000100_11110101 : OUT <= 0;  //4 / 245 = 0
    16'b00000100_11110110 : OUT <= 0;  //4 / 246 = 0
    16'b00000100_11110111 : OUT <= 0;  //4 / 247 = 0
    16'b00000100_11111000 : OUT <= 0;  //4 / 248 = 0
    16'b00000100_11111001 : OUT <= 0;  //4 / 249 = 0
    16'b00000100_11111010 : OUT <= 0;  //4 / 250 = 0
    16'b00000100_11111011 : OUT <= 0;  //4 / 251 = 0
    16'b00000100_11111100 : OUT <= 0;  //4 / 252 = 0
    16'b00000100_11111101 : OUT <= 0;  //4 / 253 = 0
    16'b00000100_11111110 : OUT <= 0;  //4 / 254 = 0
    16'b00000100_11111111 : OUT <= 0;  //4 / 255 = 0
    16'b00000101_00000000 : OUT <= 0;  //5 / 0 = 0
    16'b00000101_00000001 : OUT <= 5;  //5 / 1 = 5
    16'b00000101_00000010 : OUT <= 2;  //5 / 2 = 2
    16'b00000101_00000011 : OUT <= 1;  //5 / 3 = 1
    16'b00000101_00000100 : OUT <= 1;  //5 / 4 = 1
    16'b00000101_00000101 : OUT <= 1;  //5 / 5 = 1
    16'b00000101_00000110 : OUT <= 0;  //5 / 6 = 0
    16'b00000101_00000111 : OUT <= 0;  //5 / 7 = 0
    16'b00000101_00001000 : OUT <= 0;  //5 / 8 = 0
    16'b00000101_00001001 : OUT <= 0;  //5 / 9 = 0
    16'b00000101_00001010 : OUT <= 0;  //5 / 10 = 0
    16'b00000101_00001011 : OUT <= 0;  //5 / 11 = 0
    16'b00000101_00001100 : OUT <= 0;  //5 / 12 = 0
    16'b00000101_00001101 : OUT <= 0;  //5 / 13 = 0
    16'b00000101_00001110 : OUT <= 0;  //5 / 14 = 0
    16'b00000101_00001111 : OUT <= 0;  //5 / 15 = 0
    16'b00000101_00010000 : OUT <= 0;  //5 / 16 = 0
    16'b00000101_00010001 : OUT <= 0;  //5 / 17 = 0
    16'b00000101_00010010 : OUT <= 0;  //5 / 18 = 0
    16'b00000101_00010011 : OUT <= 0;  //5 / 19 = 0
    16'b00000101_00010100 : OUT <= 0;  //5 / 20 = 0
    16'b00000101_00010101 : OUT <= 0;  //5 / 21 = 0
    16'b00000101_00010110 : OUT <= 0;  //5 / 22 = 0
    16'b00000101_00010111 : OUT <= 0;  //5 / 23 = 0
    16'b00000101_00011000 : OUT <= 0;  //5 / 24 = 0
    16'b00000101_00011001 : OUT <= 0;  //5 / 25 = 0
    16'b00000101_00011010 : OUT <= 0;  //5 / 26 = 0
    16'b00000101_00011011 : OUT <= 0;  //5 / 27 = 0
    16'b00000101_00011100 : OUT <= 0;  //5 / 28 = 0
    16'b00000101_00011101 : OUT <= 0;  //5 / 29 = 0
    16'b00000101_00011110 : OUT <= 0;  //5 / 30 = 0
    16'b00000101_00011111 : OUT <= 0;  //5 / 31 = 0
    16'b00000101_00100000 : OUT <= 0;  //5 / 32 = 0
    16'b00000101_00100001 : OUT <= 0;  //5 / 33 = 0
    16'b00000101_00100010 : OUT <= 0;  //5 / 34 = 0
    16'b00000101_00100011 : OUT <= 0;  //5 / 35 = 0
    16'b00000101_00100100 : OUT <= 0;  //5 / 36 = 0
    16'b00000101_00100101 : OUT <= 0;  //5 / 37 = 0
    16'b00000101_00100110 : OUT <= 0;  //5 / 38 = 0
    16'b00000101_00100111 : OUT <= 0;  //5 / 39 = 0
    16'b00000101_00101000 : OUT <= 0;  //5 / 40 = 0
    16'b00000101_00101001 : OUT <= 0;  //5 / 41 = 0
    16'b00000101_00101010 : OUT <= 0;  //5 / 42 = 0
    16'b00000101_00101011 : OUT <= 0;  //5 / 43 = 0
    16'b00000101_00101100 : OUT <= 0;  //5 / 44 = 0
    16'b00000101_00101101 : OUT <= 0;  //5 / 45 = 0
    16'b00000101_00101110 : OUT <= 0;  //5 / 46 = 0
    16'b00000101_00101111 : OUT <= 0;  //5 / 47 = 0
    16'b00000101_00110000 : OUT <= 0;  //5 / 48 = 0
    16'b00000101_00110001 : OUT <= 0;  //5 / 49 = 0
    16'b00000101_00110010 : OUT <= 0;  //5 / 50 = 0
    16'b00000101_00110011 : OUT <= 0;  //5 / 51 = 0
    16'b00000101_00110100 : OUT <= 0;  //5 / 52 = 0
    16'b00000101_00110101 : OUT <= 0;  //5 / 53 = 0
    16'b00000101_00110110 : OUT <= 0;  //5 / 54 = 0
    16'b00000101_00110111 : OUT <= 0;  //5 / 55 = 0
    16'b00000101_00111000 : OUT <= 0;  //5 / 56 = 0
    16'b00000101_00111001 : OUT <= 0;  //5 / 57 = 0
    16'b00000101_00111010 : OUT <= 0;  //5 / 58 = 0
    16'b00000101_00111011 : OUT <= 0;  //5 / 59 = 0
    16'b00000101_00111100 : OUT <= 0;  //5 / 60 = 0
    16'b00000101_00111101 : OUT <= 0;  //5 / 61 = 0
    16'b00000101_00111110 : OUT <= 0;  //5 / 62 = 0
    16'b00000101_00111111 : OUT <= 0;  //5 / 63 = 0
    16'b00000101_01000000 : OUT <= 0;  //5 / 64 = 0
    16'b00000101_01000001 : OUT <= 0;  //5 / 65 = 0
    16'b00000101_01000010 : OUT <= 0;  //5 / 66 = 0
    16'b00000101_01000011 : OUT <= 0;  //5 / 67 = 0
    16'b00000101_01000100 : OUT <= 0;  //5 / 68 = 0
    16'b00000101_01000101 : OUT <= 0;  //5 / 69 = 0
    16'b00000101_01000110 : OUT <= 0;  //5 / 70 = 0
    16'b00000101_01000111 : OUT <= 0;  //5 / 71 = 0
    16'b00000101_01001000 : OUT <= 0;  //5 / 72 = 0
    16'b00000101_01001001 : OUT <= 0;  //5 / 73 = 0
    16'b00000101_01001010 : OUT <= 0;  //5 / 74 = 0
    16'b00000101_01001011 : OUT <= 0;  //5 / 75 = 0
    16'b00000101_01001100 : OUT <= 0;  //5 / 76 = 0
    16'b00000101_01001101 : OUT <= 0;  //5 / 77 = 0
    16'b00000101_01001110 : OUT <= 0;  //5 / 78 = 0
    16'b00000101_01001111 : OUT <= 0;  //5 / 79 = 0
    16'b00000101_01010000 : OUT <= 0;  //5 / 80 = 0
    16'b00000101_01010001 : OUT <= 0;  //5 / 81 = 0
    16'b00000101_01010010 : OUT <= 0;  //5 / 82 = 0
    16'b00000101_01010011 : OUT <= 0;  //5 / 83 = 0
    16'b00000101_01010100 : OUT <= 0;  //5 / 84 = 0
    16'b00000101_01010101 : OUT <= 0;  //5 / 85 = 0
    16'b00000101_01010110 : OUT <= 0;  //5 / 86 = 0
    16'b00000101_01010111 : OUT <= 0;  //5 / 87 = 0
    16'b00000101_01011000 : OUT <= 0;  //5 / 88 = 0
    16'b00000101_01011001 : OUT <= 0;  //5 / 89 = 0
    16'b00000101_01011010 : OUT <= 0;  //5 / 90 = 0
    16'b00000101_01011011 : OUT <= 0;  //5 / 91 = 0
    16'b00000101_01011100 : OUT <= 0;  //5 / 92 = 0
    16'b00000101_01011101 : OUT <= 0;  //5 / 93 = 0
    16'b00000101_01011110 : OUT <= 0;  //5 / 94 = 0
    16'b00000101_01011111 : OUT <= 0;  //5 / 95 = 0
    16'b00000101_01100000 : OUT <= 0;  //5 / 96 = 0
    16'b00000101_01100001 : OUT <= 0;  //5 / 97 = 0
    16'b00000101_01100010 : OUT <= 0;  //5 / 98 = 0
    16'b00000101_01100011 : OUT <= 0;  //5 / 99 = 0
    16'b00000101_01100100 : OUT <= 0;  //5 / 100 = 0
    16'b00000101_01100101 : OUT <= 0;  //5 / 101 = 0
    16'b00000101_01100110 : OUT <= 0;  //5 / 102 = 0
    16'b00000101_01100111 : OUT <= 0;  //5 / 103 = 0
    16'b00000101_01101000 : OUT <= 0;  //5 / 104 = 0
    16'b00000101_01101001 : OUT <= 0;  //5 / 105 = 0
    16'b00000101_01101010 : OUT <= 0;  //5 / 106 = 0
    16'b00000101_01101011 : OUT <= 0;  //5 / 107 = 0
    16'b00000101_01101100 : OUT <= 0;  //5 / 108 = 0
    16'b00000101_01101101 : OUT <= 0;  //5 / 109 = 0
    16'b00000101_01101110 : OUT <= 0;  //5 / 110 = 0
    16'b00000101_01101111 : OUT <= 0;  //5 / 111 = 0
    16'b00000101_01110000 : OUT <= 0;  //5 / 112 = 0
    16'b00000101_01110001 : OUT <= 0;  //5 / 113 = 0
    16'b00000101_01110010 : OUT <= 0;  //5 / 114 = 0
    16'b00000101_01110011 : OUT <= 0;  //5 / 115 = 0
    16'b00000101_01110100 : OUT <= 0;  //5 / 116 = 0
    16'b00000101_01110101 : OUT <= 0;  //5 / 117 = 0
    16'b00000101_01110110 : OUT <= 0;  //5 / 118 = 0
    16'b00000101_01110111 : OUT <= 0;  //5 / 119 = 0
    16'b00000101_01111000 : OUT <= 0;  //5 / 120 = 0
    16'b00000101_01111001 : OUT <= 0;  //5 / 121 = 0
    16'b00000101_01111010 : OUT <= 0;  //5 / 122 = 0
    16'b00000101_01111011 : OUT <= 0;  //5 / 123 = 0
    16'b00000101_01111100 : OUT <= 0;  //5 / 124 = 0
    16'b00000101_01111101 : OUT <= 0;  //5 / 125 = 0
    16'b00000101_01111110 : OUT <= 0;  //5 / 126 = 0
    16'b00000101_01111111 : OUT <= 0;  //5 / 127 = 0
    16'b00000101_10000000 : OUT <= 0;  //5 / 128 = 0
    16'b00000101_10000001 : OUT <= 0;  //5 / 129 = 0
    16'b00000101_10000010 : OUT <= 0;  //5 / 130 = 0
    16'b00000101_10000011 : OUT <= 0;  //5 / 131 = 0
    16'b00000101_10000100 : OUT <= 0;  //5 / 132 = 0
    16'b00000101_10000101 : OUT <= 0;  //5 / 133 = 0
    16'b00000101_10000110 : OUT <= 0;  //5 / 134 = 0
    16'b00000101_10000111 : OUT <= 0;  //5 / 135 = 0
    16'b00000101_10001000 : OUT <= 0;  //5 / 136 = 0
    16'b00000101_10001001 : OUT <= 0;  //5 / 137 = 0
    16'b00000101_10001010 : OUT <= 0;  //5 / 138 = 0
    16'b00000101_10001011 : OUT <= 0;  //5 / 139 = 0
    16'b00000101_10001100 : OUT <= 0;  //5 / 140 = 0
    16'b00000101_10001101 : OUT <= 0;  //5 / 141 = 0
    16'b00000101_10001110 : OUT <= 0;  //5 / 142 = 0
    16'b00000101_10001111 : OUT <= 0;  //5 / 143 = 0
    16'b00000101_10010000 : OUT <= 0;  //5 / 144 = 0
    16'b00000101_10010001 : OUT <= 0;  //5 / 145 = 0
    16'b00000101_10010010 : OUT <= 0;  //5 / 146 = 0
    16'b00000101_10010011 : OUT <= 0;  //5 / 147 = 0
    16'b00000101_10010100 : OUT <= 0;  //5 / 148 = 0
    16'b00000101_10010101 : OUT <= 0;  //5 / 149 = 0
    16'b00000101_10010110 : OUT <= 0;  //5 / 150 = 0
    16'b00000101_10010111 : OUT <= 0;  //5 / 151 = 0
    16'b00000101_10011000 : OUT <= 0;  //5 / 152 = 0
    16'b00000101_10011001 : OUT <= 0;  //5 / 153 = 0
    16'b00000101_10011010 : OUT <= 0;  //5 / 154 = 0
    16'b00000101_10011011 : OUT <= 0;  //5 / 155 = 0
    16'b00000101_10011100 : OUT <= 0;  //5 / 156 = 0
    16'b00000101_10011101 : OUT <= 0;  //5 / 157 = 0
    16'b00000101_10011110 : OUT <= 0;  //5 / 158 = 0
    16'b00000101_10011111 : OUT <= 0;  //5 / 159 = 0
    16'b00000101_10100000 : OUT <= 0;  //5 / 160 = 0
    16'b00000101_10100001 : OUT <= 0;  //5 / 161 = 0
    16'b00000101_10100010 : OUT <= 0;  //5 / 162 = 0
    16'b00000101_10100011 : OUT <= 0;  //5 / 163 = 0
    16'b00000101_10100100 : OUT <= 0;  //5 / 164 = 0
    16'b00000101_10100101 : OUT <= 0;  //5 / 165 = 0
    16'b00000101_10100110 : OUT <= 0;  //5 / 166 = 0
    16'b00000101_10100111 : OUT <= 0;  //5 / 167 = 0
    16'b00000101_10101000 : OUT <= 0;  //5 / 168 = 0
    16'b00000101_10101001 : OUT <= 0;  //5 / 169 = 0
    16'b00000101_10101010 : OUT <= 0;  //5 / 170 = 0
    16'b00000101_10101011 : OUT <= 0;  //5 / 171 = 0
    16'b00000101_10101100 : OUT <= 0;  //5 / 172 = 0
    16'b00000101_10101101 : OUT <= 0;  //5 / 173 = 0
    16'b00000101_10101110 : OUT <= 0;  //5 / 174 = 0
    16'b00000101_10101111 : OUT <= 0;  //5 / 175 = 0
    16'b00000101_10110000 : OUT <= 0;  //5 / 176 = 0
    16'b00000101_10110001 : OUT <= 0;  //5 / 177 = 0
    16'b00000101_10110010 : OUT <= 0;  //5 / 178 = 0
    16'b00000101_10110011 : OUT <= 0;  //5 / 179 = 0
    16'b00000101_10110100 : OUT <= 0;  //5 / 180 = 0
    16'b00000101_10110101 : OUT <= 0;  //5 / 181 = 0
    16'b00000101_10110110 : OUT <= 0;  //5 / 182 = 0
    16'b00000101_10110111 : OUT <= 0;  //5 / 183 = 0
    16'b00000101_10111000 : OUT <= 0;  //5 / 184 = 0
    16'b00000101_10111001 : OUT <= 0;  //5 / 185 = 0
    16'b00000101_10111010 : OUT <= 0;  //5 / 186 = 0
    16'b00000101_10111011 : OUT <= 0;  //5 / 187 = 0
    16'b00000101_10111100 : OUT <= 0;  //5 / 188 = 0
    16'b00000101_10111101 : OUT <= 0;  //5 / 189 = 0
    16'b00000101_10111110 : OUT <= 0;  //5 / 190 = 0
    16'b00000101_10111111 : OUT <= 0;  //5 / 191 = 0
    16'b00000101_11000000 : OUT <= 0;  //5 / 192 = 0
    16'b00000101_11000001 : OUT <= 0;  //5 / 193 = 0
    16'b00000101_11000010 : OUT <= 0;  //5 / 194 = 0
    16'b00000101_11000011 : OUT <= 0;  //5 / 195 = 0
    16'b00000101_11000100 : OUT <= 0;  //5 / 196 = 0
    16'b00000101_11000101 : OUT <= 0;  //5 / 197 = 0
    16'b00000101_11000110 : OUT <= 0;  //5 / 198 = 0
    16'b00000101_11000111 : OUT <= 0;  //5 / 199 = 0
    16'b00000101_11001000 : OUT <= 0;  //5 / 200 = 0
    16'b00000101_11001001 : OUT <= 0;  //5 / 201 = 0
    16'b00000101_11001010 : OUT <= 0;  //5 / 202 = 0
    16'b00000101_11001011 : OUT <= 0;  //5 / 203 = 0
    16'b00000101_11001100 : OUT <= 0;  //5 / 204 = 0
    16'b00000101_11001101 : OUT <= 0;  //5 / 205 = 0
    16'b00000101_11001110 : OUT <= 0;  //5 / 206 = 0
    16'b00000101_11001111 : OUT <= 0;  //5 / 207 = 0
    16'b00000101_11010000 : OUT <= 0;  //5 / 208 = 0
    16'b00000101_11010001 : OUT <= 0;  //5 / 209 = 0
    16'b00000101_11010010 : OUT <= 0;  //5 / 210 = 0
    16'b00000101_11010011 : OUT <= 0;  //5 / 211 = 0
    16'b00000101_11010100 : OUT <= 0;  //5 / 212 = 0
    16'b00000101_11010101 : OUT <= 0;  //5 / 213 = 0
    16'b00000101_11010110 : OUT <= 0;  //5 / 214 = 0
    16'b00000101_11010111 : OUT <= 0;  //5 / 215 = 0
    16'b00000101_11011000 : OUT <= 0;  //5 / 216 = 0
    16'b00000101_11011001 : OUT <= 0;  //5 / 217 = 0
    16'b00000101_11011010 : OUT <= 0;  //5 / 218 = 0
    16'b00000101_11011011 : OUT <= 0;  //5 / 219 = 0
    16'b00000101_11011100 : OUT <= 0;  //5 / 220 = 0
    16'b00000101_11011101 : OUT <= 0;  //5 / 221 = 0
    16'b00000101_11011110 : OUT <= 0;  //5 / 222 = 0
    16'b00000101_11011111 : OUT <= 0;  //5 / 223 = 0
    16'b00000101_11100000 : OUT <= 0;  //5 / 224 = 0
    16'b00000101_11100001 : OUT <= 0;  //5 / 225 = 0
    16'b00000101_11100010 : OUT <= 0;  //5 / 226 = 0
    16'b00000101_11100011 : OUT <= 0;  //5 / 227 = 0
    16'b00000101_11100100 : OUT <= 0;  //5 / 228 = 0
    16'b00000101_11100101 : OUT <= 0;  //5 / 229 = 0
    16'b00000101_11100110 : OUT <= 0;  //5 / 230 = 0
    16'b00000101_11100111 : OUT <= 0;  //5 / 231 = 0
    16'b00000101_11101000 : OUT <= 0;  //5 / 232 = 0
    16'b00000101_11101001 : OUT <= 0;  //5 / 233 = 0
    16'b00000101_11101010 : OUT <= 0;  //5 / 234 = 0
    16'b00000101_11101011 : OUT <= 0;  //5 / 235 = 0
    16'b00000101_11101100 : OUT <= 0;  //5 / 236 = 0
    16'b00000101_11101101 : OUT <= 0;  //5 / 237 = 0
    16'b00000101_11101110 : OUT <= 0;  //5 / 238 = 0
    16'b00000101_11101111 : OUT <= 0;  //5 / 239 = 0
    16'b00000101_11110000 : OUT <= 0;  //5 / 240 = 0
    16'b00000101_11110001 : OUT <= 0;  //5 / 241 = 0
    16'b00000101_11110010 : OUT <= 0;  //5 / 242 = 0
    16'b00000101_11110011 : OUT <= 0;  //5 / 243 = 0
    16'b00000101_11110100 : OUT <= 0;  //5 / 244 = 0
    16'b00000101_11110101 : OUT <= 0;  //5 / 245 = 0
    16'b00000101_11110110 : OUT <= 0;  //5 / 246 = 0
    16'b00000101_11110111 : OUT <= 0;  //5 / 247 = 0
    16'b00000101_11111000 : OUT <= 0;  //5 / 248 = 0
    16'b00000101_11111001 : OUT <= 0;  //5 / 249 = 0
    16'b00000101_11111010 : OUT <= 0;  //5 / 250 = 0
    16'b00000101_11111011 : OUT <= 0;  //5 / 251 = 0
    16'b00000101_11111100 : OUT <= 0;  //5 / 252 = 0
    16'b00000101_11111101 : OUT <= 0;  //5 / 253 = 0
    16'b00000101_11111110 : OUT <= 0;  //5 / 254 = 0
    16'b00000101_11111111 : OUT <= 0;  //5 / 255 = 0
    16'b00000110_00000000 : OUT <= 0;  //6 / 0 = 0
    16'b00000110_00000001 : OUT <= 6;  //6 / 1 = 6
    16'b00000110_00000010 : OUT <= 3;  //6 / 2 = 3
    16'b00000110_00000011 : OUT <= 2;  //6 / 3 = 2
    16'b00000110_00000100 : OUT <= 1;  //6 / 4 = 1
    16'b00000110_00000101 : OUT <= 1;  //6 / 5 = 1
    16'b00000110_00000110 : OUT <= 1;  //6 / 6 = 1
    16'b00000110_00000111 : OUT <= 0;  //6 / 7 = 0
    16'b00000110_00001000 : OUT <= 0;  //6 / 8 = 0
    16'b00000110_00001001 : OUT <= 0;  //6 / 9 = 0
    16'b00000110_00001010 : OUT <= 0;  //6 / 10 = 0
    16'b00000110_00001011 : OUT <= 0;  //6 / 11 = 0
    16'b00000110_00001100 : OUT <= 0;  //6 / 12 = 0
    16'b00000110_00001101 : OUT <= 0;  //6 / 13 = 0
    16'b00000110_00001110 : OUT <= 0;  //6 / 14 = 0
    16'b00000110_00001111 : OUT <= 0;  //6 / 15 = 0
    16'b00000110_00010000 : OUT <= 0;  //6 / 16 = 0
    16'b00000110_00010001 : OUT <= 0;  //6 / 17 = 0
    16'b00000110_00010010 : OUT <= 0;  //6 / 18 = 0
    16'b00000110_00010011 : OUT <= 0;  //6 / 19 = 0
    16'b00000110_00010100 : OUT <= 0;  //6 / 20 = 0
    16'b00000110_00010101 : OUT <= 0;  //6 / 21 = 0
    16'b00000110_00010110 : OUT <= 0;  //6 / 22 = 0
    16'b00000110_00010111 : OUT <= 0;  //6 / 23 = 0
    16'b00000110_00011000 : OUT <= 0;  //6 / 24 = 0
    16'b00000110_00011001 : OUT <= 0;  //6 / 25 = 0
    16'b00000110_00011010 : OUT <= 0;  //6 / 26 = 0
    16'b00000110_00011011 : OUT <= 0;  //6 / 27 = 0
    16'b00000110_00011100 : OUT <= 0;  //6 / 28 = 0
    16'b00000110_00011101 : OUT <= 0;  //6 / 29 = 0
    16'b00000110_00011110 : OUT <= 0;  //6 / 30 = 0
    16'b00000110_00011111 : OUT <= 0;  //6 / 31 = 0
    16'b00000110_00100000 : OUT <= 0;  //6 / 32 = 0
    16'b00000110_00100001 : OUT <= 0;  //6 / 33 = 0
    16'b00000110_00100010 : OUT <= 0;  //6 / 34 = 0
    16'b00000110_00100011 : OUT <= 0;  //6 / 35 = 0
    16'b00000110_00100100 : OUT <= 0;  //6 / 36 = 0
    16'b00000110_00100101 : OUT <= 0;  //6 / 37 = 0
    16'b00000110_00100110 : OUT <= 0;  //6 / 38 = 0
    16'b00000110_00100111 : OUT <= 0;  //6 / 39 = 0
    16'b00000110_00101000 : OUT <= 0;  //6 / 40 = 0
    16'b00000110_00101001 : OUT <= 0;  //6 / 41 = 0
    16'b00000110_00101010 : OUT <= 0;  //6 / 42 = 0
    16'b00000110_00101011 : OUT <= 0;  //6 / 43 = 0
    16'b00000110_00101100 : OUT <= 0;  //6 / 44 = 0
    16'b00000110_00101101 : OUT <= 0;  //6 / 45 = 0
    16'b00000110_00101110 : OUT <= 0;  //6 / 46 = 0
    16'b00000110_00101111 : OUT <= 0;  //6 / 47 = 0
    16'b00000110_00110000 : OUT <= 0;  //6 / 48 = 0
    16'b00000110_00110001 : OUT <= 0;  //6 / 49 = 0
    16'b00000110_00110010 : OUT <= 0;  //6 / 50 = 0
    16'b00000110_00110011 : OUT <= 0;  //6 / 51 = 0
    16'b00000110_00110100 : OUT <= 0;  //6 / 52 = 0
    16'b00000110_00110101 : OUT <= 0;  //6 / 53 = 0
    16'b00000110_00110110 : OUT <= 0;  //6 / 54 = 0
    16'b00000110_00110111 : OUT <= 0;  //6 / 55 = 0
    16'b00000110_00111000 : OUT <= 0;  //6 / 56 = 0
    16'b00000110_00111001 : OUT <= 0;  //6 / 57 = 0
    16'b00000110_00111010 : OUT <= 0;  //6 / 58 = 0
    16'b00000110_00111011 : OUT <= 0;  //6 / 59 = 0
    16'b00000110_00111100 : OUT <= 0;  //6 / 60 = 0
    16'b00000110_00111101 : OUT <= 0;  //6 / 61 = 0
    16'b00000110_00111110 : OUT <= 0;  //6 / 62 = 0
    16'b00000110_00111111 : OUT <= 0;  //6 / 63 = 0
    16'b00000110_01000000 : OUT <= 0;  //6 / 64 = 0
    16'b00000110_01000001 : OUT <= 0;  //6 / 65 = 0
    16'b00000110_01000010 : OUT <= 0;  //6 / 66 = 0
    16'b00000110_01000011 : OUT <= 0;  //6 / 67 = 0
    16'b00000110_01000100 : OUT <= 0;  //6 / 68 = 0
    16'b00000110_01000101 : OUT <= 0;  //6 / 69 = 0
    16'b00000110_01000110 : OUT <= 0;  //6 / 70 = 0
    16'b00000110_01000111 : OUT <= 0;  //6 / 71 = 0
    16'b00000110_01001000 : OUT <= 0;  //6 / 72 = 0
    16'b00000110_01001001 : OUT <= 0;  //6 / 73 = 0
    16'b00000110_01001010 : OUT <= 0;  //6 / 74 = 0
    16'b00000110_01001011 : OUT <= 0;  //6 / 75 = 0
    16'b00000110_01001100 : OUT <= 0;  //6 / 76 = 0
    16'b00000110_01001101 : OUT <= 0;  //6 / 77 = 0
    16'b00000110_01001110 : OUT <= 0;  //6 / 78 = 0
    16'b00000110_01001111 : OUT <= 0;  //6 / 79 = 0
    16'b00000110_01010000 : OUT <= 0;  //6 / 80 = 0
    16'b00000110_01010001 : OUT <= 0;  //6 / 81 = 0
    16'b00000110_01010010 : OUT <= 0;  //6 / 82 = 0
    16'b00000110_01010011 : OUT <= 0;  //6 / 83 = 0
    16'b00000110_01010100 : OUT <= 0;  //6 / 84 = 0
    16'b00000110_01010101 : OUT <= 0;  //6 / 85 = 0
    16'b00000110_01010110 : OUT <= 0;  //6 / 86 = 0
    16'b00000110_01010111 : OUT <= 0;  //6 / 87 = 0
    16'b00000110_01011000 : OUT <= 0;  //6 / 88 = 0
    16'b00000110_01011001 : OUT <= 0;  //6 / 89 = 0
    16'b00000110_01011010 : OUT <= 0;  //6 / 90 = 0
    16'b00000110_01011011 : OUT <= 0;  //6 / 91 = 0
    16'b00000110_01011100 : OUT <= 0;  //6 / 92 = 0
    16'b00000110_01011101 : OUT <= 0;  //6 / 93 = 0
    16'b00000110_01011110 : OUT <= 0;  //6 / 94 = 0
    16'b00000110_01011111 : OUT <= 0;  //6 / 95 = 0
    16'b00000110_01100000 : OUT <= 0;  //6 / 96 = 0
    16'b00000110_01100001 : OUT <= 0;  //6 / 97 = 0
    16'b00000110_01100010 : OUT <= 0;  //6 / 98 = 0
    16'b00000110_01100011 : OUT <= 0;  //6 / 99 = 0
    16'b00000110_01100100 : OUT <= 0;  //6 / 100 = 0
    16'b00000110_01100101 : OUT <= 0;  //6 / 101 = 0
    16'b00000110_01100110 : OUT <= 0;  //6 / 102 = 0
    16'b00000110_01100111 : OUT <= 0;  //6 / 103 = 0
    16'b00000110_01101000 : OUT <= 0;  //6 / 104 = 0
    16'b00000110_01101001 : OUT <= 0;  //6 / 105 = 0
    16'b00000110_01101010 : OUT <= 0;  //6 / 106 = 0
    16'b00000110_01101011 : OUT <= 0;  //6 / 107 = 0
    16'b00000110_01101100 : OUT <= 0;  //6 / 108 = 0
    16'b00000110_01101101 : OUT <= 0;  //6 / 109 = 0
    16'b00000110_01101110 : OUT <= 0;  //6 / 110 = 0
    16'b00000110_01101111 : OUT <= 0;  //6 / 111 = 0
    16'b00000110_01110000 : OUT <= 0;  //6 / 112 = 0
    16'b00000110_01110001 : OUT <= 0;  //6 / 113 = 0
    16'b00000110_01110010 : OUT <= 0;  //6 / 114 = 0
    16'b00000110_01110011 : OUT <= 0;  //6 / 115 = 0
    16'b00000110_01110100 : OUT <= 0;  //6 / 116 = 0
    16'b00000110_01110101 : OUT <= 0;  //6 / 117 = 0
    16'b00000110_01110110 : OUT <= 0;  //6 / 118 = 0
    16'b00000110_01110111 : OUT <= 0;  //6 / 119 = 0
    16'b00000110_01111000 : OUT <= 0;  //6 / 120 = 0
    16'b00000110_01111001 : OUT <= 0;  //6 / 121 = 0
    16'b00000110_01111010 : OUT <= 0;  //6 / 122 = 0
    16'b00000110_01111011 : OUT <= 0;  //6 / 123 = 0
    16'b00000110_01111100 : OUT <= 0;  //6 / 124 = 0
    16'b00000110_01111101 : OUT <= 0;  //6 / 125 = 0
    16'b00000110_01111110 : OUT <= 0;  //6 / 126 = 0
    16'b00000110_01111111 : OUT <= 0;  //6 / 127 = 0
    16'b00000110_10000000 : OUT <= 0;  //6 / 128 = 0
    16'b00000110_10000001 : OUT <= 0;  //6 / 129 = 0
    16'b00000110_10000010 : OUT <= 0;  //6 / 130 = 0
    16'b00000110_10000011 : OUT <= 0;  //6 / 131 = 0
    16'b00000110_10000100 : OUT <= 0;  //6 / 132 = 0
    16'b00000110_10000101 : OUT <= 0;  //6 / 133 = 0
    16'b00000110_10000110 : OUT <= 0;  //6 / 134 = 0
    16'b00000110_10000111 : OUT <= 0;  //6 / 135 = 0
    16'b00000110_10001000 : OUT <= 0;  //6 / 136 = 0
    16'b00000110_10001001 : OUT <= 0;  //6 / 137 = 0
    16'b00000110_10001010 : OUT <= 0;  //6 / 138 = 0
    16'b00000110_10001011 : OUT <= 0;  //6 / 139 = 0
    16'b00000110_10001100 : OUT <= 0;  //6 / 140 = 0
    16'b00000110_10001101 : OUT <= 0;  //6 / 141 = 0
    16'b00000110_10001110 : OUT <= 0;  //6 / 142 = 0
    16'b00000110_10001111 : OUT <= 0;  //6 / 143 = 0
    16'b00000110_10010000 : OUT <= 0;  //6 / 144 = 0
    16'b00000110_10010001 : OUT <= 0;  //6 / 145 = 0
    16'b00000110_10010010 : OUT <= 0;  //6 / 146 = 0
    16'b00000110_10010011 : OUT <= 0;  //6 / 147 = 0
    16'b00000110_10010100 : OUT <= 0;  //6 / 148 = 0
    16'b00000110_10010101 : OUT <= 0;  //6 / 149 = 0
    16'b00000110_10010110 : OUT <= 0;  //6 / 150 = 0
    16'b00000110_10010111 : OUT <= 0;  //6 / 151 = 0
    16'b00000110_10011000 : OUT <= 0;  //6 / 152 = 0
    16'b00000110_10011001 : OUT <= 0;  //6 / 153 = 0
    16'b00000110_10011010 : OUT <= 0;  //6 / 154 = 0
    16'b00000110_10011011 : OUT <= 0;  //6 / 155 = 0
    16'b00000110_10011100 : OUT <= 0;  //6 / 156 = 0
    16'b00000110_10011101 : OUT <= 0;  //6 / 157 = 0
    16'b00000110_10011110 : OUT <= 0;  //6 / 158 = 0
    16'b00000110_10011111 : OUT <= 0;  //6 / 159 = 0
    16'b00000110_10100000 : OUT <= 0;  //6 / 160 = 0
    16'b00000110_10100001 : OUT <= 0;  //6 / 161 = 0
    16'b00000110_10100010 : OUT <= 0;  //6 / 162 = 0
    16'b00000110_10100011 : OUT <= 0;  //6 / 163 = 0
    16'b00000110_10100100 : OUT <= 0;  //6 / 164 = 0
    16'b00000110_10100101 : OUT <= 0;  //6 / 165 = 0
    16'b00000110_10100110 : OUT <= 0;  //6 / 166 = 0
    16'b00000110_10100111 : OUT <= 0;  //6 / 167 = 0
    16'b00000110_10101000 : OUT <= 0;  //6 / 168 = 0
    16'b00000110_10101001 : OUT <= 0;  //6 / 169 = 0
    16'b00000110_10101010 : OUT <= 0;  //6 / 170 = 0
    16'b00000110_10101011 : OUT <= 0;  //6 / 171 = 0
    16'b00000110_10101100 : OUT <= 0;  //6 / 172 = 0
    16'b00000110_10101101 : OUT <= 0;  //6 / 173 = 0
    16'b00000110_10101110 : OUT <= 0;  //6 / 174 = 0
    16'b00000110_10101111 : OUT <= 0;  //6 / 175 = 0
    16'b00000110_10110000 : OUT <= 0;  //6 / 176 = 0
    16'b00000110_10110001 : OUT <= 0;  //6 / 177 = 0
    16'b00000110_10110010 : OUT <= 0;  //6 / 178 = 0
    16'b00000110_10110011 : OUT <= 0;  //6 / 179 = 0
    16'b00000110_10110100 : OUT <= 0;  //6 / 180 = 0
    16'b00000110_10110101 : OUT <= 0;  //6 / 181 = 0
    16'b00000110_10110110 : OUT <= 0;  //6 / 182 = 0
    16'b00000110_10110111 : OUT <= 0;  //6 / 183 = 0
    16'b00000110_10111000 : OUT <= 0;  //6 / 184 = 0
    16'b00000110_10111001 : OUT <= 0;  //6 / 185 = 0
    16'b00000110_10111010 : OUT <= 0;  //6 / 186 = 0
    16'b00000110_10111011 : OUT <= 0;  //6 / 187 = 0
    16'b00000110_10111100 : OUT <= 0;  //6 / 188 = 0
    16'b00000110_10111101 : OUT <= 0;  //6 / 189 = 0
    16'b00000110_10111110 : OUT <= 0;  //6 / 190 = 0
    16'b00000110_10111111 : OUT <= 0;  //6 / 191 = 0
    16'b00000110_11000000 : OUT <= 0;  //6 / 192 = 0
    16'b00000110_11000001 : OUT <= 0;  //6 / 193 = 0
    16'b00000110_11000010 : OUT <= 0;  //6 / 194 = 0
    16'b00000110_11000011 : OUT <= 0;  //6 / 195 = 0
    16'b00000110_11000100 : OUT <= 0;  //6 / 196 = 0
    16'b00000110_11000101 : OUT <= 0;  //6 / 197 = 0
    16'b00000110_11000110 : OUT <= 0;  //6 / 198 = 0
    16'b00000110_11000111 : OUT <= 0;  //6 / 199 = 0
    16'b00000110_11001000 : OUT <= 0;  //6 / 200 = 0
    16'b00000110_11001001 : OUT <= 0;  //6 / 201 = 0
    16'b00000110_11001010 : OUT <= 0;  //6 / 202 = 0
    16'b00000110_11001011 : OUT <= 0;  //6 / 203 = 0
    16'b00000110_11001100 : OUT <= 0;  //6 / 204 = 0
    16'b00000110_11001101 : OUT <= 0;  //6 / 205 = 0
    16'b00000110_11001110 : OUT <= 0;  //6 / 206 = 0
    16'b00000110_11001111 : OUT <= 0;  //6 / 207 = 0
    16'b00000110_11010000 : OUT <= 0;  //6 / 208 = 0
    16'b00000110_11010001 : OUT <= 0;  //6 / 209 = 0
    16'b00000110_11010010 : OUT <= 0;  //6 / 210 = 0
    16'b00000110_11010011 : OUT <= 0;  //6 / 211 = 0
    16'b00000110_11010100 : OUT <= 0;  //6 / 212 = 0
    16'b00000110_11010101 : OUT <= 0;  //6 / 213 = 0
    16'b00000110_11010110 : OUT <= 0;  //6 / 214 = 0
    16'b00000110_11010111 : OUT <= 0;  //6 / 215 = 0
    16'b00000110_11011000 : OUT <= 0;  //6 / 216 = 0
    16'b00000110_11011001 : OUT <= 0;  //6 / 217 = 0
    16'b00000110_11011010 : OUT <= 0;  //6 / 218 = 0
    16'b00000110_11011011 : OUT <= 0;  //6 / 219 = 0
    16'b00000110_11011100 : OUT <= 0;  //6 / 220 = 0
    16'b00000110_11011101 : OUT <= 0;  //6 / 221 = 0
    16'b00000110_11011110 : OUT <= 0;  //6 / 222 = 0
    16'b00000110_11011111 : OUT <= 0;  //6 / 223 = 0
    16'b00000110_11100000 : OUT <= 0;  //6 / 224 = 0
    16'b00000110_11100001 : OUT <= 0;  //6 / 225 = 0
    16'b00000110_11100010 : OUT <= 0;  //6 / 226 = 0
    16'b00000110_11100011 : OUT <= 0;  //6 / 227 = 0
    16'b00000110_11100100 : OUT <= 0;  //6 / 228 = 0
    16'b00000110_11100101 : OUT <= 0;  //6 / 229 = 0
    16'b00000110_11100110 : OUT <= 0;  //6 / 230 = 0
    16'b00000110_11100111 : OUT <= 0;  //6 / 231 = 0
    16'b00000110_11101000 : OUT <= 0;  //6 / 232 = 0
    16'b00000110_11101001 : OUT <= 0;  //6 / 233 = 0
    16'b00000110_11101010 : OUT <= 0;  //6 / 234 = 0
    16'b00000110_11101011 : OUT <= 0;  //6 / 235 = 0
    16'b00000110_11101100 : OUT <= 0;  //6 / 236 = 0
    16'b00000110_11101101 : OUT <= 0;  //6 / 237 = 0
    16'b00000110_11101110 : OUT <= 0;  //6 / 238 = 0
    16'b00000110_11101111 : OUT <= 0;  //6 / 239 = 0
    16'b00000110_11110000 : OUT <= 0;  //6 / 240 = 0
    16'b00000110_11110001 : OUT <= 0;  //6 / 241 = 0
    16'b00000110_11110010 : OUT <= 0;  //6 / 242 = 0
    16'b00000110_11110011 : OUT <= 0;  //6 / 243 = 0
    16'b00000110_11110100 : OUT <= 0;  //6 / 244 = 0
    16'b00000110_11110101 : OUT <= 0;  //6 / 245 = 0
    16'b00000110_11110110 : OUT <= 0;  //6 / 246 = 0
    16'b00000110_11110111 : OUT <= 0;  //6 / 247 = 0
    16'b00000110_11111000 : OUT <= 0;  //6 / 248 = 0
    16'b00000110_11111001 : OUT <= 0;  //6 / 249 = 0
    16'b00000110_11111010 : OUT <= 0;  //6 / 250 = 0
    16'b00000110_11111011 : OUT <= 0;  //6 / 251 = 0
    16'b00000110_11111100 : OUT <= 0;  //6 / 252 = 0
    16'b00000110_11111101 : OUT <= 0;  //6 / 253 = 0
    16'b00000110_11111110 : OUT <= 0;  //6 / 254 = 0
    16'b00000110_11111111 : OUT <= 0;  //6 / 255 = 0
    16'b00000111_00000000 : OUT <= 0;  //7 / 0 = 0
    16'b00000111_00000001 : OUT <= 7;  //7 / 1 = 7
    16'b00000111_00000010 : OUT <= 3;  //7 / 2 = 3
    16'b00000111_00000011 : OUT <= 2;  //7 / 3 = 2
    16'b00000111_00000100 : OUT <= 1;  //7 / 4 = 1
    16'b00000111_00000101 : OUT <= 1;  //7 / 5 = 1
    16'b00000111_00000110 : OUT <= 1;  //7 / 6 = 1
    16'b00000111_00000111 : OUT <= 1;  //7 / 7 = 1
    16'b00000111_00001000 : OUT <= 0;  //7 / 8 = 0
    16'b00000111_00001001 : OUT <= 0;  //7 / 9 = 0
    16'b00000111_00001010 : OUT <= 0;  //7 / 10 = 0
    16'b00000111_00001011 : OUT <= 0;  //7 / 11 = 0
    16'b00000111_00001100 : OUT <= 0;  //7 / 12 = 0
    16'b00000111_00001101 : OUT <= 0;  //7 / 13 = 0
    16'b00000111_00001110 : OUT <= 0;  //7 / 14 = 0
    16'b00000111_00001111 : OUT <= 0;  //7 / 15 = 0
    16'b00000111_00010000 : OUT <= 0;  //7 / 16 = 0
    16'b00000111_00010001 : OUT <= 0;  //7 / 17 = 0
    16'b00000111_00010010 : OUT <= 0;  //7 / 18 = 0
    16'b00000111_00010011 : OUT <= 0;  //7 / 19 = 0
    16'b00000111_00010100 : OUT <= 0;  //7 / 20 = 0
    16'b00000111_00010101 : OUT <= 0;  //7 / 21 = 0
    16'b00000111_00010110 : OUT <= 0;  //7 / 22 = 0
    16'b00000111_00010111 : OUT <= 0;  //7 / 23 = 0
    16'b00000111_00011000 : OUT <= 0;  //7 / 24 = 0
    16'b00000111_00011001 : OUT <= 0;  //7 / 25 = 0
    16'b00000111_00011010 : OUT <= 0;  //7 / 26 = 0
    16'b00000111_00011011 : OUT <= 0;  //7 / 27 = 0
    16'b00000111_00011100 : OUT <= 0;  //7 / 28 = 0
    16'b00000111_00011101 : OUT <= 0;  //7 / 29 = 0
    16'b00000111_00011110 : OUT <= 0;  //7 / 30 = 0
    16'b00000111_00011111 : OUT <= 0;  //7 / 31 = 0
    16'b00000111_00100000 : OUT <= 0;  //7 / 32 = 0
    16'b00000111_00100001 : OUT <= 0;  //7 / 33 = 0
    16'b00000111_00100010 : OUT <= 0;  //7 / 34 = 0
    16'b00000111_00100011 : OUT <= 0;  //7 / 35 = 0
    16'b00000111_00100100 : OUT <= 0;  //7 / 36 = 0
    16'b00000111_00100101 : OUT <= 0;  //7 / 37 = 0
    16'b00000111_00100110 : OUT <= 0;  //7 / 38 = 0
    16'b00000111_00100111 : OUT <= 0;  //7 / 39 = 0
    16'b00000111_00101000 : OUT <= 0;  //7 / 40 = 0
    16'b00000111_00101001 : OUT <= 0;  //7 / 41 = 0
    16'b00000111_00101010 : OUT <= 0;  //7 / 42 = 0
    16'b00000111_00101011 : OUT <= 0;  //7 / 43 = 0
    16'b00000111_00101100 : OUT <= 0;  //7 / 44 = 0
    16'b00000111_00101101 : OUT <= 0;  //7 / 45 = 0
    16'b00000111_00101110 : OUT <= 0;  //7 / 46 = 0
    16'b00000111_00101111 : OUT <= 0;  //7 / 47 = 0
    16'b00000111_00110000 : OUT <= 0;  //7 / 48 = 0
    16'b00000111_00110001 : OUT <= 0;  //7 / 49 = 0
    16'b00000111_00110010 : OUT <= 0;  //7 / 50 = 0
    16'b00000111_00110011 : OUT <= 0;  //7 / 51 = 0
    16'b00000111_00110100 : OUT <= 0;  //7 / 52 = 0
    16'b00000111_00110101 : OUT <= 0;  //7 / 53 = 0
    16'b00000111_00110110 : OUT <= 0;  //7 / 54 = 0
    16'b00000111_00110111 : OUT <= 0;  //7 / 55 = 0
    16'b00000111_00111000 : OUT <= 0;  //7 / 56 = 0
    16'b00000111_00111001 : OUT <= 0;  //7 / 57 = 0
    16'b00000111_00111010 : OUT <= 0;  //7 / 58 = 0
    16'b00000111_00111011 : OUT <= 0;  //7 / 59 = 0
    16'b00000111_00111100 : OUT <= 0;  //7 / 60 = 0
    16'b00000111_00111101 : OUT <= 0;  //7 / 61 = 0
    16'b00000111_00111110 : OUT <= 0;  //7 / 62 = 0
    16'b00000111_00111111 : OUT <= 0;  //7 / 63 = 0
    16'b00000111_01000000 : OUT <= 0;  //7 / 64 = 0
    16'b00000111_01000001 : OUT <= 0;  //7 / 65 = 0
    16'b00000111_01000010 : OUT <= 0;  //7 / 66 = 0
    16'b00000111_01000011 : OUT <= 0;  //7 / 67 = 0
    16'b00000111_01000100 : OUT <= 0;  //7 / 68 = 0
    16'b00000111_01000101 : OUT <= 0;  //7 / 69 = 0
    16'b00000111_01000110 : OUT <= 0;  //7 / 70 = 0
    16'b00000111_01000111 : OUT <= 0;  //7 / 71 = 0
    16'b00000111_01001000 : OUT <= 0;  //7 / 72 = 0
    16'b00000111_01001001 : OUT <= 0;  //7 / 73 = 0
    16'b00000111_01001010 : OUT <= 0;  //7 / 74 = 0
    16'b00000111_01001011 : OUT <= 0;  //7 / 75 = 0
    16'b00000111_01001100 : OUT <= 0;  //7 / 76 = 0
    16'b00000111_01001101 : OUT <= 0;  //7 / 77 = 0
    16'b00000111_01001110 : OUT <= 0;  //7 / 78 = 0
    16'b00000111_01001111 : OUT <= 0;  //7 / 79 = 0
    16'b00000111_01010000 : OUT <= 0;  //7 / 80 = 0
    16'b00000111_01010001 : OUT <= 0;  //7 / 81 = 0
    16'b00000111_01010010 : OUT <= 0;  //7 / 82 = 0
    16'b00000111_01010011 : OUT <= 0;  //7 / 83 = 0
    16'b00000111_01010100 : OUT <= 0;  //7 / 84 = 0
    16'b00000111_01010101 : OUT <= 0;  //7 / 85 = 0
    16'b00000111_01010110 : OUT <= 0;  //7 / 86 = 0
    16'b00000111_01010111 : OUT <= 0;  //7 / 87 = 0
    16'b00000111_01011000 : OUT <= 0;  //7 / 88 = 0
    16'b00000111_01011001 : OUT <= 0;  //7 / 89 = 0
    16'b00000111_01011010 : OUT <= 0;  //7 / 90 = 0
    16'b00000111_01011011 : OUT <= 0;  //7 / 91 = 0
    16'b00000111_01011100 : OUT <= 0;  //7 / 92 = 0
    16'b00000111_01011101 : OUT <= 0;  //7 / 93 = 0
    16'b00000111_01011110 : OUT <= 0;  //7 / 94 = 0
    16'b00000111_01011111 : OUT <= 0;  //7 / 95 = 0
    16'b00000111_01100000 : OUT <= 0;  //7 / 96 = 0
    16'b00000111_01100001 : OUT <= 0;  //7 / 97 = 0
    16'b00000111_01100010 : OUT <= 0;  //7 / 98 = 0
    16'b00000111_01100011 : OUT <= 0;  //7 / 99 = 0
    16'b00000111_01100100 : OUT <= 0;  //7 / 100 = 0
    16'b00000111_01100101 : OUT <= 0;  //7 / 101 = 0
    16'b00000111_01100110 : OUT <= 0;  //7 / 102 = 0
    16'b00000111_01100111 : OUT <= 0;  //7 / 103 = 0
    16'b00000111_01101000 : OUT <= 0;  //7 / 104 = 0
    16'b00000111_01101001 : OUT <= 0;  //7 / 105 = 0
    16'b00000111_01101010 : OUT <= 0;  //7 / 106 = 0
    16'b00000111_01101011 : OUT <= 0;  //7 / 107 = 0
    16'b00000111_01101100 : OUT <= 0;  //7 / 108 = 0
    16'b00000111_01101101 : OUT <= 0;  //7 / 109 = 0
    16'b00000111_01101110 : OUT <= 0;  //7 / 110 = 0
    16'b00000111_01101111 : OUT <= 0;  //7 / 111 = 0
    16'b00000111_01110000 : OUT <= 0;  //7 / 112 = 0
    16'b00000111_01110001 : OUT <= 0;  //7 / 113 = 0
    16'b00000111_01110010 : OUT <= 0;  //7 / 114 = 0
    16'b00000111_01110011 : OUT <= 0;  //7 / 115 = 0
    16'b00000111_01110100 : OUT <= 0;  //7 / 116 = 0
    16'b00000111_01110101 : OUT <= 0;  //7 / 117 = 0
    16'b00000111_01110110 : OUT <= 0;  //7 / 118 = 0
    16'b00000111_01110111 : OUT <= 0;  //7 / 119 = 0
    16'b00000111_01111000 : OUT <= 0;  //7 / 120 = 0
    16'b00000111_01111001 : OUT <= 0;  //7 / 121 = 0
    16'b00000111_01111010 : OUT <= 0;  //7 / 122 = 0
    16'b00000111_01111011 : OUT <= 0;  //7 / 123 = 0
    16'b00000111_01111100 : OUT <= 0;  //7 / 124 = 0
    16'b00000111_01111101 : OUT <= 0;  //7 / 125 = 0
    16'b00000111_01111110 : OUT <= 0;  //7 / 126 = 0
    16'b00000111_01111111 : OUT <= 0;  //7 / 127 = 0
    16'b00000111_10000000 : OUT <= 0;  //7 / 128 = 0
    16'b00000111_10000001 : OUT <= 0;  //7 / 129 = 0
    16'b00000111_10000010 : OUT <= 0;  //7 / 130 = 0
    16'b00000111_10000011 : OUT <= 0;  //7 / 131 = 0
    16'b00000111_10000100 : OUT <= 0;  //7 / 132 = 0
    16'b00000111_10000101 : OUT <= 0;  //7 / 133 = 0
    16'b00000111_10000110 : OUT <= 0;  //7 / 134 = 0
    16'b00000111_10000111 : OUT <= 0;  //7 / 135 = 0
    16'b00000111_10001000 : OUT <= 0;  //7 / 136 = 0
    16'b00000111_10001001 : OUT <= 0;  //7 / 137 = 0
    16'b00000111_10001010 : OUT <= 0;  //7 / 138 = 0
    16'b00000111_10001011 : OUT <= 0;  //7 / 139 = 0
    16'b00000111_10001100 : OUT <= 0;  //7 / 140 = 0
    16'b00000111_10001101 : OUT <= 0;  //7 / 141 = 0
    16'b00000111_10001110 : OUT <= 0;  //7 / 142 = 0
    16'b00000111_10001111 : OUT <= 0;  //7 / 143 = 0
    16'b00000111_10010000 : OUT <= 0;  //7 / 144 = 0
    16'b00000111_10010001 : OUT <= 0;  //7 / 145 = 0
    16'b00000111_10010010 : OUT <= 0;  //7 / 146 = 0
    16'b00000111_10010011 : OUT <= 0;  //7 / 147 = 0
    16'b00000111_10010100 : OUT <= 0;  //7 / 148 = 0
    16'b00000111_10010101 : OUT <= 0;  //7 / 149 = 0
    16'b00000111_10010110 : OUT <= 0;  //7 / 150 = 0
    16'b00000111_10010111 : OUT <= 0;  //7 / 151 = 0
    16'b00000111_10011000 : OUT <= 0;  //7 / 152 = 0
    16'b00000111_10011001 : OUT <= 0;  //7 / 153 = 0
    16'b00000111_10011010 : OUT <= 0;  //7 / 154 = 0
    16'b00000111_10011011 : OUT <= 0;  //7 / 155 = 0
    16'b00000111_10011100 : OUT <= 0;  //7 / 156 = 0
    16'b00000111_10011101 : OUT <= 0;  //7 / 157 = 0
    16'b00000111_10011110 : OUT <= 0;  //7 / 158 = 0
    16'b00000111_10011111 : OUT <= 0;  //7 / 159 = 0
    16'b00000111_10100000 : OUT <= 0;  //7 / 160 = 0
    16'b00000111_10100001 : OUT <= 0;  //7 / 161 = 0
    16'b00000111_10100010 : OUT <= 0;  //7 / 162 = 0
    16'b00000111_10100011 : OUT <= 0;  //7 / 163 = 0
    16'b00000111_10100100 : OUT <= 0;  //7 / 164 = 0
    16'b00000111_10100101 : OUT <= 0;  //7 / 165 = 0
    16'b00000111_10100110 : OUT <= 0;  //7 / 166 = 0
    16'b00000111_10100111 : OUT <= 0;  //7 / 167 = 0
    16'b00000111_10101000 : OUT <= 0;  //7 / 168 = 0
    16'b00000111_10101001 : OUT <= 0;  //7 / 169 = 0
    16'b00000111_10101010 : OUT <= 0;  //7 / 170 = 0
    16'b00000111_10101011 : OUT <= 0;  //7 / 171 = 0
    16'b00000111_10101100 : OUT <= 0;  //7 / 172 = 0
    16'b00000111_10101101 : OUT <= 0;  //7 / 173 = 0
    16'b00000111_10101110 : OUT <= 0;  //7 / 174 = 0
    16'b00000111_10101111 : OUT <= 0;  //7 / 175 = 0
    16'b00000111_10110000 : OUT <= 0;  //7 / 176 = 0
    16'b00000111_10110001 : OUT <= 0;  //7 / 177 = 0
    16'b00000111_10110010 : OUT <= 0;  //7 / 178 = 0
    16'b00000111_10110011 : OUT <= 0;  //7 / 179 = 0
    16'b00000111_10110100 : OUT <= 0;  //7 / 180 = 0
    16'b00000111_10110101 : OUT <= 0;  //7 / 181 = 0
    16'b00000111_10110110 : OUT <= 0;  //7 / 182 = 0
    16'b00000111_10110111 : OUT <= 0;  //7 / 183 = 0
    16'b00000111_10111000 : OUT <= 0;  //7 / 184 = 0
    16'b00000111_10111001 : OUT <= 0;  //7 / 185 = 0
    16'b00000111_10111010 : OUT <= 0;  //7 / 186 = 0
    16'b00000111_10111011 : OUT <= 0;  //7 / 187 = 0
    16'b00000111_10111100 : OUT <= 0;  //7 / 188 = 0
    16'b00000111_10111101 : OUT <= 0;  //7 / 189 = 0
    16'b00000111_10111110 : OUT <= 0;  //7 / 190 = 0
    16'b00000111_10111111 : OUT <= 0;  //7 / 191 = 0
    16'b00000111_11000000 : OUT <= 0;  //7 / 192 = 0
    16'b00000111_11000001 : OUT <= 0;  //7 / 193 = 0
    16'b00000111_11000010 : OUT <= 0;  //7 / 194 = 0
    16'b00000111_11000011 : OUT <= 0;  //7 / 195 = 0
    16'b00000111_11000100 : OUT <= 0;  //7 / 196 = 0
    16'b00000111_11000101 : OUT <= 0;  //7 / 197 = 0
    16'b00000111_11000110 : OUT <= 0;  //7 / 198 = 0
    16'b00000111_11000111 : OUT <= 0;  //7 / 199 = 0
    16'b00000111_11001000 : OUT <= 0;  //7 / 200 = 0
    16'b00000111_11001001 : OUT <= 0;  //7 / 201 = 0
    16'b00000111_11001010 : OUT <= 0;  //7 / 202 = 0
    16'b00000111_11001011 : OUT <= 0;  //7 / 203 = 0
    16'b00000111_11001100 : OUT <= 0;  //7 / 204 = 0
    16'b00000111_11001101 : OUT <= 0;  //7 / 205 = 0
    16'b00000111_11001110 : OUT <= 0;  //7 / 206 = 0
    16'b00000111_11001111 : OUT <= 0;  //7 / 207 = 0
    16'b00000111_11010000 : OUT <= 0;  //7 / 208 = 0
    16'b00000111_11010001 : OUT <= 0;  //7 / 209 = 0
    16'b00000111_11010010 : OUT <= 0;  //7 / 210 = 0
    16'b00000111_11010011 : OUT <= 0;  //7 / 211 = 0
    16'b00000111_11010100 : OUT <= 0;  //7 / 212 = 0
    16'b00000111_11010101 : OUT <= 0;  //7 / 213 = 0
    16'b00000111_11010110 : OUT <= 0;  //7 / 214 = 0
    16'b00000111_11010111 : OUT <= 0;  //7 / 215 = 0
    16'b00000111_11011000 : OUT <= 0;  //7 / 216 = 0
    16'b00000111_11011001 : OUT <= 0;  //7 / 217 = 0
    16'b00000111_11011010 : OUT <= 0;  //7 / 218 = 0
    16'b00000111_11011011 : OUT <= 0;  //7 / 219 = 0
    16'b00000111_11011100 : OUT <= 0;  //7 / 220 = 0
    16'b00000111_11011101 : OUT <= 0;  //7 / 221 = 0
    16'b00000111_11011110 : OUT <= 0;  //7 / 222 = 0
    16'b00000111_11011111 : OUT <= 0;  //7 / 223 = 0
    16'b00000111_11100000 : OUT <= 0;  //7 / 224 = 0
    16'b00000111_11100001 : OUT <= 0;  //7 / 225 = 0
    16'b00000111_11100010 : OUT <= 0;  //7 / 226 = 0
    16'b00000111_11100011 : OUT <= 0;  //7 / 227 = 0
    16'b00000111_11100100 : OUT <= 0;  //7 / 228 = 0
    16'b00000111_11100101 : OUT <= 0;  //7 / 229 = 0
    16'b00000111_11100110 : OUT <= 0;  //7 / 230 = 0
    16'b00000111_11100111 : OUT <= 0;  //7 / 231 = 0
    16'b00000111_11101000 : OUT <= 0;  //7 / 232 = 0
    16'b00000111_11101001 : OUT <= 0;  //7 / 233 = 0
    16'b00000111_11101010 : OUT <= 0;  //7 / 234 = 0
    16'b00000111_11101011 : OUT <= 0;  //7 / 235 = 0
    16'b00000111_11101100 : OUT <= 0;  //7 / 236 = 0
    16'b00000111_11101101 : OUT <= 0;  //7 / 237 = 0
    16'b00000111_11101110 : OUT <= 0;  //7 / 238 = 0
    16'b00000111_11101111 : OUT <= 0;  //7 / 239 = 0
    16'b00000111_11110000 : OUT <= 0;  //7 / 240 = 0
    16'b00000111_11110001 : OUT <= 0;  //7 / 241 = 0
    16'b00000111_11110010 : OUT <= 0;  //7 / 242 = 0
    16'b00000111_11110011 : OUT <= 0;  //7 / 243 = 0
    16'b00000111_11110100 : OUT <= 0;  //7 / 244 = 0
    16'b00000111_11110101 : OUT <= 0;  //7 / 245 = 0
    16'b00000111_11110110 : OUT <= 0;  //7 / 246 = 0
    16'b00000111_11110111 : OUT <= 0;  //7 / 247 = 0
    16'b00000111_11111000 : OUT <= 0;  //7 / 248 = 0
    16'b00000111_11111001 : OUT <= 0;  //7 / 249 = 0
    16'b00000111_11111010 : OUT <= 0;  //7 / 250 = 0
    16'b00000111_11111011 : OUT <= 0;  //7 / 251 = 0
    16'b00000111_11111100 : OUT <= 0;  //7 / 252 = 0
    16'b00000111_11111101 : OUT <= 0;  //7 / 253 = 0
    16'b00000111_11111110 : OUT <= 0;  //7 / 254 = 0
    16'b00000111_11111111 : OUT <= 0;  //7 / 255 = 0
    16'b00001000_00000000 : OUT <= 0;  //8 / 0 = 0
    16'b00001000_00000001 : OUT <= 8;  //8 / 1 = 8
    16'b00001000_00000010 : OUT <= 4;  //8 / 2 = 4
    16'b00001000_00000011 : OUT <= 2;  //8 / 3 = 2
    16'b00001000_00000100 : OUT <= 2;  //8 / 4 = 2
    16'b00001000_00000101 : OUT <= 1;  //8 / 5 = 1
    16'b00001000_00000110 : OUT <= 1;  //8 / 6 = 1
    16'b00001000_00000111 : OUT <= 1;  //8 / 7 = 1
    16'b00001000_00001000 : OUT <= 1;  //8 / 8 = 1
    16'b00001000_00001001 : OUT <= 0;  //8 / 9 = 0
    16'b00001000_00001010 : OUT <= 0;  //8 / 10 = 0
    16'b00001000_00001011 : OUT <= 0;  //8 / 11 = 0
    16'b00001000_00001100 : OUT <= 0;  //8 / 12 = 0
    16'b00001000_00001101 : OUT <= 0;  //8 / 13 = 0
    16'b00001000_00001110 : OUT <= 0;  //8 / 14 = 0
    16'b00001000_00001111 : OUT <= 0;  //8 / 15 = 0
    16'b00001000_00010000 : OUT <= 0;  //8 / 16 = 0
    16'b00001000_00010001 : OUT <= 0;  //8 / 17 = 0
    16'b00001000_00010010 : OUT <= 0;  //8 / 18 = 0
    16'b00001000_00010011 : OUT <= 0;  //8 / 19 = 0
    16'b00001000_00010100 : OUT <= 0;  //8 / 20 = 0
    16'b00001000_00010101 : OUT <= 0;  //8 / 21 = 0
    16'b00001000_00010110 : OUT <= 0;  //8 / 22 = 0
    16'b00001000_00010111 : OUT <= 0;  //8 / 23 = 0
    16'b00001000_00011000 : OUT <= 0;  //8 / 24 = 0
    16'b00001000_00011001 : OUT <= 0;  //8 / 25 = 0
    16'b00001000_00011010 : OUT <= 0;  //8 / 26 = 0
    16'b00001000_00011011 : OUT <= 0;  //8 / 27 = 0
    16'b00001000_00011100 : OUT <= 0;  //8 / 28 = 0
    16'b00001000_00011101 : OUT <= 0;  //8 / 29 = 0
    16'b00001000_00011110 : OUT <= 0;  //8 / 30 = 0
    16'b00001000_00011111 : OUT <= 0;  //8 / 31 = 0
    16'b00001000_00100000 : OUT <= 0;  //8 / 32 = 0
    16'b00001000_00100001 : OUT <= 0;  //8 / 33 = 0
    16'b00001000_00100010 : OUT <= 0;  //8 / 34 = 0
    16'b00001000_00100011 : OUT <= 0;  //8 / 35 = 0
    16'b00001000_00100100 : OUT <= 0;  //8 / 36 = 0
    16'b00001000_00100101 : OUT <= 0;  //8 / 37 = 0
    16'b00001000_00100110 : OUT <= 0;  //8 / 38 = 0
    16'b00001000_00100111 : OUT <= 0;  //8 / 39 = 0
    16'b00001000_00101000 : OUT <= 0;  //8 / 40 = 0
    16'b00001000_00101001 : OUT <= 0;  //8 / 41 = 0
    16'b00001000_00101010 : OUT <= 0;  //8 / 42 = 0
    16'b00001000_00101011 : OUT <= 0;  //8 / 43 = 0
    16'b00001000_00101100 : OUT <= 0;  //8 / 44 = 0
    16'b00001000_00101101 : OUT <= 0;  //8 / 45 = 0
    16'b00001000_00101110 : OUT <= 0;  //8 / 46 = 0
    16'b00001000_00101111 : OUT <= 0;  //8 / 47 = 0
    16'b00001000_00110000 : OUT <= 0;  //8 / 48 = 0
    16'b00001000_00110001 : OUT <= 0;  //8 / 49 = 0
    16'b00001000_00110010 : OUT <= 0;  //8 / 50 = 0
    16'b00001000_00110011 : OUT <= 0;  //8 / 51 = 0
    16'b00001000_00110100 : OUT <= 0;  //8 / 52 = 0
    16'b00001000_00110101 : OUT <= 0;  //8 / 53 = 0
    16'b00001000_00110110 : OUT <= 0;  //8 / 54 = 0
    16'b00001000_00110111 : OUT <= 0;  //8 / 55 = 0
    16'b00001000_00111000 : OUT <= 0;  //8 / 56 = 0
    16'b00001000_00111001 : OUT <= 0;  //8 / 57 = 0
    16'b00001000_00111010 : OUT <= 0;  //8 / 58 = 0
    16'b00001000_00111011 : OUT <= 0;  //8 / 59 = 0
    16'b00001000_00111100 : OUT <= 0;  //8 / 60 = 0
    16'b00001000_00111101 : OUT <= 0;  //8 / 61 = 0
    16'b00001000_00111110 : OUT <= 0;  //8 / 62 = 0
    16'b00001000_00111111 : OUT <= 0;  //8 / 63 = 0
    16'b00001000_01000000 : OUT <= 0;  //8 / 64 = 0
    16'b00001000_01000001 : OUT <= 0;  //8 / 65 = 0
    16'b00001000_01000010 : OUT <= 0;  //8 / 66 = 0
    16'b00001000_01000011 : OUT <= 0;  //8 / 67 = 0
    16'b00001000_01000100 : OUT <= 0;  //8 / 68 = 0
    16'b00001000_01000101 : OUT <= 0;  //8 / 69 = 0
    16'b00001000_01000110 : OUT <= 0;  //8 / 70 = 0
    16'b00001000_01000111 : OUT <= 0;  //8 / 71 = 0
    16'b00001000_01001000 : OUT <= 0;  //8 / 72 = 0
    16'b00001000_01001001 : OUT <= 0;  //8 / 73 = 0
    16'b00001000_01001010 : OUT <= 0;  //8 / 74 = 0
    16'b00001000_01001011 : OUT <= 0;  //8 / 75 = 0
    16'b00001000_01001100 : OUT <= 0;  //8 / 76 = 0
    16'b00001000_01001101 : OUT <= 0;  //8 / 77 = 0
    16'b00001000_01001110 : OUT <= 0;  //8 / 78 = 0
    16'b00001000_01001111 : OUT <= 0;  //8 / 79 = 0
    16'b00001000_01010000 : OUT <= 0;  //8 / 80 = 0
    16'b00001000_01010001 : OUT <= 0;  //8 / 81 = 0
    16'b00001000_01010010 : OUT <= 0;  //8 / 82 = 0
    16'b00001000_01010011 : OUT <= 0;  //8 / 83 = 0
    16'b00001000_01010100 : OUT <= 0;  //8 / 84 = 0
    16'b00001000_01010101 : OUT <= 0;  //8 / 85 = 0
    16'b00001000_01010110 : OUT <= 0;  //8 / 86 = 0
    16'b00001000_01010111 : OUT <= 0;  //8 / 87 = 0
    16'b00001000_01011000 : OUT <= 0;  //8 / 88 = 0
    16'b00001000_01011001 : OUT <= 0;  //8 / 89 = 0
    16'b00001000_01011010 : OUT <= 0;  //8 / 90 = 0
    16'b00001000_01011011 : OUT <= 0;  //8 / 91 = 0
    16'b00001000_01011100 : OUT <= 0;  //8 / 92 = 0
    16'b00001000_01011101 : OUT <= 0;  //8 / 93 = 0
    16'b00001000_01011110 : OUT <= 0;  //8 / 94 = 0
    16'b00001000_01011111 : OUT <= 0;  //8 / 95 = 0
    16'b00001000_01100000 : OUT <= 0;  //8 / 96 = 0
    16'b00001000_01100001 : OUT <= 0;  //8 / 97 = 0
    16'b00001000_01100010 : OUT <= 0;  //8 / 98 = 0
    16'b00001000_01100011 : OUT <= 0;  //8 / 99 = 0
    16'b00001000_01100100 : OUT <= 0;  //8 / 100 = 0
    16'b00001000_01100101 : OUT <= 0;  //8 / 101 = 0
    16'b00001000_01100110 : OUT <= 0;  //8 / 102 = 0
    16'b00001000_01100111 : OUT <= 0;  //8 / 103 = 0
    16'b00001000_01101000 : OUT <= 0;  //8 / 104 = 0
    16'b00001000_01101001 : OUT <= 0;  //8 / 105 = 0
    16'b00001000_01101010 : OUT <= 0;  //8 / 106 = 0
    16'b00001000_01101011 : OUT <= 0;  //8 / 107 = 0
    16'b00001000_01101100 : OUT <= 0;  //8 / 108 = 0
    16'b00001000_01101101 : OUT <= 0;  //8 / 109 = 0
    16'b00001000_01101110 : OUT <= 0;  //8 / 110 = 0
    16'b00001000_01101111 : OUT <= 0;  //8 / 111 = 0
    16'b00001000_01110000 : OUT <= 0;  //8 / 112 = 0
    16'b00001000_01110001 : OUT <= 0;  //8 / 113 = 0
    16'b00001000_01110010 : OUT <= 0;  //8 / 114 = 0
    16'b00001000_01110011 : OUT <= 0;  //8 / 115 = 0
    16'b00001000_01110100 : OUT <= 0;  //8 / 116 = 0
    16'b00001000_01110101 : OUT <= 0;  //8 / 117 = 0
    16'b00001000_01110110 : OUT <= 0;  //8 / 118 = 0
    16'b00001000_01110111 : OUT <= 0;  //8 / 119 = 0
    16'b00001000_01111000 : OUT <= 0;  //8 / 120 = 0
    16'b00001000_01111001 : OUT <= 0;  //8 / 121 = 0
    16'b00001000_01111010 : OUT <= 0;  //8 / 122 = 0
    16'b00001000_01111011 : OUT <= 0;  //8 / 123 = 0
    16'b00001000_01111100 : OUT <= 0;  //8 / 124 = 0
    16'b00001000_01111101 : OUT <= 0;  //8 / 125 = 0
    16'b00001000_01111110 : OUT <= 0;  //8 / 126 = 0
    16'b00001000_01111111 : OUT <= 0;  //8 / 127 = 0
    16'b00001000_10000000 : OUT <= 0;  //8 / 128 = 0
    16'b00001000_10000001 : OUT <= 0;  //8 / 129 = 0
    16'b00001000_10000010 : OUT <= 0;  //8 / 130 = 0
    16'b00001000_10000011 : OUT <= 0;  //8 / 131 = 0
    16'b00001000_10000100 : OUT <= 0;  //8 / 132 = 0
    16'b00001000_10000101 : OUT <= 0;  //8 / 133 = 0
    16'b00001000_10000110 : OUT <= 0;  //8 / 134 = 0
    16'b00001000_10000111 : OUT <= 0;  //8 / 135 = 0
    16'b00001000_10001000 : OUT <= 0;  //8 / 136 = 0
    16'b00001000_10001001 : OUT <= 0;  //8 / 137 = 0
    16'b00001000_10001010 : OUT <= 0;  //8 / 138 = 0
    16'b00001000_10001011 : OUT <= 0;  //8 / 139 = 0
    16'b00001000_10001100 : OUT <= 0;  //8 / 140 = 0
    16'b00001000_10001101 : OUT <= 0;  //8 / 141 = 0
    16'b00001000_10001110 : OUT <= 0;  //8 / 142 = 0
    16'b00001000_10001111 : OUT <= 0;  //8 / 143 = 0
    16'b00001000_10010000 : OUT <= 0;  //8 / 144 = 0
    16'b00001000_10010001 : OUT <= 0;  //8 / 145 = 0
    16'b00001000_10010010 : OUT <= 0;  //8 / 146 = 0
    16'b00001000_10010011 : OUT <= 0;  //8 / 147 = 0
    16'b00001000_10010100 : OUT <= 0;  //8 / 148 = 0
    16'b00001000_10010101 : OUT <= 0;  //8 / 149 = 0
    16'b00001000_10010110 : OUT <= 0;  //8 / 150 = 0
    16'b00001000_10010111 : OUT <= 0;  //8 / 151 = 0
    16'b00001000_10011000 : OUT <= 0;  //8 / 152 = 0
    16'b00001000_10011001 : OUT <= 0;  //8 / 153 = 0
    16'b00001000_10011010 : OUT <= 0;  //8 / 154 = 0
    16'b00001000_10011011 : OUT <= 0;  //8 / 155 = 0
    16'b00001000_10011100 : OUT <= 0;  //8 / 156 = 0
    16'b00001000_10011101 : OUT <= 0;  //8 / 157 = 0
    16'b00001000_10011110 : OUT <= 0;  //8 / 158 = 0
    16'b00001000_10011111 : OUT <= 0;  //8 / 159 = 0
    16'b00001000_10100000 : OUT <= 0;  //8 / 160 = 0
    16'b00001000_10100001 : OUT <= 0;  //8 / 161 = 0
    16'b00001000_10100010 : OUT <= 0;  //8 / 162 = 0
    16'b00001000_10100011 : OUT <= 0;  //8 / 163 = 0
    16'b00001000_10100100 : OUT <= 0;  //8 / 164 = 0
    16'b00001000_10100101 : OUT <= 0;  //8 / 165 = 0
    16'b00001000_10100110 : OUT <= 0;  //8 / 166 = 0
    16'b00001000_10100111 : OUT <= 0;  //8 / 167 = 0
    16'b00001000_10101000 : OUT <= 0;  //8 / 168 = 0
    16'b00001000_10101001 : OUT <= 0;  //8 / 169 = 0
    16'b00001000_10101010 : OUT <= 0;  //8 / 170 = 0
    16'b00001000_10101011 : OUT <= 0;  //8 / 171 = 0
    16'b00001000_10101100 : OUT <= 0;  //8 / 172 = 0
    16'b00001000_10101101 : OUT <= 0;  //8 / 173 = 0
    16'b00001000_10101110 : OUT <= 0;  //8 / 174 = 0
    16'b00001000_10101111 : OUT <= 0;  //8 / 175 = 0
    16'b00001000_10110000 : OUT <= 0;  //8 / 176 = 0
    16'b00001000_10110001 : OUT <= 0;  //8 / 177 = 0
    16'b00001000_10110010 : OUT <= 0;  //8 / 178 = 0
    16'b00001000_10110011 : OUT <= 0;  //8 / 179 = 0
    16'b00001000_10110100 : OUT <= 0;  //8 / 180 = 0
    16'b00001000_10110101 : OUT <= 0;  //8 / 181 = 0
    16'b00001000_10110110 : OUT <= 0;  //8 / 182 = 0
    16'b00001000_10110111 : OUT <= 0;  //8 / 183 = 0
    16'b00001000_10111000 : OUT <= 0;  //8 / 184 = 0
    16'b00001000_10111001 : OUT <= 0;  //8 / 185 = 0
    16'b00001000_10111010 : OUT <= 0;  //8 / 186 = 0
    16'b00001000_10111011 : OUT <= 0;  //8 / 187 = 0
    16'b00001000_10111100 : OUT <= 0;  //8 / 188 = 0
    16'b00001000_10111101 : OUT <= 0;  //8 / 189 = 0
    16'b00001000_10111110 : OUT <= 0;  //8 / 190 = 0
    16'b00001000_10111111 : OUT <= 0;  //8 / 191 = 0
    16'b00001000_11000000 : OUT <= 0;  //8 / 192 = 0
    16'b00001000_11000001 : OUT <= 0;  //8 / 193 = 0
    16'b00001000_11000010 : OUT <= 0;  //8 / 194 = 0
    16'b00001000_11000011 : OUT <= 0;  //8 / 195 = 0
    16'b00001000_11000100 : OUT <= 0;  //8 / 196 = 0
    16'b00001000_11000101 : OUT <= 0;  //8 / 197 = 0
    16'b00001000_11000110 : OUT <= 0;  //8 / 198 = 0
    16'b00001000_11000111 : OUT <= 0;  //8 / 199 = 0
    16'b00001000_11001000 : OUT <= 0;  //8 / 200 = 0
    16'b00001000_11001001 : OUT <= 0;  //8 / 201 = 0
    16'b00001000_11001010 : OUT <= 0;  //8 / 202 = 0
    16'b00001000_11001011 : OUT <= 0;  //8 / 203 = 0
    16'b00001000_11001100 : OUT <= 0;  //8 / 204 = 0
    16'b00001000_11001101 : OUT <= 0;  //8 / 205 = 0
    16'b00001000_11001110 : OUT <= 0;  //8 / 206 = 0
    16'b00001000_11001111 : OUT <= 0;  //8 / 207 = 0
    16'b00001000_11010000 : OUT <= 0;  //8 / 208 = 0
    16'b00001000_11010001 : OUT <= 0;  //8 / 209 = 0
    16'b00001000_11010010 : OUT <= 0;  //8 / 210 = 0
    16'b00001000_11010011 : OUT <= 0;  //8 / 211 = 0
    16'b00001000_11010100 : OUT <= 0;  //8 / 212 = 0
    16'b00001000_11010101 : OUT <= 0;  //8 / 213 = 0
    16'b00001000_11010110 : OUT <= 0;  //8 / 214 = 0
    16'b00001000_11010111 : OUT <= 0;  //8 / 215 = 0
    16'b00001000_11011000 : OUT <= 0;  //8 / 216 = 0
    16'b00001000_11011001 : OUT <= 0;  //8 / 217 = 0
    16'b00001000_11011010 : OUT <= 0;  //8 / 218 = 0
    16'b00001000_11011011 : OUT <= 0;  //8 / 219 = 0
    16'b00001000_11011100 : OUT <= 0;  //8 / 220 = 0
    16'b00001000_11011101 : OUT <= 0;  //8 / 221 = 0
    16'b00001000_11011110 : OUT <= 0;  //8 / 222 = 0
    16'b00001000_11011111 : OUT <= 0;  //8 / 223 = 0
    16'b00001000_11100000 : OUT <= 0;  //8 / 224 = 0
    16'b00001000_11100001 : OUT <= 0;  //8 / 225 = 0
    16'b00001000_11100010 : OUT <= 0;  //8 / 226 = 0
    16'b00001000_11100011 : OUT <= 0;  //8 / 227 = 0
    16'b00001000_11100100 : OUT <= 0;  //8 / 228 = 0
    16'b00001000_11100101 : OUT <= 0;  //8 / 229 = 0
    16'b00001000_11100110 : OUT <= 0;  //8 / 230 = 0
    16'b00001000_11100111 : OUT <= 0;  //8 / 231 = 0
    16'b00001000_11101000 : OUT <= 0;  //8 / 232 = 0
    16'b00001000_11101001 : OUT <= 0;  //8 / 233 = 0
    16'b00001000_11101010 : OUT <= 0;  //8 / 234 = 0
    16'b00001000_11101011 : OUT <= 0;  //8 / 235 = 0
    16'b00001000_11101100 : OUT <= 0;  //8 / 236 = 0
    16'b00001000_11101101 : OUT <= 0;  //8 / 237 = 0
    16'b00001000_11101110 : OUT <= 0;  //8 / 238 = 0
    16'b00001000_11101111 : OUT <= 0;  //8 / 239 = 0
    16'b00001000_11110000 : OUT <= 0;  //8 / 240 = 0
    16'b00001000_11110001 : OUT <= 0;  //8 / 241 = 0
    16'b00001000_11110010 : OUT <= 0;  //8 / 242 = 0
    16'b00001000_11110011 : OUT <= 0;  //8 / 243 = 0
    16'b00001000_11110100 : OUT <= 0;  //8 / 244 = 0
    16'b00001000_11110101 : OUT <= 0;  //8 / 245 = 0
    16'b00001000_11110110 : OUT <= 0;  //8 / 246 = 0
    16'b00001000_11110111 : OUT <= 0;  //8 / 247 = 0
    16'b00001000_11111000 : OUT <= 0;  //8 / 248 = 0
    16'b00001000_11111001 : OUT <= 0;  //8 / 249 = 0
    16'b00001000_11111010 : OUT <= 0;  //8 / 250 = 0
    16'b00001000_11111011 : OUT <= 0;  //8 / 251 = 0
    16'b00001000_11111100 : OUT <= 0;  //8 / 252 = 0
    16'b00001000_11111101 : OUT <= 0;  //8 / 253 = 0
    16'b00001000_11111110 : OUT <= 0;  //8 / 254 = 0
    16'b00001000_11111111 : OUT <= 0;  //8 / 255 = 0
    16'b00001001_00000000 : OUT <= 0;  //9 / 0 = 0
    16'b00001001_00000001 : OUT <= 9;  //9 / 1 = 9
    16'b00001001_00000010 : OUT <= 4;  //9 / 2 = 4
    16'b00001001_00000011 : OUT <= 3;  //9 / 3 = 3
    16'b00001001_00000100 : OUT <= 2;  //9 / 4 = 2
    16'b00001001_00000101 : OUT <= 1;  //9 / 5 = 1
    16'b00001001_00000110 : OUT <= 1;  //9 / 6 = 1
    16'b00001001_00000111 : OUT <= 1;  //9 / 7 = 1
    16'b00001001_00001000 : OUT <= 1;  //9 / 8 = 1
    16'b00001001_00001001 : OUT <= 1;  //9 / 9 = 1
    16'b00001001_00001010 : OUT <= 0;  //9 / 10 = 0
    16'b00001001_00001011 : OUT <= 0;  //9 / 11 = 0
    16'b00001001_00001100 : OUT <= 0;  //9 / 12 = 0
    16'b00001001_00001101 : OUT <= 0;  //9 / 13 = 0
    16'b00001001_00001110 : OUT <= 0;  //9 / 14 = 0
    16'b00001001_00001111 : OUT <= 0;  //9 / 15 = 0
    16'b00001001_00010000 : OUT <= 0;  //9 / 16 = 0
    16'b00001001_00010001 : OUT <= 0;  //9 / 17 = 0
    16'b00001001_00010010 : OUT <= 0;  //9 / 18 = 0
    16'b00001001_00010011 : OUT <= 0;  //9 / 19 = 0
    16'b00001001_00010100 : OUT <= 0;  //9 / 20 = 0
    16'b00001001_00010101 : OUT <= 0;  //9 / 21 = 0
    16'b00001001_00010110 : OUT <= 0;  //9 / 22 = 0
    16'b00001001_00010111 : OUT <= 0;  //9 / 23 = 0
    16'b00001001_00011000 : OUT <= 0;  //9 / 24 = 0
    16'b00001001_00011001 : OUT <= 0;  //9 / 25 = 0
    16'b00001001_00011010 : OUT <= 0;  //9 / 26 = 0
    16'b00001001_00011011 : OUT <= 0;  //9 / 27 = 0
    16'b00001001_00011100 : OUT <= 0;  //9 / 28 = 0
    16'b00001001_00011101 : OUT <= 0;  //9 / 29 = 0
    16'b00001001_00011110 : OUT <= 0;  //9 / 30 = 0
    16'b00001001_00011111 : OUT <= 0;  //9 / 31 = 0
    16'b00001001_00100000 : OUT <= 0;  //9 / 32 = 0
    16'b00001001_00100001 : OUT <= 0;  //9 / 33 = 0
    16'b00001001_00100010 : OUT <= 0;  //9 / 34 = 0
    16'b00001001_00100011 : OUT <= 0;  //9 / 35 = 0
    16'b00001001_00100100 : OUT <= 0;  //9 / 36 = 0
    16'b00001001_00100101 : OUT <= 0;  //9 / 37 = 0
    16'b00001001_00100110 : OUT <= 0;  //9 / 38 = 0
    16'b00001001_00100111 : OUT <= 0;  //9 / 39 = 0
    16'b00001001_00101000 : OUT <= 0;  //9 / 40 = 0
    16'b00001001_00101001 : OUT <= 0;  //9 / 41 = 0
    16'b00001001_00101010 : OUT <= 0;  //9 / 42 = 0
    16'b00001001_00101011 : OUT <= 0;  //9 / 43 = 0
    16'b00001001_00101100 : OUT <= 0;  //9 / 44 = 0
    16'b00001001_00101101 : OUT <= 0;  //9 / 45 = 0
    16'b00001001_00101110 : OUT <= 0;  //9 / 46 = 0
    16'b00001001_00101111 : OUT <= 0;  //9 / 47 = 0
    16'b00001001_00110000 : OUT <= 0;  //9 / 48 = 0
    16'b00001001_00110001 : OUT <= 0;  //9 / 49 = 0
    16'b00001001_00110010 : OUT <= 0;  //9 / 50 = 0
    16'b00001001_00110011 : OUT <= 0;  //9 / 51 = 0
    16'b00001001_00110100 : OUT <= 0;  //9 / 52 = 0
    16'b00001001_00110101 : OUT <= 0;  //9 / 53 = 0
    16'b00001001_00110110 : OUT <= 0;  //9 / 54 = 0
    16'b00001001_00110111 : OUT <= 0;  //9 / 55 = 0
    16'b00001001_00111000 : OUT <= 0;  //9 / 56 = 0
    16'b00001001_00111001 : OUT <= 0;  //9 / 57 = 0
    16'b00001001_00111010 : OUT <= 0;  //9 / 58 = 0
    16'b00001001_00111011 : OUT <= 0;  //9 / 59 = 0
    16'b00001001_00111100 : OUT <= 0;  //9 / 60 = 0
    16'b00001001_00111101 : OUT <= 0;  //9 / 61 = 0
    16'b00001001_00111110 : OUT <= 0;  //9 / 62 = 0
    16'b00001001_00111111 : OUT <= 0;  //9 / 63 = 0
    16'b00001001_01000000 : OUT <= 0;  //9 / 64 = 0
    16'b00001001_01000001 : OUT <= 0;  //9 / 65 = 0
    16'b00001001_01000010 : OUT <= 0;  //9 / 66 = 0
    16'b00001001_01000011 : OUT <= 0;  //9 / 67 = 0
    16'b00001001_01000100 : OUT <= 0;  //9 / 68 = 0
    16'b00001001_01000101 : OUT <= 0;  //9 / 69 = 0
    16'b00001001_01000110 : OUT <= 0;  //9 / 70 = 0
    16'b00001001_01000111 : OUT <= 0;  //9 / 71 = 0
    16'b00001001_01001000 : OUT <= 0;  //9 / 72 = 0
    16'b00001001_01001001 : OUT <= 0;  //9 / 73 = 0
    16'b00001001_01001010 : OUT <= 0;  //9 / 74 = 0
    16'b00001001_01001011 : OUT <= 0;  //9 / 75 = 0
    16'b00001001_01001100 : OUT <= 0;  //9 / 76 = 0
    16'b00001001_01001101 : OUT <= 0;  //9 / 77 = 0
    16'b00001001_01001110 : OUT <= 0;  //9 / 78 = 0
    16'b00001001_01001111 : OUT <= 0;  //9 / 79 = 0
    16'b00001001_01010000 : OUT <= 0;  //9 / 80 = 0
    16'b00001001_01010001 : OUT <= 0;  //9 / 81 = 0
    16'b00001001_01010010 : OUT <= 0;  //9 / 82 = 0
    16'b00001001_01010011 : OUT <= 0;  //9 / 83 = 0
    16'b00001001_01010100 : OUT <= 0;  //9 / 84 = 0
    16'b00001001_01010101 : OUT <= 0;  //9 / 85 = 0
    16'b00001001_01010110 : OUT <= 0;  //9 / 86 = 0
    16'b00001001_01010111 : OUT <= 0;  //9 / 87 = 0
    16'b00001001_01011000 : OUT <= 0;  //9 / 88 = 0
    16'b00001001_01011001 : OUT <= 0;  //9 / 89 = 0
    16'b00001001_01011010 : OUT <= 0;  //9 / 90 = 0
    16'b00001001_01011011 : OUT <= 0;  //9 / 91 = 0
    16'b00001001_01011100 : OUT <= 0;  //9 / 92 = 0
    16'b00001001_01011101 : OUT <= 0;  //9 / 93 = 0
    16'b00001001_01011110 : OUT <= 0;  //9 / 94 = 0
    16'b00001001_01011111 : OUT <= 0;  //9 / 95 = 0
    16'b00001001_01100000 : OUT <= 0;  //9 / 96 = 0
    16'b00001001_01100001 : OUT <= 0;  //9 / 97 = 0
    16'b00001001_01100010 : OUT <= 0;  //9 / 98 = 0
    16'b00001001_01100011 : OUT <= 0;  //9 / 99 = 0
    16'b00001001_01100100 : OUT <= 0;  //9 / 100 = 0
    16'b00001001_01100101 : OUT <= 0;  //9 / 101 = 0
    16'b00001001_01100110 : OUT <= 0;  //9 / 102 = 0
    16'b00001001_01100111 : OUT <= 0;  //9 / 103 = 0
    16'b00001001_01101000 : OUT <= 0;  //9 / 104 = 0
    16'b00001001_01101001 : OUT <= 0;  //9 / 105 = 0
    16'b00001001_01101010 : OUT <= 0;  //9 / 106 = 0
    16'b00001001_01101011 : OUT <= 0;  //9 / 107 = 0
    16'b00001001_01101100 : OUT <= 0;  //9 / 108 = 0
    16'b00001001_01101101 : OUT <= 0;  //9 / 109 = 0
    16'b00001001_01101110 : OUT <= 0;  //9 / 110 = 0
    16'b00001001_01101111 : OUT <= 0;  //9 / 111 = 0
    16'b00001001_01110000 : OUT <= 0;  //9 / 112 = 0
    16'b00001001_01110001 : OUT <= 0;  //9 / 113 = 0
    16'b00001001_01110010 : OUT <= 0;  //9 / 114 = 0
    16'b00001001_01110011 : OUT <= 0;  //9 / 115 = 0
    16'b00001001_01110100 : OUT <= 0;  //9 / 116 = 0
    16'b00001001_01110101 : OUT <= 0;  //9 / 117 = 0
    16'b00001001_01110110 : OUT <= 0;  //9 / 118 = 0
    16'b00001001_01110111 : OUT <= 0;  //9 / 119 = 0
    16'b00001001_01111000 : OUT <= 0;  //9 / 120 = 0
    16'b00001001_01111001 : OUT <= 0;  //9 / 121 = 0
    16'b00001001_01111010 : OUT <= 0;  //9 / 122 = 0
    16'b00001001_01111011 : OUT <= 0;  //9 / 123 = 0
    16'b00001001_01111100 : OUT <= 0;  //9 / 124 = 0
    16'b00001001_01111101 : OUT <= 0;  //9 / 125 = 0
    16'b00001001_01111110 : OUT <= 0;  //9 / 126 = 0
    16'b00001001_01111111 : OUT <= 0;  //9 / 127 = 0
    16'b00001001_10000000 : OUT <= 0;  //9 / 128 = 0
    16'b00001001_10000001 : OUT <= 0;  //9 / 129 = 0
    16'b00001001_10000010 : OUT <= 0;  //9 / 130 = 0
    16'b00001001_10000011 : OUT <= 0;  //9 / 131 = 0
    16'b00001001_10000100 : OUT <= 0;  //9 / 132 = 0
    16'b00001001_10000101 : OUT <= 0;  //9 / 133 = 0
    16'b00001001_10000110 : OUT <= 0;  //9 / 134 = 0
    16'b00001001_10000111 : OUT <= 0;  //9 / 135 = 0
    16'b00001001_10001000 : OUT <= 0;  //9 / 136 = 0
    16'b00001001_10001001 : OUT <= 0;  //9 / 137 = 0
    16'b00001001_10001010 : OUT <= 0;  //9 / 138 = 0
    16'b00001001_10001011 : OUT <= 0;  //9 / 139 = 0
    16'b00001001_10001100 : OUT <= 0;  //9 / 140 = 0
    16'b00001001_10001101 : OUT <= 0;  //9 / 141 = 0
    16'b00001001_10001110 : OUT <= 0;  //9 / 142 = 0
    16'b00001001_10001111 : OUT <= 0;  //9 / 143 = 0
    16'b00001001_10010000 : OUT <= 0;  //9 / 144 = 0
    16'b00001001_10010001 : OUT <= 0;  //9 / 145 = 0
    16'b00001001_10010010 : OUT <= 0;  //9 / 146 = 0
    16'b00001001_10010011 : OUT <= 0;  //9 / 147 = 0
    16'b00001001_10010100 : OUT <= 0;  //9 / 148 = 0
    16'b00001001_10010101 : OUT <= 0;  //9 / 149 = 0
    16'b00001001_10010110 : OUT <= 0;  //9 / 150 = 0
    16'b00001001_10010111 : OUT <= 0;  //9 / 151 = 0
    16'b00001001_10011000 : OUT <= 0;  //9 / 152 = 0
    16'b00001001_10011001 : OUT <= 0;  //9 / 153 = 0
    16'b00001001_10011010 : OUT <= 0;  //9 / 154 = 0
    16'b00001001_10011011 : OUT <= 0;  //9 / 155 = 0
    16'b00001001_10011100 : OUT <= 0;  //9 / 156 = 0
    16'b00001001_10011101 : OUT <= 0;  //9 / 157 = 0
    16'b00001001_10011110 : OUT <= 0;  //9 / 158 = 0
    16'b00001001_10011111 : OUT <= 0;  //9 / 159 = 0
    16'b00001001_10100000 : OUT <= 0;  //9 / 160 = 0
    16'b00001001_10100001 : OUT <= 0;  //9 / 161 = 0
    16'b00001001_10100010 : OUT <= 0;  //9 / 162 = 0
    16'b00001001_10100011 : OUT <= 0;  //9 / 163 = 0
    16'b00001001_10100100 : OUT <= 0;  //9 / 164 = 0
    16'b00001001_10100101 : OUT <= 0;  //9 / 165 = 0
    16'b00001001_10100110 : OUT <= 0;  //9 / 166 = 0
    16'b00001001_10100111 : OUT <= 0;  //9 / 167 = 0
    16'b00001001_10101000 : OUT <= 0;  //9 / 168 = 0
    16'b00001001_10101001 : OUT <= 0;  //9 / 169 = 0
    16'b00001001_10101010 : OUT <= 0;  //9 / 170 = 0
    16'b00001001_10101011 : OUT <= 0;  //9 / 171 = 0
    16'b00001001_10101100 : OUT <= 0;  //9 / 172 = 0
    16'b00001001_10101101 : OUT <= 0;  //9 / 173 = 0
    16'b00001001_10101110 : OUT <= 0;  //9 / 174 = 0
    16'b00001001_10101111 : OUT <= 0;  //9 / 175 = 0
    16'b00001001_10110000 : OUT <= 0;  //9 / 176 = 0
    16'b00001001_10110001 : OUT <= 0;  //9 / 177 = 0
    16'b00001001_10110010 : OUT <= 0;  //9 / 178 = 0
    16'b00001001_10110011 : OUT <= 0;  //9 / 179 = 0
    16'b00001001_10110100 : OUT <= 0;  //9 / 180 = 0
    16'b00001001_10110101 : OUT <= 0;  //9 / 181 = 0
    16'b00001001_10110110 : OUT <= 0;  //9 / 182 = 0
    16'b00001001_10110111 : OUT <= 0;  //9 / 183 = 0
    16'b00001001_10111000 : OUT <= 0;  //9 / 184 = 0
    16'b00001001_10111001 : OUT <= 0;  //9 / 185 = 0
    16'b00001001_10111010 : OUT <= 0;  //9 / 186 = 0
    16'b00001001_10111011 : OUT <= 0;  //9 / 187 = 0
    16'b00001001_10111100 : OUT <= 0;  //9 / 188 = 0
    16'b00001001_10111101 : OUT <= 0;  //9 / 189 = 0
    16'b00001001_10111110 : OUT <= 0;  //9 / 190 = 0
    16'b00001001_10111111 : OUT <= 0;  //9 / 191 = 0
    16'b00001001_11000000 : OUT <= 0;  //9 / 192 = 0
    16'b00001001_11000001 : OUT <= 0;  //9 / 193 = 0
    16'b00001001_11000010 : OUT <= 0;  //9 / 194 = 0
    16'b00001001_11000011 : OUT <= 0;  //9 / 195 = 0
    16'b00001001_11000100 : OUT <= 0;  //9 / 196 = 0
    16'b00001001_11000101 : OUT <= 0;  //9 / 197 = 0
    16'b00001001_11000110 : OUT <= 0;  //9 / 198 = 0
    16'b00001001_11000111 : OUT <= 0;  //9 / 199 = 0
    16'b00001001_11001000 : OUT <= 0;  //9 / 200 = 0
    16'b00001001_11001001 : OUT <= 0;  //9 / 201 = 0
    16'b00001001_11001010 : OUT <= 0;  //9 / 202 = 0
    16'b00001001_11001011 : OUT <= 0;  //9 / 203 = 0
    16'b00001001_11001100 : OUT <= 0;  //9 / 204 = 0
    16'b00001001_11001101 : OUT <= 0;  //9 / 205 = 0
    16'b00001001_11001110 : OUT <= 0;  //9 / 206 = 0
    16'b00001001_11001111 : OUT <= 0;  //9 / 207 = 0
    16'b00001001_11010000 : OUT <= 0;  //9 / 208 = 0
    16'b00001001_11010001 : OUT <= 0;  //9 / 209 = 0
    16'b00001001_11010010 : OUT <= 0;  //9 / 210 = 0
    16'b00001001_11010011 : OUT <= 0;  //9 / 211 = 0
    16'b00001001_11010100 : OUT <= 0;  //9 / 212 = 0
    16'b00001001_11010101 : OUT <= 0;  //9 / 213 = 0
    16'b00001001_11010110 : OUT <= 0;  //9 / 214 = 0
    16'b00001001_11010111 : OUT <= 0;  //9 / 215 = 0
    16'b00001001_11011000 : OUT <= 0;  //9 / 216 = 0
    16'b00001001_11011001 : OUT <= 0;  //9 / 217 = 0
    16'b00001001_11011010 : OUT <= 0;  //9 / 218 = 0
    16'b00001001_11011011 : OUT <= 0;  //9 / 219 = 0
    16'b00001001_11011100 : OUT <= 0;  //9 / 220 = 0
    16'b00001001_11011101 : OUT <= 0;  //9 / 221 = 0
    16'b00001001_11011110 : OUT <= 0;  //9 / 222 = 0
    16'b00001001_11011111 : OUT <= 0;  //9 / 223 = 0
    16'b00001001_11100000 : OUT <= 0;  //9 / 224 = 0
    16'b00001001_11100001 : OUT <= 0;  //9 / 225 = 0
    16'b00001001_11100010 : OUT <= 0;  //9 / 226 = 0
    16'b00001001_11100011 : OUT <= 0;  //9 / 227 = 0
    16'b00001001_11100100 : OUT <= 0;  //9 / 228 = 0
    16'b00001001_11100101 : OUT <= 0;  //9 / 229 = 0
    16'b00001001_11100110 : OUT <= 0;  //9 / 230 = 0
    16'b00001001_11100111 : OUT <= 0;  //9 / 231 = 0
    16'b00001001_11101000 : OUT <= 0;  //9 / 232 = 0
    16'b00001001_11101001 : OUT <= 0;  //9 / 233 = 0
    16'b00001001_11101010 : OUT <= 0;  //9 / 234 = 0
    16'b00001001_11101011 : OUT <= 0;  //9 / 235 = 0
    16'b00001001_11101100 : OUT <= 0;  //9 / 236 = 0
    16'b00001001_11101101 : OUT <= 0;  //9 / 237 = 0
    16'b00001001_11101110 : OUT <= 0;  //9 / 238 = 0
    16'b00001001_11101111 : OUT <= 0;  //9 / 239 = 0
    16'b00001001_11110000 : OUT <= 0;  //9 / 240 = 0
    16'b00001001_11110001 : OUT <= 0;  //9 / 241 = 0
    16'b00001001_11110010 : OUT <= 0;  //9 / 242 = 0
    16'b00001001_11110011 : OUT <= 0;  //9 / 243 = 0
    16'b00001001_11110100 : OUT <= 0;  //9 / 244 = 0
    16'b00001001_11110101 : OUT <= 0;  //9 / 245 = 0
    16'b00001001_11110110 : OUT <= 0;  //9 / 246 = 0
    16'b00001001_11110111 : OUT <= 0;  //9 / 247 = 0
    16'b00001001_11111000 : OUT <= 0;  //9 / 248 = 0
    16'b00001001_11111001 : OUT <= 0;  //9 / 249 = 0
    16'b00001001_11111010 : OUT <= 0;  //9 / 250 = 0
    16'b00001001_11111011 : OUT <= 0;  //9 / 251 = 0
    16'b00001001_11111100 : OUT <= 0;  //9 / 252 = 0
    16'b00001001_11111101 : OUT <= 0;  //9 / 253 = 0
    16'b00001001_11111110 : OUT <= 0;  //9 / 254 = 0
    16'b00001001_11111111 : OUT <= 0;  //9 / 255 = 0
    16'b00001010_00000000 : OUT <= 0;  //10 / 0 = 0
    16'b00001010_00000001 : OUT <= 10;  //10 / 1 = 10
    16'b00001010_00000010 : OUT <= 5;  //10 / 2 = 5
    16'b00001010_00000011 : OUT <= 3;  //10 / 3 = 3
    16'b00001010_00000100 : OUT <= 2;  //10 / 4 = 2
    16'b00001010_00000101 : OUT <= 2;  //10 / 5 = 2
    16'b00001010_00000110 : OUT <= 1;  //10 / 6 = 1
    16'b00001010_00000111 : OUT <= 1;  //10 / 7 = 1
    16'b00001010_00001000 : OUT <= 1;  //10 / 8 = 1
    16'b00001010_00001001 : OUT <= 1;  //10 / 9 = 1
    16'b00001010_00001010 : OUT <= 1;  //10 / 10 = 1
    16'b00001010_00001011 : OUT <= 0;  //10 / 11 = 0
    16'b00001010_00001100 : OUT <= 0;  //10 / 12 = 0
    16'b00001010_00001101 : OUT <= 0;  //10 / 13 = 0
    16'b00001010_00001110 : OUT <= 0;  //10 / 14 = 0
    16'b00001010_00001111 : OUT <= 0;  //10 / 15 = 0
    16'b00001010_00010000 : OUT <= 0;  //10 / 16 = 0
    16'b00001010_00010001 : OUT <= 0;  //10 / 17 = 0
    16'b00001010_00010010 : OUT <= 0;  //10 / 18 = 0
    16'b00001010_00010011 : OUT <= 0;  //10 / 19 = 0
    16'b00001010_00010100 : OUT <= 0;  //10 / 20 = 0
    16'b00001010_00010101 : OUT <= 0;  //10 / 21 = 0
    16'b00001010_00010110 : OUT <= 0;  //10 / 22 = 0
    16'b00001010_00010111 : OUT <= 0;  //10 / 23 = 0
    16'b00001010_00011000 : OUT <= 0;  //10 / 24 = 0
    16'b00001010_00011001 : OUT <= 0;  //10 / 25 = 0
    16'b00001010_00011010 : OUT <= 0;  //10 / 26 = 0
    16'b00001010_00011011 : OUT <= 0;  //10 / 27 = 0
    16'b00001010_00011100 : OUT <= 0;  //10 / 28 = 0
    16'b00001010_00011101 : OUT <= 0;  //10 / 29 = 0
    16'b00001010_00011110 : OUT <= 0;  //10 / 30 = 0
    16'b00001010_00011111 : OUT <= 0;  //10 / 31 = 0
    16'b00001010_00100000 : OUT <= 0;  //10 / 32 = 0
    16'b00001010_00100001 : OUT <= 0;  //10 / 33 = 0
    16'b00001010_00100010 : OUT <= 0;  //10 / 34 = 0
    16'b00001010_00100011 : OUT <= 0;  //10 / 35 = 0
    16'b00001010_00100100 : OUT <= 0;  //10 / 36 = 0
    16'b00001010_00100101 : OUT <= 0;  //10 / 37 = 0
    16'b00001010_00100110 : OUT <= 0;  //10 / 38 = 0
    16'b00001010_00100111 : OUT <= 0;  //10 / 39 = 0
    16'b00001010_00101000 : OUT <= 0;  //10 / 40 = 0
    16'b00001010_00101001 : OUT <= 0;  //10 / 41 = 0
    16'b00001010_00101010 : OUT <= 0;  //10 / 42 = 0
    16'b00001010_00101011 : OUT <= 0;  //10 / 43 = 0
    16'b00001010_00101100 : OUT <= 0;  //10 / 44 = 0
    16'b00001010_00101101 : OUT <= 0;  //10 / 45 = 0
    16'b00001010_00101110 : OUT <= 0;  //10 / 46 = 0
    16'b00001010_00101111 : OUT <= 0;  //10 / 47 = 0
    16'b00001010_00110000 : OUT <= 0;  //10 / 48 = 0
    16'b00001010_00110001 : OUT <= 0;  //10 / 49 = 0
    16'b00001010_00110010 : OUT <= 0;  //10 / 50 = 0
    16'b00001010_00110011 : OUT <= 0;  //10 / 51 = 0
    16'b00001010_00110100 : OUT <= 0;  //10 / 52 = 0
    16'b00001010_00110101 : OUT <= 0;  //10 / 53 = 0
    16'b00001010_00110110 : OUT <= 0;  //10 / 54 = 0
    16'b00001010_00110111 : OUT <= 0;  //10 / 55 = 0
    16'b00001010_00111000 : OUT <= 0;  //10 / 56 = 0
    16'b00001010_00111001 : OUT <= 0;  //10 / 57 = 0
    16'b00001010_00111010 : OUT <= 0;  //10 / 58 = 0
    16'b00001010_00111011 : OUT <= 0;  //10 / 59 = 0
    16'b00001010_00111100 : OUT <= 0;  //10 / 60 = 0
    16'b00001010_00111101 : OUT <= 0;  //10 / 61 = 0
    16'b00001010_00111110 : OUT <= 0;  //10 / 62 = 0
    16'b00001010_00111111 : OUT <= 0;  //10 / 63 = 0
    16'b00001010_01000000 : OUT <= 0;  //10 / 64 = 0
    16'b00001010_01000001 : OUT <= 0;  //10 / 65 = 0
    16'b00001010_01000010 : OUT <= 0;  //10 / 66 = 0
    16'b00001010_01000011 : OUT <= 0;  //10 / 67 = 0
    16'b00001010_01000100 : OUT <= 0;  //10 / 68 = 0
    16'b00001010_01000101 : OUT <= 0;  //10 / 69 = 0
    16'b00001010_01000110 : OUT <= 0;  //10 / 70 = 0
    16'b00001010_01000111 : OUT <= 0;  //10 / 71 = 0
    16'b00001010_01001000 : OUT <= 0;  //10 / 72 = 0
    16'b00001010_01001001 : OUT <= 0;  //10 / 73 = 0
    16'b00001010_01001010 : OUT <= 0;  //10 / 74 = 0
    16'b00001010_01001011 : OUT <= 0;  //10 / 75 = 0
    16'b00001010_01001100 : OUT <= 0;  //10 / 76 = 0
    16'b00001010_01001101 : OUT <= 0;  //10 / 77 = 0
    16'b00001010_01001110 : OUT <= 0;  //10 / 78 = 0
    16'b00001010_01001111 : OUT <= 0;  //10 / 79 = 0
    16'b00001010_01010000 : OUT <= 0;  //10 / 80 = 0
    16'b00001010_01010001 : OUT <= 0;  //10 / 81 = 0
    16'b00001010_01010010 : OUT <= 0;  //10 / 82 = 0
    16'b00001010_01010011 : OUT <= 0;  //10 / 83 = 0
    16'b00001010_01010100 : OUT <= 0;  //10 / 84 = 0
    16'b00001010_01010101 : OUT <= 0;  //10 / 85 = 0
    16'b00001010_01010110 : OUT <= 0;  //10 / 86 = 0
    16'b00001010_01010111 : OUT <= 0;  //10 / 87 = 0
    16'b00001010_01011000 : OUT <= 0;  //10 / 88 = 0
    16'b00001010_01011001 : OUT <= 0;  //10 / 89 = 0
    16'b00001010_01011010 : OUT <= 0;  //10 / 90 = 0
    16'b00001010_01011011 : OUT <= 0;  //10 / 91 = 0
    16'b00001010_01011100 : OUT <= 0;  //10 / 92 = 0
    16'b00001010_01011101 : OUT <= 0;  //10 / 93 = 0
    16'b00001010_01011110 : OUT <= 0;  //10 / 94 = 0
    16'b00001010_01011111 : OUT <= 0;  //10 / 95 = 0
    16'b00001010_01100000 : OUT <= 0;  //10 / 96 = 0
    16'b00001010_01100001 : OUT <= 0;  //10 / 97 = 0
    16'b00001010_01100010 : OUT <= 0;  //10 / 98 = 0
    16'b00001010_01100011 : OUT <= 0;  //10 / 99 = 0
    16'b00001010_01100100 : OUT <= 0;  //10 / 100 = 0
    16'b00001010_01100101 : OUT <= 0;  //10 / 101 = 0
    16'b00001010_01100110 : OUT <= 0;  //10 / 102 = 0
    16'b00001010_01100111 : OUT <= 0;  //10 / 103 = 0
    16'b00001010_01101000 : OUT <= 0;  //10 / 104 = 0
    16'b00001010_01101001 : OUT <= 0;  //10 / 105 = 0
    16'b00001010_01101010 : OUT <= 0;  //10 / 106 = 0
    16'b00001010_01101011 : OUT <= 0;  //10 / 107 = 0
    16'b00001010_01101100 : OUT <= 0;  //10 / 108 = 0
    16'b00001010_01101101 : OUT <= 0;  //10 / 109 = 0
    16'b00001010_01101110 : OUT <= 0;  //10 / 110 = 0
    16'b00001010_01101111 : OUT <= 0;  //10 / 111 = 0
    16'b00001010_01110000 : OUT <= 0;  //10 / 112 = 0
    16'b00001010_01110001 : OUT <= 0;  //10 / 113 = 0
    16'b00001010_01110010 : OUT <= 0;  //10 / 114 = 0
    16'b00001010_01110011 : OUT <= 0;  //10 / 115 = 0
    16'b00001010_01110100 : OUT <= 0;  //10 / 116 = 0
    16'b00001010_01110101 : OUT <= 0;  //10 / 117 = 0
    16'b00001010_01110110 : OUT <= 0;  //10 / 118 = 0
    16'b00001010_01110111 : OUT <= 0;  //10 / 119 = 0
    16'b00001010_01111000 : OUT <= 0;  //10 / 120 = 0
    16'b00001010_01111001 : OUT <= 0;  //10 / 121 = 0
    16'b00001010_01111010 : OUT <= 0;  //10 / 122 = 0
    16'b00001010_01111011 : OUT <= 0;  //10 / 123 = 0
    16'b00001010_01111100 : OUT <= 0;  //10 / 124 = 0
    16'b00001010_01111101 : OUT <= 0;  //10 / 125 = 0
    16'b00001010_01111110 : OUT <= 0;  //10 / 126 = 0
    16'b00001010_01111111 : OUT <= 0;  //10 / 127 = 0
    16'b00001010_10000000 : OUT <= 0;  //10 / 128 = 0
    16'b00001010_10000001 : OUT <= 0;  //10 / 129 = 0
    16'b00001010_10000010 : OUT <= 0;  //10 / 130 = 0
    16'b00001010_10000011 : OUT <= 0;  //10 / 131 = 0
    16'b00001010_10000100 : OUT <= 0;  //10 / 132 = 0
    16'b00001010_10000101 : OUT <= 0;  //10 / 133 = 0
    16'b00001010_10000110 : OUT <= 0;  //10 / 134 = 0
    16'b00001010_10000111 : OUT <= 0;  //10 / 135 = 0
    16'b00001010_10001000 : OUT <= 0;  //10 / 136 = 0
    16'b00001010_10001001 : OUT <= 0;  //10 / 137 = 0
    16'b00001010_10001010 : OUT <= 0;  //10 / 138 = 0
    16'b00001010_10001011 : OUT <= 0;  //10 / 139 = 0
    16'b00001010_10001100 : OUT <= 0;  //10 / 140 = 0
    16'b00001010_10001101 : OUT <= 0;  //10 / 141 = 0
    16'b00001010_10001110 : OUT <= 0;  //10 / 142 = 0
    16'b00001010_10001111 : OUT <= 0;  //10 / 143 = 0
    16'b00001010_10010000 : OUT <= 0;  //10 / 144 = 0
    16'b00001010_10010001 : OUT <= 0;  //10 / 145 = 0
    16'b00001010_10010010 : OUT <= 0;  //10 / 146 = 0
    16'b00001010_10010011 : OUT <= 0;  //10 / 147 = 0
    16'b00001010_10010100 : OUT <= 0;  //10 / 148 = 0
    16'b00001010_10010101 : OUT <= 0;  //10 / 149 = 0
    16'b00001010_10010110 : OUT <= 0;  //10 / 150 = 0
    16'b00001010_10010111 : OUT <= 0;  //10 / 151 = 0
    16'b00001010_10011000 : OUT <= 0;  //10 / 152 = 0
    16'b00001010_10011001 : OUT <= 0;  //10 / 153 = 0
    16'b00001010_10011010 : OUT <= 0;  //10 / 154 = 0
    16'b00001010_10011011 : OUT <= 0;  //10 / 155 = 0
    16'b00001010_10011100 : OUT <= 0;  //10 / 156 = 0
    16'b00001010_10011101 : OUT <= 0;  //10 / 157 = 0
    16'b00001010_10011110 : OUT <= 0;  //10 / 158 = 0
    16'b00001010_10011111 : OUT <= 0;  //10 / 159 = 0
    16'b00001010_10100000 : OUT <= 0;  //10 / 160 = 0
    16'b00001010_10100001 : OUT <= 0;  //10 / 161 = 0
    16'b00001010_10100010 : OUT <= 0;  //10 / 162 = 0
    16'b00001010_10100011 : OUT <= 0;  //10 / 163 = 0
    16'b00001010_10100100 : OUT <= 0;  //10 / 164 = 0
    16'b00001010_10100101 : OUT <= 0;  //10 / 165 = 0
    16'b00001010_10100110 : OUT <= 0;  //10 / 166 = 0
    16'b00001010_10100111 : OUT <= 0;  //10 / 167 = 0
    16'b00001010_10101000 : OUT <= 0;  //10 / 168 = 0
    16'b00001010_10101001 : OUT <= 0;  //10 / 169 = 0
    16'b00001010_10101010 : OUT <= 0;  //10 / 170 = 0
    16'b00001010_10101011 : OUT <= 0;  //10 / 171 = 0
    16'b00001010_10101100 : OUT <= 0;  //10 / 172 = 0
    16'b00001010_10101101 : OUT <= 0;  //10 / 173 = 0
    16'b00001010_10101110 : OUT <= 0;  //10 / 174 = 0
    16'b00001010_10101111 : OUT <= 0;  //10 / 175 = 0
    16'b00001010_10110000 : OUT <= 0;  //10 / 176 = 0
    16'b00001010_10110001 : OUT <= 0;  //10 / 177 = 0
    16'b00001010_10110010 : OUT <= 0;  //10 / 178 = 0
    16'b00001010_10110011 : OUT <= 0;  //10 / 179 = 0
    16'b00001010_10110100 : OUT <= 0;  //10 / 180 = 0
    16'b00001010_10110101 : OUT <= 0;  //10 / 181 = 0
    16'b00001010_10110110 : OUT <= 0;  //10 / 182 = 0
    16'b00001010_10110111 : OUT <= 0;  //10 / 183 = 0
    16'b00001010_10111000 : OUT <= 0;  //10 / 184 = 0
    16'b00001010_10111001 : OUT <= 0;  //10 / 185 = 0
    16'b00001010_10111010 : OUT <= 0;  //10 / 186 = 0
    16'b00001010_10111011 : OUT <= 0;  //10 / 187 = 0
    16'b00001010_10111100 : OUT <= 0;  //10 / 188 = 0
    16'b00001010_10111101 : OUT <= 0;  //10 / 189 = 0
    16'b00001010_10111110 : OUT <= 0;  //10 / 190 = 0
    16'b00001010_10111111 : OUT <= 0;  //10 / 191 = 0
    16'b00001010_11000000 : OUT <= 0;  //10 / 192 = 0
    16'b00001010_11000001 : OUT <= 0;  //10 / 193 = 0
    16'b00001010_11000010 : OUT <= 0;  //10 / 194 = 0
    16'b00001010_11000011 : OUT <= 0;  //10 / 195 = 0
    16'b00001010_11000100 : OUT <= 0;  //10 / 196 = 0
    16'b00001010_11000101 : OUT <= 0;  //10 / 197 = 0
    16'b00001010_11000110 : OUT <= 0;  //10 / 198 = 0
    16'b00001010_11000111 : OUT <= 0;  //10 / 199 = 0
    16'b00001010_11001000 : OUT <= 0;  //10 / 200 = 0
    16'b00001010_11001001 : OUT <= 0;  //10 / 201 = 0
    16'b00001010_11001010 : OUT <= 0;  //10 / 202 = 0
    16'b00001010_11001011 : OUT <= 0;  //10 / 203 = 0
    16'b00001010_11001100 : OUT <= 0;  //10 / 204 = 0
    16'b00001010_11001101 : OUT <= 0;  //10 / 205 = 0
    16'b00001010_11001110 : OUT <= 0;  //10 / 206 = 0
    16'b00001010_11001111 : OUT <= 0;  //10 / 207 = 0
    16'b00001010_11010000 : OUT <= 0;  //10 / 208 = 0
    16'b00001010_11010001 : OUT <= 0;  //10 / 209 = 0
    16'b00001010_11010010 : OUT <= 0;  //10 / 210 = 0
    16'b00001010_11010011 : OUT <= 0;  //10 / 211 = 0
    16'b00001010_11010100 : OUT <= 0;  //10 / 212 = 0
    16'b00001010_11010101 : OUT <= 0;  //10 / 213 = 0
    16'b00001010_11010110 : OUT <= 0;  //10 / 214 = 0
    16'b00001010_11010111 : OUT <= 0;  //10 / 215 = 0
    16'b00001010_11011000 : OUT <= 0;  //10 / 216 = 0
    16'b00001010_11011001 : OUT <= 0;  //10 / 217 = 0
    16'b00001010_11011010 : OUT <= 0;  //10 / 218 = 0
    16'b00001010_11011011 : OUT <= 0;  //10 / 219 = 0
    16'b00001010_11011100 : OUT <= 0;  //10 / 220 = 0
    16'b00001010_11011101 : OUT <= 0;  //10 / 221 = 0
    16'b00001010_11011110 : OUT <= 0;  //10 / 222 = 0
    16'b00001010_11011111 : OUT <= 0;  //10 / 223 = 0
    16'b00001010_11100000 : OUT <= 0;  //10 / 224 = 0
    16'b00001010_11100001 : OUT <= 0;  //10 / 225 = 0
    16'b00001010_11100010 : OUT <= 0;  //10 / 226 = 0
    16'b00001010_11100011 : OUT <= 0;  //10 / 227 = 0
    16'b00001010_11100100 : OUT <= 0;  //10 / 228 = 0
    16'b00001010_11100101 : OUT <= 0;  //10 / 229 = 0
    16'b00001010_11100110 : OUT <= 0;  //10 / 230 = 0
    16'b00001010_11100111 : OUT <= 0;  //10 / 231 = 0
    16'b00001010_11101000 : OUT <= 0;  //10 / 232 = 0
    16'b00001010_11101001 : OUT <= 0;  //10 / 233 = 0
    16'b00001010_11101010 : OUT <= 0;  //10 / 234 = 0
    16'b00001010_11101011 : OUT <= 0;  //10 / 235 = 0
    16'b00001010_11101100 : OUT <= 0;  //10 / 236 = 0
    16'b00001010_11101101 : OUT <= 0;  //10 / 237 = 0
    16'b00001010_11101110 : OUT <= 0;  //10 / 238 = 0
    16'b00001010_11101111 : OUT <= 0;  //10 / 239 = 0
    16'b00001010_11110000 : OUT <= 0;  //10 / 240 = 0
    16'b00001010_11110001 : OUT <= 0;  //10 / 241 = 0
    16'b00001010_11110010 : OUT <= 0;  //10 / 242 = 0
    16'b00001010_11110011 : OUT <= 0;  //10 / 243 = 0
    16'b00001010_11110100 : OUT <= 0;  //10 / 244 = 0
    16'b00001010_11110101 : OUT <= 0;  //10 / 245 = 0
    16'b00001010_11110110 : OUT <= 0;  //10 / 246 = 0
    16'b00001010_11110111 : OUT <= 0;  //10 / 247 = 0
    16'b00001010_11111000 : OUT <= 0;  //10 / 248 = 0
    16'b00001010_11111001 : OUT <= 0;  //10 / 249 = 0
    16'b00001010_11111010 : OUT <= 0;  //10 / 250 = 0
    16'b00001010_11111011 : OUT <= 0;  //10 / 251 = 0
    16'b00001010_11111100 : OUT <= 0;  //10 / 252 = 0
    16'b00001010_11111101 : OUT <= 0;  //10 / 253 = 0
    16'b00001010_11111110 : OUT <= 0;  //10 / 254 = 0
    16'b00001010_11111111 : OUT <= 0;  //10 / 255 = 0
    16'b00001011_00000000 : OUT <= 0;  //11 / 0 = 0
    16'b00001011_00000001 : OUT <= 11;  //11 / 1 = 11
    16'b00001011_00000010 : OUT <= 5;  //11 / 2 = 5
    16'b00001011_00000011 : OUT <= 3;  //11 / 3 = 3
    16'b00001011_00000100 : OUT <= 2;  //11 / 4 = 2
    16'b00001011_00000101 : OUT <= 2;  //11 / 5 = 2
    16'b00001011_00000110 : OUT <= 1;  //11 / 6 = 1
    16'b00001011_00000111 : OUT <= 1;  //11 / 7 = 1
    16'b00001011_00001000 : OUT <= 1;  //11 / 8 = 1
    16'b00001011_00001001 : OUT <= 1;  //11 / 9 = 1
    16'b00001011_00001010 : OUT <= 1;  //11 / 10 = 1
    16'b00001011_00001011 : OUT <= 1;  //11 / 11 = 1
    16'b00001011_00001100 : OUT <= 0;  //11 / 12 = 0
    16'b00001011_00001101 : OUT <= 0;  //11 / 13 = 0
    16'b00001011_00001110 : OUT <= 0;  //11 / 14 = 0
    16'b00001011_00001111 : OUT <= 0;  //11 / 15 = 0
    16'b00001011_00010000 : OUT <= 0;  //11 / 16 = 0
    16'b00001011_00010001 : OUT <= 0;  //11 / 17 = 0
    16'b00001011_00010010 : OUT <= 0;  //11 / 18 = 0
    16'b00001011_00010011 : OUT <= 0;  //11 / 19 = 0
    16'b00001011_00010100 : OUT <= 0;  //11 / 20 = 0
    16'b00001011_00010101 : OUT <= 0;  //11 / 21 = 0
    16'b00001011_00010110 : OUT <= 0;  //11 / 22 = 0
    16'b00001011_00010111 : OUT <= 0;  //11 / 23 = 0
    16'b00001011_00011000 : OUT <= 0;  //11 / 24 = 0
    16'b00001011_00011001 : OUT <= 0;  //11 / 25 = 0
    16'b00001011_00011010 : OUT <= 0;  //11 / 26 = 0
    16'b00001011_00011011 : OUT <= 0;  //11 / 27 = 0
    16'b00001011_00011100 : OUT <= 0;  //11 / 28 = 0
    16'b00001011_00011101 : OUT <= 0;  //11 / 29 = 0
    16'b00001011_00011110 : OUT <= 0;  //11 / 30 = 0
    16'b00001011_00011111 : OUT <= 0;  //11 / 31 = 0
    16'b00001011_00100000 : OUT <= 0;  //11 / 32 = 0
    16'b00001011_00100001 : OUT <= 0;  //11 / 33 = 0
    16'b00001011_00100010 : OUT <= 0;  //11 / 34 = 0
    16'b00001011_00100011 : OUT <= 0;  //11 / 35 = 0
    16'b00001011_00100100 : OUT <= 0;  //11 / 36 = 0
    16'b00001011_00100101 : OUT <= 0;  //11 / 37 = 0
    16'b00001011_00100110 : OUT <= 0;  //11 / 38 = 0
    16'b00001011_00100111 : OUT <= 0;  //11 / 39 = 0
    16'b00001011_00101000 : OUT <= 0;  //11 / 40 = 0
    16'b00001011_00101001 : OUT <= 0;  //11 / 41 = 0
    16'b00001011_00101010 : OUT <= 0;  //11 / 42 = 0
    16'b00001011_00101011 : OUT <= 0;  //11 / 43 = 0
    16'b00001011_00101100 : OUT <= 0;  //11 / 44 = 0
    16'b00001011_00101101 : OUT <= 0;  //11 / 45 = 0
    16'b00001011_00101110 : OUT <= 0;  //11 / 46 = 0
    16'b00001011_00101111 : OUT <= 0;  //11 / 47 = 0
    16'b00001011_00110000 : OUT <= 0;  //11 / 48 = 0
    16'b00001011_00110001 : OUT <= 0;  //11 / 49 = 0
    16'b00001011_00110010 : OUT <= 0;  //11 / 50 = 0
    16'b00001011_00110011 : OUT <= 0;  //11 / 51 = 0
    16'b00001011_00110100 : OUT <= 0;  //11 / 52 = 0
    16'b00001011_00110101 : OUT <= 0;  //11 / 53 = 0
    16'b00001011_00110110 : OUT <= 0;  //11 / 54 = 0
    16'b00001011_00110111 : OUT <= 0;  //11 / 55 = 0
    16'b00001011_00111000 : OUT <= 0;  //11 / 56 = 0
    16'b00001011_00111001 : OUT <= 0;  //11 / 57 = 0
    16'b00001011_00111010 : OUT <= 0;  //11 / 58 = 0
    16'b00001011_00111011 : OUT <= 0;  //11 / 59 = 0
    16'b00001011_00111100 : OUT <= 0;  //11 / 60 = 0
    16'b00001011_00111101 : OUT <= 0;  //11 / 61 = 0
    16'b00001011_00111110 : OUT <= 0;  //11 / 62 = 0
    16'b00001011_00111111 : OUT <= 0;  //11 / 63 = 0
    16'b00001011_01000000 : OUT <= 0;  //11 / 64 = 0
    16'b00001011_01000001 : OUT <= 0;  //11 / 65 = 0
    16'b00001011_01000010 : OUT <= 0;  //11 / 66 = 0
    16'b00001011_01000011 : OUT <= 0;  //11 / 67 = 0
    16'b00001011_01000100 : OUT <= 0;  //11 / 68 = 0
    16'b00001011_01000101 : OUT <= 0;  //11 / 69 = 0
    16'b00001011_01000110 : OUT <= 0;  //11 / 70 = 0
    16'b00001011_01000111 : OUT <= 0;  //11 / 71 = 0
    16'b00001011_01001000 : OUT <= 0;  //11 / 72 = 0
    16'b00001011_01001001 : OUT <= 0;  //11 / 73 = 0
    16'b00001011_01001010 : OUT <= 0;  //11 / 74 = 0
    16'b00001011_01001011 : OUT <= 0;  //11 / 75 = 0
    16'b00001011_01001100 : OUT <= 0;  //11 / 76 = 0
    16'b00001011_01001101 : OUT <= 0;  //11 / 77 = 0
    16'b00001011_01001110 : OUT <= 0;  //11 / 78 = 0
    16'b00001011_01001111 : OUT <= 0;  //11 / 79 = 0
    16'b00001011_01010000 : OUT <= 0;  //11 / 80 = 0
    16'b00001011_01010001 : OUT <= 0;  //11 / 81 = 0
    16'b00001011_01010010 : OUT <= 0;  //11 / 82 = 0
    16'b00001011_01010011 : OUT <= 0;  //11 / 83 = 0
    16'b00001011_01010100 : OUT <= 0;  //11 / 84 = 0
    16'b00001011_01010101 : OUT <= 0;  //11 / 85 = 0
    16'b00001011_01010110 : OUT <= 0;  //11 / 86 = 0
    16'b00001011_01010111 : OUT <= 0;  //11 / 87 = 0
    16'b00001011_01011000 : OUT <= 0;  //11 / 88 = 0
    16'b00001011_01011001 : OUT <= 0;  //11 / 89 = 0
    16'b00001011_01011010 : OUT <= 0;  //11 / 90 = 0
    16'b00001011_01011011 : OUT <= 0;  //11 / 91 = 0
    16'b00001011_01011100 : OUT <= 0;  //11 / 92 = 0
    16'b00001011_01011101 : OUT <= 0;  //11 / 93 = 0
    16'b00001011_01011110 : OUT <= 0;  //11 / 94 = 0
    16'b00001011_01011111 : OUT <= 0;  //11 / 95 = 0
    16'b00001011_01100000 : OUT <= 0;  //11 / 96 = 0
    16'b00001011_01100001 : OUT <= 0;  //11 / 97 = 0
    16'b00001011_01100010 : OUT <= 0;  //11 / 98 = 0
    16'b00001011_01100011 : OUT <= 0;  //11 / 99 = 0
    16'b00001011_01100100 : OUT <= 0;  //11 / 100 = 0
    16'b00001011_01100101 : OUT <= 0;  //11 / 101 = 0
    16'b00001011_01100110 : OUT <= 0;  //11 / 102 = 0
    16'b00001011_01100111 : OUT <= 0;  //11 / 103 = 0
    16'b00001011_01101000 : OUT <= 0;  //11 / 104 = 0
    16'b00001011_01101001 : OUT <= 0;  //11 / 105 = 0
    16'b00001011_01101010 : OUT <= 0;  //11 / 106 = 0
    16'b00001011_01101011 : OUT <= 0;  //11 / 107 = 0
    16'b00001011_01101100 : OUT <= 0;  //11 / 108 = 0
    16'b00001011_01101101 : OUT <= 0;  //11 / 109 = 0
    16'b00001011_01101110 : OUT <= 0;  //11 / 110 = 0
    16'b00001011_01101111 : OUT <= 0;  //11 / 111 = 0
    16'b00001011_01110000 : OUT <= 0;  //11 / 112 = 0
    16'b00001011_01110001 : OUT <= 0;  //11 / 113 = 0
    16'b00001011_01110010 : OUT <= 0;  //11 / 114 = 0
    16'b00001011_01110011 : OUT <= 0;  //11 / 115 = 0
    16'b00001011_01110100 : OUT <= 0;  //11 / 116 = 0
    16'b00001011_01110101 : OUT <= 0;  //11 / 117 = 0
    16'b00001011_01110110 : OUT <= 0;  //11 / 118 = 0
    16'b00001011_01110111 : OUT <= 0;  //11 / 119 = 0
    16'b00001011_01111000 : OUT <= 0;  //11 / 120 = 0
    16'b00001011_01111001 : OUT <= 0;  //11 / 121 = 0
    16'b00001011_01111010 : OUT <= 0;  //11 / 122 = 0
    16'b00001011_01111011 : OUT <= 0;  //11 / 123 = 0
    16'b00001011_01111100 : OUT <= 0;  //11 / 124 = 0
    16'b00001011_01111101 : OUT <= 0;  //11 / 125 = 0
    16'b00001011_01111110 : OUT <= 0;  //11 / 126 = 0
    16'b00001011_01111111 : OUT <= 0;  //11 / 127 = 0
    16'b00001011_10000000 : OUT <= 0;  //11 / 128 = 0
    16'b00001011_10000001 : OUT <= 0;  //11 / 129 = 0
    16'b00001011_10000010 : OUT <= 0;  //11 / 130 = 0
    16'b00001011_10000011 : OUT <= 0;  //11 / 131 = 0
    16'b00001011_10000100 : OUT <= 0;  //11 / 132 = 0
    16'b00001011_10000101 : OUT <= 0;  //11 / 133 = 0
    16'b00001011_10000110 : OUT <= 0;  //11 / 134 = 0
    16'b00001011_10000111 : OUT <= 0;  //11 / 135 = 0
    16'b00001011_10001000 : OUT <= 0;  //11 / 136 = 0
    16'b00001011_10001001 : OUT <= 0;  //11 / 137 = 0
    16'b00001011_10001010 : OUT <= 0;  //11 / 138 = 0
    16'b00001011_10001011 : OUT <= 0;  //11 / 139 = 0
    16'b00001011_10001100 : OUT <= 0;  //11 / 140 = 0
    16'b00001011_10001101 : OUT <= 0;  //11 / 141 = 0
    16'b00001011_10001110 : OUT <= 0;  //11 / 142 = 0
    16'b00001011_10001111 : OUT <= 0;  //11 / 143 = 0
    16'b00001011_10010000 : OUT <= 0;  //11 / 144 = 0
    16'b00001011_10010001 : OUT <= 0;  //11 / 145 = 0
    16'b00001011_10010010 : OUT <= 0;  //11 / 146 = 0
    16'b00001011_10010011 : OUT <= 0;  //11 / 147 = 0
    16'b00001011_10010100 : OUT <= 0;  //11 / 148 = 0
    16'b00001011_10010101 : OUT <= 0;  //11 / 149 = 0
    16'b00001011_10010110 : OUT <= 0;  //11 / 150 = 0
    16'b00001011_10010111 : OUT <= 0;  //11 / 151 = 0
    16'b00001011_10011000 : OUT <= 0;  //11 / 152 = 0
    16'b00001011_10011001 : OUT <= 0;  //11 / 153 = 0
    16'b00001011_10011010 : OUT <= 0;  //11 / 154 = 0
    16'b00001011_10011011 : OUT <= 0;  //11 / 155 = 0
    16'b00001011_10011100 : OUT <= 0;  //11 / 156 = 0
    16'b00001011_10011101 : OUT <= 0;  //11 / 157 = 0
    16'b00001011_10011110 : OUT <= 0;  //11 / 158 = 0
    16'b00001011_10011111 : OUT <= 0;  //11 / 159 = 0
    16'b00001011_10100000 : OUT <= 0;  //11 / 160 = 0
    16'b00001011_10100001 : OUT <= 0;  //11 / 161 = 0
    16'b00001011_10100010 : OUT <= 0;  //11 / 162 = 0
    16'b00001011_10100011 : OUT <= 0;  //11 / 163 = 0
    16'b00001011_10100100 : OUT <= 0;  //11 / 164 = 0
    16'b00001011_10100101 : OUT <= 0;  //11 / 165 = 0
    16'b00001011_10100110 : OUT <= 0;  //11 / 166 = 0
    16'b00001011_10100111 : OUT <= 0;  //11 / 167 = 0
    16'b00001011_10101000 : OUT <= 0;  //11 / 168 = 0
    16'b00001011_10101001 : OUT <= 0;  //11 / 169 = 0
    16'b00001011_10101010 : OUT <= 0;  //11 / 170 = 0
    16'b00001011_10101011 : OUT <= 0;  //11 / 171 = 0
    16'b00001011_10101100 : OUT <= 0;  //11 / 172 = 0
    16'b00001011_10101101 : OUT <= 0;  //11 / 173 = 0
    16'b00001011_10101110 : OUT <= 0;  //11 / 174 = 0
    16'b00001011_10101111 : OUT <= 0;  //11 / 175 = 0
    16'b00001011_10110000 : OUT <= 0;  //11 / 176 = 0
    16'b00001011_10110001 : OUT <= 0;  //11 / 177 = 0
    16'b00001011_10110010 : OUT <= 0;  //11 / 178 = 0
    16'b00001011_10110011 : OUT <= 0;  //11 / 179 = 0
    16'b00001011_10110100 : OUT <= 0;  //11 / 180 = 0
    16'b00001011_10110101 : OUT <= 0;  //11 / 181 = 0
    16'b00001011_10110110 : OUT <= 0;  //11 / 182 = 0
    16'b00001011_10110111 : OUT <= 0;  //11 / 183 = 0
    16'b00001011_10111000 : OUT <= 0;  //11 / 184 = 0
    16'b00001011_10111001 : OUT <= 0;  //11 / 185 = 0
    16'b00001011_10111010 : OUT <= 0;  //11 / 186 = 0
    16'b00001011_10111011 : OUT <= 0;  //11 / 187 = 0
    16'b00001011_10111100 : OUT <= 0;  //11 / 188 = 0
    16'b00001011_10111101 : OUT <= 0;  //11 / 189 = 0
    16'b00001011_10111110 : OUT <= 0;  //11 / 190 = 0
    16'b00001011_10111111 : OUT <= 0;  //11 / 191 = 0
    16'b00001011_11000000 : OUT <= 0;  //11 / 192 = 0
    16'b00001011_11000001 : OUT <= 0;  //11 / 193 = 0
    16'b00001011_11000010 : OUT <= 0;  //11 / 194 = 0
    16'b00001011_11000011 : OUT <= 0;  //11 / 195 = 0
    16'b00001011_11000100 : OUT <= 0;  //11 / 196 = 0
    16'b00001011_11000101 : OUT <= 0;  //11 / 197 = 0
    16'b00001011_11000110 : OUT <= 0;  //11 / 198 = 0
    16'b00001011_11000111 : OUT <= 0;  //11 / 199 = 0
    16'b00001011_11001000 : OUT <= 0;  //11 / 200 = 0
    16'b00001011_11001001 : OUT <= 0;  //11 / 201 = 0
    16'b00001011_11001010 : OUT <= 0;  //11 / 202 = 0
    16'b00001011_11001011 : OUT <= 0;  //11 / 203 = 0
    16'b00001011_11001100 : OUT <= 0;  //11 / 204 = 0
    16'b00001011_11001101 : OUT <= 0;  //11 / 205 = 0
    16'b00001011_11001110 : OUT <= 0;  //11 / 206 = 0
    16'b00001011_11001111 : OUT <= 0;  //11 / 207 = 0
    16'b00001011_11010000 : OUT <= 0;  //11 / 208 = 0
    16'b00001011_11010001 : OUT <= 0;  //11 / 209 = 0
    16'b00001011_11010010 : OUT <= 0;  //11 / 210 = 0
    16'b00001011_11010011 : OUT <= 0;  //11 / 211 = 0
    16'b00001011_11010100 : OUT <= 0;  //11 / 212 = 0
    16'b00001011_11010101 : OUT <= 0;  //11 / 213 = 0
    16'b00001011_11010110 : OUT <= 0;  //11 / 214 = 0
    16'b00001011_11010111 : OUT <= 0;  //11 / 215 = 0
    16'b00001011_11011000 : OUT <= 0;  //11 / 216 = 0
    16'b00001011_11011001 : OUT <= 0;  //11 / 217 = 0
    16'b00001011_11011010 : OUT <= 0;  //11 / 218 = 0
    16'b00001011_11011011 : OUT <= 0;  //11 / 219 = 0
    16'b00001011_11011100 : OUT <= 0;  //11 / 220 = 0
    16'b00001011_11011101 : OUT <= 0;  //11 / 221 = 0
    16'b00001011_11011110 : OUT <= 0;  //11 / 222 = 0
    16'b00001011_11011111 : OUT <= 0;  //11 / 223 = 0
    16'b00001011_11100000 : OUT <= 0;  //11 / 224 = 0
    16'b00001011_11100001 : OUT <= 0;  //11 / 225 = 0
    16'b00001011_11100010 : OUT <= 0;  //11 / 226 = 0
    16'b00001011_11100011 : OUT <= 0;  //11 / 227 = 0
    16'b00001011_11100100 : OUT <= 0;  //11 / 228 = 0
    16'b00001011_11100101 : OUT <= 0;  //11 / 229 = 0
    16'b00001011_11100110 : OUT <= 0;  //11 / 230 = 0
    16'b00001011_11100111 : OUT <= 0;  //11 / 231 = 0
    16'b00001011_11101000 : OUT <= 0;  //11 / 232 = 0
    16'b00001011_11101001 : OUT <= 0;  //11 / 233 = 0
    16'b00001011_11101010 : OUT <= 0;  //11 / 234 = 0
    16'b00001011_11101011 : OUT <= 0;  //11 / 235 = 0
    16'b00001011_11101100 : OUT <= 0;  //11 / 236 = 0
    16'b00001011_11101101 : OUT <= 0;  //11 / 237 = 0
    16'b00001011_11101110 : OUT <= 0;  //11 / 238 = 0
    16'b00001011_11101111 : OUT <= 0;  //11 / 239 = 0
    16'b00001011_11110000 : OUT <= 0;  //11 / 240 = 0
    16'b00001011_11110001 : OUT <= 0;  //11 / 241 = 0
    16'b00001011_11110010 : OUT <= 0;  //11 / 242 = 0
    16'b00001011_11110011 : OUT <= 0;  //11 / 243 = 0
    16'b00001011_11110100 : OUT <= 0;  //11 / 244 = 0
    16'b00001011_11110101 : OUT <= 0;  //11 / 245 = 0
    16'b00001011_11110110 : OUT <= 0;  //11 / 246 = 0
    16'b00001011_11110111 : OUT <= 0;  //11 / 247 = 0
    16'b00001011_11111000 : OUT <= 0;  //11 / 248 = 0
    16'b00001011_11111001 : OUT <= 0;  //11 / 249 = 0
    16'b00001011_11111010 : OUT <= 0;  //11 / 250 = 0
    16'b00001011_11111011 : OUT <= 0;  //11 / 251 = 0
    16'b00001011_11111100 : OUT <= 0;  //11 / 252 = 0
    16'b00001011_11111101 : OUT <= 0;  //11 / 253 = 0
    16'b00001011_11111110 : OUT <= 0;  //11 / 254 = 0
    16'b00001011_11111111 : OUT <= 0;  //11 / 255 = 0
    16'b00001100_00000000 : OUT <= 0;  //12 / 0 = 0
    16'b00001100_00000001 : OUT <= 12;  //12 / 1 = 12
    16'b00001100_00000010 : OUT <= 6;  //12 / 2 = 6
    16'b00001100_00000011 : OUT <= 4;  //12 / 3 = 4
    16'b00001100_00000100 : OUT <= 3;  //12 / 4 = 3
    16'b00001100_00000101 : OUT <= 2;  //12 / 5 = 2
    16'b00001100_00000110 : OUT <= 2;  //12 / 6 = 2
    16'b00001100_00000111 : OUT <= 1;  //12 / 7 = 1
    16'b00001100_00001000 : OUT <= 1;  //12 / 8 = 1
    16'b00001100_00001001 : OUT <= 1;  //12 / 9 = 1
    16'b00001100_00001010 : OUT <= 1;  //12 / 10 = 1
    16'b00001100_00001011 : OUT <= 1;  //12 / 11 = 1
    16'b00001100_00001100 : OUT <= 1;  //12 / 12 = 1
    16'b00001100_00001101 : OUT <= 0;  //12 / 13 = 0
    16'b00001100_00001110 : OUT <= 0;  //12 / 14 = 0
    16'b00001100_00001111 : OUT <= 0;  //12 / 15 = 0
    16'b00001100_00010000 : OUT <= 0;  //12 / 16 = 0
    16'b00001100_00010001 : OUT <= 0;  //12 / 17 = 0
    16'b00001100_00010010 : OUT <= 0;  //12 / 18 = 0
    16'b00001100_00010011 : OUT <= 0;  //12 / 19 = 0
    16'b00001100_00010100 : OUT <= 0;  //12 / 20 = 0
    16'b00001100_00010101 : OUT <= 0;  //12 / 21 = 0
    16'b00001100_00010110 : OUT <= 0;  //12 / 22 = 0
    16'b00001100_00010111 : OUT <= 0;  //12 / 23 = 0
    16'b00001100_00011000 : OUT <= 0;  //12 / 24 = 0
    16'b00001100_00011001 : OUT <= 0;  //12 / 25 = 0
    16'b00001100_00011010 : OUT <= 0;  //12 / 26 = 0
    16'b00001100_00011011 : OUT <= 0;  //12 / 27 = 0
    16'b00001100_00011100 : OUT <= 0;  //12 / 28 = 0
    16'b00001100_00011101 : OUT <= 0;  //12 / 29 = 0
    16'b00001100_00011110 : OUT <= 0;  //12 / 30 = 0
    16'b00001100_00011111 : OUT <= 0;  //12 / 31 = 0
    16'b00001100_00100000 : OUT <= 0;  //12 / 32 = 0
    16'b00001100_00100001 : OUT <= 0;  //12 / 33 = 0
    16'b00001100_00100010 : OUT <= 0;  //12 / 34 = 0
    16'b00001100_00100011 : OUT <= 0;  //12 / 35 = 0
    16'b00001100_00100100 : OUT <= 0;  //12 / 36 = 0
    16'b00001100_00100101 : OUT <= 0;  //12 / 37 = 0
    16'b00001100_00100110 : OUT <= 0;  //12 / 38 = 0
    16'b00001100_00100111 : OUT <= 0;  //12 / 39 = 0
    16'b00001100_00101000 : OUT <= 0;  //12 / 40 = 0
    16'b00001100_00101001 : OUT <= 0;  //12 / 41 = 0
    16'b00001100_00101010 : OUT <= 0;  //12 / 42 = 0
    16'b00001100_00101011 : OUT <= 0;  //12 / 43 = 0
    16'b00001100_00101100 : OUT <= 0;  //12 / 44 = 0
    16'b00001100_00101101 : OUT <= 0;  //12 / 45 = 0
    16'b00001100_00101110 : OUT <= 0;  //12 / 46 = 0
    16'b00001100_00101111 : OUT <= 0;  //12 / 47 = 0
    16'b00001100_00110000 : OUT <= 0;  //12 / 48 = 0
    16'b00001100_00110001 : OUT <= 0;  //12 / 49 = 0
    16'b00001100_00110010 : OUT <= 0;  //12 / 50 = 0
    16'b00001100_00110011 : OUT <= 0;  //12 / 51 = 0
    16'b00001100_00110100 : OUT <= 0;  //12 / 52 = 0
    16'b00001100_00110101 : OUT <= 0;  //12 / 53 = 0
    16'b00001100_00110110 : OUT <= 0;  //12 / 54 = 0
    16'b00001100_00110111 : OUT <= 0;  //12 / 55 = 0
    16'b00001100_00111000 : OUT <= 0;  //12 / 56 = 0
    16'b00001100_00111001 : OUT <= 0;  //12 / 57 = 0
    16'b00001100_00111010 : OUT <= 0;  //12 / 58 = 0
    16'b00001100_00111011 : OUT <= 0;  //12 / 59 = 0
    16'b00001100_00111100 : OUT <= 0;  //12 / 60 = 0
    16'b00001100_00111101 : OUT <= 0;  //12 / 61 = 0
    16'b00001100_00111110 : OUT <= 0;  //12 / 62 = 0
    16'b00001100_00111111 : OUT <= 0;  //12 / 63 = 0
    16'b00001100_01000000 : OUT <= 0;  //12 / 64 = 0
    16'b00001100_01000001 : OUT <= 0;  //12 / 65 = 0
    16'b00001100_01000010 : OUT <= 0;  //12 / 66 = 0
    16'b00001100_01000011 : OUT <= 0;  //12 / 67 = 0
    16'b00001100_01000100 : OUT <= 0;  //12 / 68 = 0
    16'b00001100_01000101 : OUT <= 0;  //12 / 69 = 0
    16'b00001100_01000110 : OUT <= 0;  //12 / 70 = 0
    16'b00001100_01000111 : OUT <= 0;  //12 / 71 = 0
    16'b00001100_01001000 : OUT <= 0;  //12 / 72 = 0
    16'b00001100_01001001 : OUT <= 0;  //12 / 73 = 0
    16'b00001100_01001010 : OUT <= 0;  //12 / 74 = 0
    16'b00001100_01001011 : OUT <= 0;  //12 / 75 = 0
    16'b00001100_01001100 : OUT <= 0;  //12 / 76 = 0
    16'b00001100_01001101 : OUT <= 0;  //12 / 77 = 0
    16'b00001100_01001110 : OUT <= 0;  //12 / 78 = 0
    16'b00001100_01001111 : OUT <= 0;  //12 / 79 = 0
    16'b00001100_01010000 : OUT <= 0;  //12 / 80 = 0
    16'b00001100_01010001 : OUT <= 0;  //12 / 81 = 0
    16'b00001100_01010010 : OUT <= 0;  //12 / 82 = 0
    16'b00001100_01010011 : OUT <= 0;  //12 / 83 = 0
    16'b00001100_01010100 : OUT <= 0;  //12 / 84 = 0
    16'b00001100_01010101 : OUT <= 0;  //12 / 85 = 0
    16'b00001100_01010110 : OUT <= 0;  //12 / 86 = 0
    16'b00001100_01010111 : OUT <= 0;  //12 / 87 = 0
    16'b00001100_01011000 : OUT <= 0;  //12 / 88 = 0
    16'b00001100_01011001 : OUT <= 0;  //12 / 89 = 0
    16'b00001100_01011010 : OUT <= 0;  //12 / 90 = 0
    16'b00001100_01011011 : OUT <= 0;  //12 / 91 = 0
    16'b00001100_01011100 : OUT <= 0;  //12 / 92 = 0
    16'b00001100_01011101 : OUT <= 0;  //12 / 93 = 0
    16'b00001100_01011110 : OUT <= 0;  //12 / 94 = 0
    16'b00001100_01011111 : OUT <= 0;  //12 / 95 = 0
    16'b00001100_01100000 : OUT <= 0;  //12 / 96 = 0
    16'b00001100_01100001 : OUT <= 0;  //12 / 97 = 0
    16'b00001100_01100010 : OUT <= 0;  //12 / 98 = 0
    16'b00001100_01100011 : OUT <= 0;  //12 / 99 = 0
    16'b00001100_01100100 : OUT <= 0;  //12 / 100 = 0
    16'b00001100_01100101 : OUT <= 0;  //12 / 101 = 0
    16'b00001100_01100110 : OUT <= 0;  //12 / 102 = 0
    16'b00001100_01100111 : OUT <= 0;  //12 / 103 = 0
    16'b00001100_01101000 : OUT <= 0;  //12 / 104 = 0
    16'b00001100_01101001 : OUT <= 0;  //12 / 105 = 0
    16'b00001100_01101010 : OUT <= 0;  //12 / 106 = 0
    16'b00001100_01101011 : OUT <= 0;  //12 / 107 = 0
    16'b00001100_01101100 : OUT <= 0;  //12 / 108 = 0
    16'b00001100_01101101 : OUT <= 0;  //12 / 109 = 0
    16'b00001100_01101110 : OUT <= 0;  //12 / 110 = 0
    16'b00001100_01101111 : OUT <= 0;  //12 / 111 = 0
    16'b00001100_01110000 : OUT <= 0;  //12 / 112 = 0
    16'b00001100_01110001 : OUT <= 0;  //12 / 113 = 0
    16'b00001100_01110010 : OUT <= 0;  //12 / 114 = 0
    16'b00001100_01110011 : OUT <= 0;  //12 / 115 = 0
    16'b00001100_01110100 : OUT <= 0;  //12 / 116 = 0
    16'b00001100_01110101 : OUT <= 0;  //12 / 117 = 0
    16'b00001100_01110110 : OUT <= 0;  //12 / 118 = 0
    16'b00001100_01110111 : OUT <= 0;  //12 / 119 = 0
    16'b00001100_01111000 : OUT <= 0;  //12 / 120 = 0
    16'b00001100_01111001 : OUT <= 0;  //12 / 121 = 0
    16'b00001100_01111010 : OUT <= 0;  //12 / 122 = 0
    16'b00001100_01111011 : OUT <= 0;  //12 / 123 = 0
    16'b00001100_01111100 : OUT <= 0;  //12 / 124 = 0
    16'b00001100_01111101 : OUT <= 0;  //12 / 125 = 0
    16'b00001100_01111110 : OUT <= 0;  //12 / 126 = 0
    16'b00001100_01111111 : OUT <= 0;  //12 / 127 = 0
    16'b00001100_10000000 : OUT <= 0;  //12 / 128 = 0
    16'b00001100_10000001 : OUT <= 0;  //12 / 129 = 0
    16'b00001100_10000010 : OUT <= 0;  //12 / 130 = 0
    16'b00001100_10000011 : OUT <= 0;  //12 / 131 = 0
    16'b00001100_10000100 : OUT <= 0;  //12 / 132 = 0
    16'b00001100_10000101 : OUT <= 0;  //12 / 133 = 0
    16'b00001100_10000110 : OUT <= 0;  //12 / 134 = 0
    16'b00001100_10000111 : OUT <= 0;  //12 / 135 = 0
    16'b00001100_10001000 : OUT <= 0;  //12 / 136 = 0
    16'b00001100_10001001 : OUT <= 0;  //12 / 137 = 0
    16'b00001100_10001010 : OUT <= 0;  //12 / 138 = 0
    16'b00001100_10001011 : OUT <= 0;  //12 / 139 = 0
    16'b00001100_10001100 : OUT <= 0;  //12 / 140 = 0
    16'b00001100_10001101 : OUT <= 0;  //12 / 141 = 0
    16'b00001100_10001110 : OUT <= 0;  //12 / 142 = 0
    16'b00001100_10001111 : OUT <= 0;  //12 / 143 = 0
    16'b00001100_10010000 : OUT <= 0;  //12 / 144 = 0
    16'b00001100_10010001 : OUT <= 0;  //12 / 145 = 0
    16'b00001100_10010010 : OUT <= 0;  //12 / 146 = 0
    16'b00001100_10010011 : OUT <= 0;  //12 / 147 = 0
    16'b00001100_10010100 : OUT <= 0;  //12 / 148 = 0
    16'b00001100_10010101 : OUT <= 0;  //12 / 149 = 0
    16'b00001100_10010110 : OUT <= 0;  //12 / 150 = 0
    16'b00001100_10010111 : OUT <= 0;  //12 / 151 = 0
    16'b00001100_10011000 : OUT <= 0;  //12 / 152 = 0
    16'b00001100_10011001 : OUT <= 0;  //12 / 153 = 0
    16'b00001100_10011010 : OUT <= 0;  //12 / 154 = 0
    16'b00001100_10011011 : OUT <= 0;  //12 / 155 = 0
    16'b00001100_10011100 : OUT <= 0;  //12 / 156 = 0
    16'b00001100_10011101 : OUT <= 0;  //12 / 157 = 0
    16'b00001100_10011110 : OUT <= 0;  //12 / 158 = 0
    16'b00001100_10011111 : OUT <= 0;  //12 / 159 = 0
    16'b00001100_10100000 : OUT <= 0;  //12 / 160 = 0
    16'b00001100_10100001 : OUT <= 0;  //12 / 161 = 0
    16'b00001100_10100010 : OUT <= 0;  //12 / 162 = 0
    16'b00001100_10100011 : OUT <= 0;  //12 / 163 = 0
    16'b00001100_10100100 : OUT <= 0;  //12 / 164 = 0
    16'b00001100_10100101 : OUT <= 0;  //12 / 165 = 0
    16'b00001100_10100110 : OUT <= 0;  //12 / 166 = 0
    16'b00001100_10100111 : OUT <= 0;  //12 / 167 = 0
    16'b00001100_10101000 : OUT <= 0;  //12 / 168 = 0
    16'b00001100_10101001 : OUT <= 0;  //12 / 169 = 0
    16'b00001100_10101010 : OUT <= 0;  //12 / 170 = 0
    16'b00001100_10101011 : OUT <= 0;  //12 / 171 = 0
    16'b00001100_10101100 : OUT <= 0;  //12 / 172 = 0
    16'b00001100_10101101 : OUT <= 0;  //12 / 173 = 0
    16'b00001100_10101110 : OUT <= 0;  //12 / 174 = 0
    16'b00001100_10101111 : OUT <= 0;  //12 / 175 = 0
    16'b00001100_10110000 : OUT <= 0;  //12 / 176 = 0
    16'b00001100_10110001 : OUT <= 0;  //12 / 177 = 0
    16'b00001100_10110010 : OUT <= 0;  //12 / 178 = 0
    16'b00001100_10110011 : OUT <= 0;  //12 / 179 = 0
    16'b00001100_10110100 : OUT <= 0;  //12 / 180 = 0
    16'b00001100_10110101 : OUT <= 0;  //12 / 181 = 0
    16'b00001100_10110110 : OUT <= 0;  //12 / 182 = 0
    16'b00001100_10110111 : OUT <= 0;  //12 / 183 = 0
    16'b00001100_10111000 : OUT <= 0;  //12 / 184 = 0
    16'b00001100_10111001 : OUT <= 0;  //12 / 185 = 0
    16'b00001100_10111010 : OUT <= 0;  //12 / 186 = 0
    16'b00001100_10111011 : OUT <= 0;  //12 / 187 = 0
    16'b00001100_10111100 : OUT <= 0;  //12 / 188 = 0
    16'b00001100_10111101 : OUT <= 0;  //12 / 189 = 0
    16'b00001100_10111110 : OUT <= 0;  //12 / 190 = 0
    16'b00001100_10111111 : OUT <= 0;  //12 / 191 = 0
    16'b00001100_11000000 : OUT <= 0;  //12 / 192 = 0
    16'b00001100_11000001 : OUT <= 0;  //12 / 193 = 0
    16'b00001100_11000010 : OUT <= 0;  //12 / 194 = 0
    16'b00001100_11000011 : OUT <= 0;  //12 / 195 = 0
    16'b00001100_11000100 : OUT <= 0;  //12 / 196 = 0
    16'b00001100_11000101 : OUT <= 0;  //12 / 197 = 0
    16'b00001100_11000110 : OUT <= 0;  //12 / 198 = 0
    16'b00001100_11000111 : OUT <= 0;  //12 / 199 = 0
    16'b00001100_11001000 : OUT <= 0;  //12 / 200 = 0
    16'b00001100_11001001 : OUT <= 0;  //12 / 201 = 0
    16'b00001100_11001010 : OUT <= 0;  //12 / 202 = 0
    16'b00001100_11001011 : OUT <= 0;  //12 / 203 = 0
    16'b00001100_11001100 : OUT <= 0;  //12 / 204 = 0
    16'b00001100_11001101 : OUT <= 0;  //12 / 205 = 0
    16'b00001100_11001110 : OUT <= 0;  //12 / 206 = 0
    16'b00001100_11001111 : OUT <= 0;  //12 / 207 = 0
    16'b00001100_11010000 : OUT <= 0;  //12 / 208 = 0
    16'b00001100_11010001 : OUT <= 0;  //12 / 209 = 0
    16'b00001100_11010010 : OUT <= 0;  //12 / 210 = 0
    16'b00001100_11010011 : OUT <= 0;  //12 / 211 = 0
    16'b00001100_11010100 : OUT <= 0;  //12 / 212 = 0
    16'b00001100_11010101 : OUT <= 0;  //12 / 213 = 0
    16'b00001100_11010110 : OUT <= 0;  //12 / 214 = 0
    16'b00001100_11010111 : OUT <= 0;  //12 / 215 = 0
    16'b00001100_11011000 : OUT <= 0;  //12 / 216 = 0
    16'b00001100_11011001 : OUT <= 0;  //12 / 217 = 0
    16'b00001100_11011010 : OUT <= 0;  //12 / 218 = 0
    16'b00001100_11011011 : OUT <= 0;  //12 / 219 = 0
    16'b00001100_11011100 : OUT <= 0;  //12 / 220 = 0
    16'b00001100_11011101 : OUT <= 0;  //12 / 221 = 0
    16'b00001100_11011110 : OUT <= 0;  //12 / 222 = 0
    16'b00001100_11011111 : OUT <= 0;  //12 / 223 = 0
    16'b00001100_11100000 : OUT <= 0;  //12 / 224 = 0
    16'b00001100_11100001 : OUT <= 0;  //12 / 225 = 0
    16'b00001100_11100010 : OUT <= 0;  //12 / 226 = 0
    16'b00001100_11100011 : OUT <= 0;  //12 / 227 = 0
    16'b00001100_11100100 : OUT <= 0;  //12 / 228 = 0
    16'b00001100_11100101 : OUT <= 0;  //12 / 229 = 0
    16'b00001100_11100110 : OUT <= 0;  //12 / 230 = 0
    16'b00001100_11100111 : OUT <= 0;  //12 / 231 = 0
    16'b00001100_11101000 : OUT <= 0;  //12 / 232 = 0
    16'b00001100_11101001 : OUT <= 0;  //12 / 233 = 0
    16'b00001100_11101010 : OUT <= 0;  //12 / 234 = 0
    16'b00001100_11101011 : OUT <= 0;  //12 / 235 = 0
    16'b00001100_11101100 : OUT <= 0;  //12 / 236 = 0
    16'b00001100_11101101 : OUT <= 0;  //12 / 237 = 0
    16'b00001100_11101110 : OUT <= 0;  //12 / 238 = 0
    16'b00001100_11101111 : OUT <= 0;  //12 / 239 = 0
    16'b00001100_11110000 : OUT <= 0;  //12 / 240 = 0
    16'b00001100_11110001 : OUT <= 0;  //12 / 241 = 0
    16'b00001100_11110010 : OUT <= 0;  //12 / 242 = 0
    16'b00001100_11110011 : OUT <= 0;  //12 / 243 = 0
    16'b00001100_11110100 : OUT <= 0;  //12 / 244 = 0
    16'b00001100_11110101 : OUT <= 0;  //12 / 245 = 0
    16'b00001100_11110110 : OUT <= 0;  //12 / 246 = 0
    16'b00001100_11110111 : OUT <= 0;  //12 / 247 = 0
    16'b00001100_11111000 : OUT <= 0;  //12 / 248 = 0
    16'b00001100_11111001 : OUT <= 0;  //12 / 249 = 0
    16'b00001100_11111010 : OUT <= 0;  //12 / 250 = 0
    16'b00001100_11111011 : OUT <= 0;  //12 / 251 = 0
    16'b00001100_11111100 : OUT <= 0;  //12 / 252 = 0
    16'b00001100_11111101 : OUT <= 0;  //12 / 253 = 0
    16'b00001100_11111110 : OUT <= 0;  //12 / 254 = 0
    16'b00001100_11111111 : OUT <= 0;  //12 / 255 = 0
    16'b00001101_00000000 : OUT <= 0;  //13 / 0 = 0
    16'b00001101_00000001 : OUT <= 13;  //13 / 1 = 13
    16'b00001101_00000010 : OUT <= 6;  //13 / 2 = 6
    16'b00001101_00000011 : OUT <= 4;  //13 / 3 = 4
    16'b00001101_00000100 : OUT <= 3;  //13 / 4 = 3
    16'b00001101_00000101 : OUT <= 2;  //13 / 5 = 2
    16'b00001101_00000110 : OUT <= 2;  //13 / 6 = 2
    16'b00001101_00000111 : OUT <= 1;  //13 / 7 = 1
    16'b00001101_00001000 : OUT <= 1;  //13 / 8 = 1
    16'b00001101_00001001 : OUT <= 1;  //13 / 9 = 1
    16'b00001101_00001010 : OUT <= 1;  //13 / 10 = 1
    16'b00001101_00001011 : OUT <= 1;  //13 / 11 = 1
    16'b00001101_00001100 : OUT <= 1;  //13 / 12 = 1
    16'b00001101_00001101 : OUT <= 1;  //13 / 13 = 1
    16'b00001101_00001110 : OUT <= 0;  //13 / 14 = 0
    16'b00001101_00001111 : OUT <= 0;  //13 / 15 = 0
    16'b00001101_00010000 : OUT <= 0;  //13 / 16 = 0
    16'b00001101_00010001 : OUT <= 0;  //13 / 17 = 0
    16'b00001101_00010010 : OUT <= 0;  //13 / 18 = 0
    16'b00001101_00010011 : OUT <= 0;  //13 / 19 = 0
    16'b00001101_00010100 : OUT <= 0;  //13 / 20 = 0
    16'b00001101_00010101 : OUT <= 0;  //13 / 21 = 0
    16'b00001101_00010110 : OUT <= 0;  //13 / 22 = 0
    16'b00001101_00010111 : OUT <= 0;  //13 / 23 = 0
    16'b00001101_00011000 : OUT <= 0;  //13 / 24 = 0
    16'b00001101_00011001 : OUT <= 0;  //13 / 25 = 0
    16'b00001101_00011010 : OUT <= 0;  //13 / 26 = 0
    16'b00001101_00011011 : OUT <= 0;  //13 / 27 = 0
    16'b00001101_00011100 : OUT <= 0;  //13 / 28 = 0
    16'b00001101_00011101 : OUT <= 0;  //13 / 29 = 0
    16'b00001101_00011110 : OUT <= 0;  //13 / 30 = 0
    16'b00001101_00011111 : OUT <= 0;  //13 / 31 = 0
    16'b00001101_00100000 : OUT <= 0;  //13 / 32 = 0
    16'b00001101_00100001 : OUT <= 0;  //13 / 33 = 0
    16'b00001101_00100010 : OUT <= 0;  //13 / 34 = 0
    16'b00001101_00100011 : OUT <= 0;  //13 / 35 = 0
    16'b00001101_00100100 : OUT <= 0;  //13 / 36 = 0
    16'b00001101_00100101 : OUT <= 0;  //13 / 37 = 0
    16'b00001101_00100110 : OUT <= 0;  //13 / 38 = 0
    16'b00001101_00100111 : OUT <= 0;  //13 / 39 = 0
    16'b00001101_00101000 : OUT <= 0;  //13 / 40 = 0
    16'b00001101_00101001 : OUT <= 0;  //13 / 41 = 0
    16'b00001101_00101010 : OUT <= 0;  //13 / 42 = 0
    16'b00001101_00101011 : OUT <= 0;  //13 / 43 = 0
    16'b00001101_00101100 : OUT <= 0;  //13 / 44 = 0
    16'b00001101_00101101 : OUT <= 0;  //13 / 45 = 0
    16'b00001101_00101110 : OUT <= 0;  //13 / 46 = 0
    16'b00001101_00101111 : OUT <= 0;  //13 / 47 = 0
    16'b00001101_00110000 : OUT <= 0;  //13 / 48 = 0
    16'b00001101_00110001 : OUT <= 0;  //13 / 49 = 0
    16'b00001101_00110010 : OUT <= 0;  //13 / 50 = 0
    16'b00001101_00110011 : OUT <= 0;  //13 / 51 = 0
    16'b00001101_00110100 : OUT <= 0;  //13 / 52 = 0
    16'b00001101_00110101 : OUT <= 0;  //13 / 53 = 0
    16'b00001101_00110110 : OUT <= 0;  //13 / 54 = 0
    16'b00001101_00110111 : OUT <= 0;  //13 / 55 = 0
    16'b00001101_00111000 : OUT <= 0;  //13 / 56 = 0
    16'b00001101_00111001 : OUT <= 0;  //13 / 57 = 0
    16'b00001101_00111010 : OUT <= 0;  //13 / 58 = 0
    16'b00001101_00111011 : OUT <= 0;  //13 / 59 = 0
    16'b00001101_00111100 : OUT <= 0;  //13 / 60 = 0
    16'b00001101_00111101 : OUT <= 0;  //13 / 61 = 0
    16'b00001101_00111110 : OUT <= 0;  //13 / 62 = 0
    16'b00001101_00111111 : OUT <= 0;  //13 / 63 = 0
    16'b00001101_01000000 : OUT <= 0;  //13 / 64 = 0
    16'b00001101_01000001 : OUT <= 0;  //13 / 65 = 0
    16'b00001101_01000010 : OUT <= 0;  //13 / 66 = 0
    16'b00001101_01000011 : OUT <= 0;  //13 / 67 = 0
    16'b00001101_01000100 : OUT <= 0;  //13 / 68 = 0
    16'b00001101_01000101 : OUT <= 0;  //13 / 69 = 0
    16'b00001101_01000110 : OUT <= 0;  //13 / 70 = 0
    16'b00001101_01000111 : OUT <= 0;  //13 / 71 = 0
    16'b00001101_01001000 : OUT <= 0;  //13 / 72 = 0
    16'b00001101_01001001 : OUT <= 0;  //13 / 73 = 0
    16'b00001101_01001010 : OUT <= 0;  //13 / 74 = 0
    16'b00001101_01001011 : OUT <= 0;  //13 / 75 = 0
    16'b00001101_01001100 : OUT <= 0;  //13 / 76 = 0
    16'b00001101_01001101 : OUT <= 0;  //13 / 77 = 0
    16'b00001101_01001110 : OUT <= 0;  //13 / 78 = 0
    16'b00001101_01001111 : OUT <= 0;  //13 / 79 = 0
    16'b00001101_01010000 : OUT <= 0;  //13 / 80 = 0
    16'b00001101_01010001 : OUT <= 0;  //13 / 81 = 0
    16'b00001101_01010010 : OUT <= 0;  //13 / 82 = 0
    16'b00001101_01010011 : OUT <= 0;  //13 / 83 = 0
    16'b00001101_01010100 : OUT <= 0;  //13 / 84 = 0
    16'b00001101_01010101 : OUT <= 0;  //13 / 85 = 0
    16'b00001101_01010110 : OUT <= 0;  //13 / 86 = 0
    16'b00001101_01010111 : OUT <= 0;  //13 / 87 = 0
    16'b00001101_01011000 : OUT <= 0;  //13 / 88 = 0
    16'b00001101_01011001 : OUT <= 0;  //13 / 89 = 0
    16'b00001101_01011010 : OUT <= 0;  //13 / 90 = 0
    16'b00001101_01011011 : OUT <= 0;  //13 / 91 = 0
    16'b00001101_01011100 : OUT <= 0;  //13 / 92 = 0
    16'b00001101_01011101 : OUT <= 0;  //13 / 93 = 0
    16'b00001101_01011110 : OUT <= 0;  //13 / 94 = 0
    16'b00001101_01011111 : OUT <= 0;  //13 / 95 = 0
    16'b00001101_01100000 : OUT <= 0;  //13 / 96 = 0
    16'b00001101_01100001 : OUT <= 0;  //13 / 97 = 0
    16'b00001101_01100010 : OUT <= 0;  //13 / 98 = 0
    16'b00001101_01100011 : OUT <= 0;  //13 / 99 = 0
    16'b00001101_01100100 : OUT <= 0;  //13 / 100 = 0
    16'b00001101_01100101 : OUT <= 0;  //13 / 101 = 0
    16'b00001101_01100110 : OUT <= 0;  //13 / 102 = 0
    16'b00001101_01100111 : OUT <= 0;  //13 / 103 = 0
    16'b00001101_01101000 : OUT <= 0;  //13 / 104 = 0
    16'b00001101_01101001 : OUT <= 0;  //13 / 105 = 0
    16'b00001101_01101010 : OUT <= 0;  //13 / 106 = 0
    16'b00001101_01101011 : OUT <= 0;  //13 / 107 = 0
    16'b00001101_01101100 : OUT <= 0;  //13 / 108 = 0
    16'b00001101_01101101 : OUT <= 0;  //13 / 109 = 0
    16'b00001101_01101110 : OUT <= 0;  //13 / 110 = 0
    16'b00001101_01101111 : OUT <= 0;  //13 / 111 = 0
    16'b00001101_01110000 : OUT <= 0;  //13 / 112 = 0
    16'b00001101_01110001 : OUT <= 0;  //13 / 113 = 0
    16'b00001101_01110010 : OUT <= 0;  //13 / 114 = 0
    16'b00001101_01110011 : OUT <= 0;  //13 / 115 = 0
    16'b00001101_01110100 : OUT <= 0;  //13 / 116 = 0
    16'b00001101_01110101 : OUT <= 0;  //13 / 117 = 0
    16'b00001101_01110110 : OUT <= 0;  //13 / 118 = 0
    16'b00001101_01110111 : OUT <= 0;  //13 / 119 = 0
    16'b00001101_01111000 : OUT <= 0;  //13 / 120 = 0
    16'b00001101_01111001 : OUT <= 0;  //13 / 121 = 0
    16'b00001101_01111010 : OUT <= 0;  //13 / 122 = 0
    16'b00001101_01111011 : OUT <= 0;  //13 / 123 = 0
    16'b00001101_01111100 : OUT <= 0;  //13 / 124 = 0
    16'b00001101_01111101 : OUT <= 0;  //13 / 125 = 0
    16'b00001101_01111110 : OUT <= 0;  //13 / 126 = 0
    16'b00001101_01111111 : OUT <= 0;  //13 / 127 = 0
    16'b00001101_10000000 : OUT <= 0;  //13 / 128 = 0
    16'b00001101_10000001 : OUT <= 0;  //13 / 129 = 0
    16'b00001101_10000010 : OUT <= 0;  //13 / 130 = 0
    16'b00001101_10000011 : OUT <= 0;  //13 / 131 = 0
    16'b00001101_10000100 : OUT <= 0;  //13 / 132 = 0
    16'b00001101_10000101 : OUT <= 0;  //13 / 133 = 0
    16'b00001101_10000110 : OUT <= 0;  //13 / 134 = 0
    16'b00001101_10000111 : OUT <= 0;  //13 / 135 = 0
    16'b00001101_10001000 : OUT <= 0;  //13 / 136 = 0
    16'b00001101_10001001 : OUT <= 0;  //13 / 137 = 0
    16'b00001101_10001010 : OUT <= 0;  //13 / 138 = 0
    16'b00001101_10001011 : OUT <= 0;  //13 / 139 = 0
    16'b00001101_10001100 : OUT <= 0;  //13 / 140 = 0
    16'b00001101_10001101 : OUT <= 0;  //13 / 141 = 0
    16'b00001101_10001110 : OUT <= 0;  //13 / 142 = 0
    16'b00001101_10001111 : OUT <= 0;  //13 / 143 = 0
    16'b00001101_10010000 : OUT <= 0;  //13 / 144 = 0
    16'b00001101_10010001 : OUT <= 0;  //13 / 145 = 0
    16'b00001101_10010010 : OUT <= 0;  //13 / 146 = 0
    16'b00001101_10010011 : OUT <= 0;  //13 / 147 = 0
    16'b00001101_10010100 : OUT <= 0;  //13 / 148 = 0
    16'b00001101_10010101 : OUT <= 0;  //13 / 149 = 0
    16'b00001101_10010110 : OUT <= 0;  //13 / 150 = 0
    16'b00001101_10010111 : OUT <= 0;  //13 / 151 = 0
    16'b00001101_10011000 : OUT <= 0;  //13 / 152 = 0
    16'b00001101_10011001 : OUT <= 0;  //13 / 153 = 0
    16'b00001101_10011010 : OUT <= 0;  //13 / 154 = 0
    16'b00001101_10011011 : OUT <= 0;  //13 / 155 = 0
    16'b00001101_10011100 : OUT <= 0;  //13 / 156 = 0
    16'b00001101_10011101 : OUT <= 0;  //13 / 157 = 0
    16'b00001101_10011110 : OUT <= 0;  //13 / 158 = 0
    16'b00001101_10011111 : OUT <= 0;  //13 / 159 = 0
    16'b00001101_10100000 : OUT <= 0;  //13 / 160 = 0
    16'b00001101_10100001 : OUT <= 0;  //13 / 161 = 0
    16'b00001101_10100010 : OUT <= 0;  //13 / 162 = 0
    16'b00001101_10100011 : OUT <= 0;  //13 / 163 = 0
    16'b00001101_10100100 : OUT <= 0;  //13 / 164 = 0
    16'b00001101_10100101 : OUT <= 0;  //13 / 165 = 0
    16'b00001101_10100110 : OUT <= 0;  //13 / 166 = 0
    16'b00001101_10100111 : OUT <= 0;  //13 / 167 = 0
    16'b00001101_10101000 : OUT <= 0;  //13 / 168 = 0
    16'b00001101_10101001 : OUT <= 0;  //13 / 169 = 0
    16'b00001101_10101010 : OUT <= 0;  //13 / 170 = 0
    16'b00001101_10101011 : OUT <= 0;  //13 / 171 = 0
    16'b00001101_10101100 : OUT <= 0;  //13 / 172 = 0
    16'b00001101_10101101 : OUT <= 0;  //13 / 173 = 0
    16'b00001101_10101110 : OUT <= 0;  //13 / 174 = 0
    16'b00001101_10101111 : OUT <= 0;  //13 / 175 = 0
    16'b00001101_10110000 : OUT <= 0;  //13 / 176 = 0
    16'b00001101_10110001 : OUT <= 0;  //13 / 177 = 0
    16'b00001101_10110010 : OUT <= 0;  //13 / 178 = 0
    16'b00001101_10110011 : OUT <= 0;  //13 / 179 = 0
    16'b00001101_10110100 : OUT <= 0;  //13 / 180 = 0
    16'b00001101_10110101 : OUT <= 0;  //13 / 181 = 0
    16'b00001101_10110110 : OUT <= 0;  //13 / 182 = 0
    16'b00001101_10110111 : OUT <= 0;  //13 / 183 = 0
    16'b00001101_10111000 : OUT <= 0;  //13 / 184 = 0
    16'b00001101_10111001 : OUT <= 0;  //13 / 185 = 0
    16'b00001101_10111010 : OUT <= 0;  //13 / 186 = 0
    16'b00001101_10111011 : OUT <= 0;  //13 / 187 = 0
    16'b00001101_10111100 : OUT <= 0;  //13 / 188 = 0
    16'b00001101_10111101 : OUT <= 0;  //13 / 189 = 0
    16'b00001101_10111110 : OUT <= 0;  //13 / 190 = 0
    16'b00001101_10111111 : OUT <= 0;  //13 / 191 = 0
    16'b00001101_11000000 : OUT <= 0;  //13 / 192 = 0
    16'b00001101_11000001 : OUT <= 0;  //13 / 193 = 0
    16'b00001101_11000010 : OUT <= 0;  //13 / 194 = 0
    16'b00001101_11000011 : OUT <= 0;  //13 / 195 = 0
    16'b00001101_11000100 : OUT <= 0;  //13 / 196 = 0
    16'b00001101_11000101 : OUT <= 0;  //13 / 197 = 0
    16'b00001101_11000110 : OUT <= 0;  //13 / 198 = 0
    16'b00001101_11000111 : OUT <= 0;  //13 / 199 = 0
    16'b00001101_11001000 : OUT <= 0;  //13 / 200 = 0
    16'b00001101_11001001 : OUT <= 0;  //13 / 201 = 0
    16'b00001101_11001010 : OUT <= 0;  //13 / 202 = 0
    16'b00001101_11001011 : OUT <= 0;  //13 / 203 = 0
    16'b00001101_11001100 : OUT <= 0;  //13 / 204 = 0
    16'b00001101_11001101 : OUT <= 0;  //13 / 205 = 0
    16'b00001101_11001110 : OUT <= 0;  //13 / 206 = 0
    16'b00001101_11001111 : OUT <= 0;  //13 / 207 = 0
    16'b00001101_11010000 : OUT <= 0;  //13 / 208 = 0
    16'b00001101_11010001 : OUT <= 0;  //13 / 209 = 0
    16'b00001101_11010010 : OUT <= 0;  //13 / 210 = 0
    16'b00001101_11010011 : OUT <= 0;  //13 / 211 = 0
    16'b00001101_11010100 : OUT <= 0;  //13 / 212 = 0
    16'b00001101_11010101 : OUT <= 0;  //13 / 213 = 0
    16'b00001101_11010110 : OUT <= 0;  //13 / 214 = 0
    16'b00001101_11010111 : OUT <= 0;  //13 / 215 = 0
    16'b00001101_11011000 : OUT <= 0;  //13 / 216 = 0
    16'b00001101_11011001 : OUT <= 0;  //13 / 217 = 0
    16'b00001101_11011010 : OUT <= 0;  //13 / 218 = 0
    16'b00001101_11011011 : OUT <= 0;  //13 / 219 = 0
    16'b00001101_11011100 : OUT <= 0;  //13 / 220 = 0
    16'b00001101_11011101 : OUT <= 0;  //13 / 221 = 0
    16'b00001101_11011110 : OUT <= 0;  //13 / 222 = 0
    16'b00001101_11011111 : OUT <= 0;  //13 / 223 = 0
    16'b00001101_11100000 : OUT <= 0;  //13 / 224 = 0
    16'b00001101_11100001 : OUT <= 0;  //13 / 225 = 0
    16'b00001101_11100010 : OUT <= 0;  //13 / 226 = 0
    16'b00001101_11100011 : OUT <= 0;  //13 / 227 = 0
    16'b00001101_11100100 : OUT <= 0;  //13 / 228 = 0
    16'b00001101_11100101 : OUT <= 0;  //13 / 229 = 0
    16'b00001101_11100110 : OUT <= 0;  //13 / 230 = 0
    16'b00001101_11100111 : OUT <= 0;  //13 / 231 = 0
    16'b00001101_11101000 : OUT <= 0;  //13 / 232 = 0
    16'b00001101_11101001 : OUT <= 0;  //13 / 233 = 0
    16'b00001101_11101010 : OUT <= 0;  //13 / 234 = 0
    16'b00001101_11101011 : OUT <= 0;  //13 / 235 = 0
    16'b00001101_11101100 : OUT <= 0;  //13 / 236 = 0
    16'b00001101_11101101 : OUT <= 0;  //13 / 237 = 0
    16'b00001101_11101110 : OUT <= 0;  //13 / 238 = 0
    16'b00001101_11101111 : OUT <= 0;  //13 / 239 = 0
    16'b00001101_11110000 : OUT <= 0;  //13 / 240 = 0
    16'b00001101_11110001 : OUT <= 0;  //13 / 241 = 0
    16'b00001101_11110010 : OUT <= 0;  //13 / 242 = 0
    16'b00001101_11110011 : OUT <= 0;  //13 / 243 = 0
    16'b00001101_11110100 : OUT <= 0;  //13 / 244 = 0
    16'b00001101_11110101 : OUT <= 0;  //13 / 245 = 0
    16'b00001101_11110110 : OUT <= 0;  //13 / 246 = 0
    16'b00001101_11110111 : OUT <= 0;  //13 / 247 = 0
    16'b00001101_11111000 : OUT <= 0;  //13 / 248 = 0
    16'b00001101_11111001 : OUT <= 0;  //13 / 249 = 0
    16'b00001101_11111010 : OUT <= 0;  //13 / 250 = 0
    16'b00001101_11111011 : OUT <= 0;  //13 / 251 = 0
    16'b00001101_11111100 : OUT <= 0;  //13 / 252 = 0
    16'b00001101_11111101 : OUT <= 0;  //13 / 253 = 0
    16'b00001101_11111110 : OUT <= 0;  //13 / 254 = 0
    16'b00001101_11111111 : OUT <= 0;  //13 / 255 = 0
    16'b00001110_00000000 : OUT <= 0;  //14 / 0 = 0
    16'b00001110_00000001 : OUT <= 14;  //14 / 1 = 14
    16'b00001110_00000010 : OUT <= 7;  //14 / 2 = 7
    16'b00001110_00000011 : OUT <= 4;  //14 / 3 = 4
    16'b00001110_00000100 : OUT <= 3;  //14 / 4 = 3
    16'b00001110_00000101 : OUT <= 2;  //14 / 5 = 2
    16'b00001110_00000110 : OUT <= 2;  //14 / 6 = 2
    16'b00001110_00000111 : OUT <= 2;  //14 / 7 = 2
    16'b00001110_00001000 : OUT <= 1;  //14 / 8 = 1
    16'b00001110_00001001 : OUT <= 1;  //14 / 9 = 1
    16'b00001110_00001010 : OUT <= 1;  //14 / 10 = 1
    16'b00001110_00001011 : OUT <= 1;  //14 / 11 = 1
    16'b00001110_00001100 : OUT <= 1;  //14 / 12 = 1
    16'b00001110_00001101 : OUT <= 1;  //14 / 13 = 1
    16'b00001110_00001110 : OUT <= 1;  //14 / 14 = 1
    16'b00001110_00001111 : OUT <= 0;  //14 / 15 = 0
    16'b00001110_00010000 : OUT <= 0;  //14 / 16 = 0
    16'b00001110_00010001 : OUT <= 0;  //14 / 17 = 0
    16'b00001110_00010010 : OUT <= 0;  //14 / 18 = 0
    16'b00001110_00010011 : OUT <= 0;  //14 / 19 = 0
    16'b00001110_00010100 : OUT <= 0;  //14 / 20 = 0
    16'b00001110_00010101 : OUT <= 0;  //14 / 21 = 0
    16'b00001110_00010110 : OUT <= 0;  //14 / 22 = 0
    16'b00001110_00010111 : OUT <= 0;  //14 / 23 = 0
    16'b00001110_00011000 : OUT <= 0;  //14 / 24 = 0
    16'b00001110_00011001 : OUT <= 0;  //14 / 25 = 0
    16'b00001110_00011010 : OUT <= 0;  //14 / 26 = 0
    16'b00001110_00011011 : OUT <= 0;  //14 / 27 = 0
    16'b00001110_00011100 : OUT <= 0;  //14 / 28 = 0
    16'b00001110_00011101 : OUT <= 0;  //14 / 29 = 0
    16'b00001110_00011110 : OUT <= 0;  //14 / 30 = 0
    16'b00001110_00011111 : OUT <= 0;  //14 / 31 = 0
    16'b00001110_00100000 : OUT <= 0;  //14 / 32 = 0
    16'b00001110_00100001 : OUT <= 0;  //14 / 33 = 0
    16'b00001110_00100010 : OUT <= 0;  //14 / 34 = 0
    16'b00001110_00100011 : OUT <= 0;  //14 / 35 = 0
    16'b00001110_00100100 : OUT <= 0;  //14 / 36 = 0
    16'b00001110_00100101 : OUT <= 0;  //14 / 37 = 0
    16'b00001110_00100110 : OUT <= 0;  //14 / 38 = 0
    16'b00001110_00100111 : OUT <= 0;  //14 / 39 = 0
    16'b00001110_00101000 : OUT <= 0;  //14 / 40 = 0
    16'b00001110_00101001 : OUT <= 0;  //14 / 41 = 0
    16'b00001110_00101010 : OUT <= 0;  //14 / 42 = 0
    16'b00001110_00101011 : OUT <= 0;  //14 / 43 = 0
    16'b00001110_00101100 : OUT <= 0;  //14 / 44 = 0
    16'b00001110_00101101 : OUT <= 0;  //14 / 45 = 0
    16'b00001110_00101110 : OUT <= 0;  //14 / 46 = 0
    16'b00001110_00101111 : OUT <= 0;  //14 / 47 = 0
    16'b00001110_00110000 : OUT <= 0;  //14 / 48 = 0
    16'b00001110_00110001 : OUT <= 0;  //14 / 49 = 0
    16'b00001110_00110010 : OUT <= 0;  //14 / 50 = 0
    16'b00001110_00110011 : OUT <= 0;  //14 / 51 = 0
    16'b00001110_00110100 : OUT <= 0;  //14 / 52 = 0
    16'b00001110_00110101 : OUT <= 0;  //14 / 53 = 0
    16'b00001110_00110110 : OUT <= 0;  //14 / 54 = 0
    16'b00001110_00110111 : OUT <= 0;  //14 / 55 = 0
    16'b00001110_00111000 : OUT <= 0;  //14 / 56 = 0
    16'b00001110_00111001 : OUT <= 0;  //14 / 57 = 0
    16'b00001110_00111010 : OUT <= 0;  //14 / 58 = 0
    16'b00001110_00111011 : OUT <= 0;  //14 / 59 = 0
    16'b00001110_00111100 : OUT <= 0;  //14 / 60 = 0
    16'b00001110_00111101 : OUT <= 0;  //14 / 61 = 0
    16'b00001110_00111110 : OUT <= 0;  //14 / 62 = 0
    16'b00001110_00111111 : OUT <= 0;  //14 / 63 = 0
    16'b00001110_01000000 : OUT <= 0;  //14 / 64 = 0
    16'b00001110_01000001 : OUT <= 0;  //14 / 65 = 0
    16'b00001110_01000010 : OUT <= 0;  //14 / 66 = 0
    16'b00001110_01000011 : OUT <= 0;  //14 / 67 = 0
    16'b00001110_01000100 : OUT <= 0;  //14 / 68 = 0
    16'b00001110_01000101 : OUT <= 0;  //14 / 69 = 0
    16'b00001110_01000110 : OUT <= 0;  //14 / 70 = 0
    16'b00001110_01000111 : OUT <= 0;  //14 / 71 = 0
    16'b00001110_01001000 : OUT <= 0;  //14 / 72 = 0
    16'b00001110_01001001 : OUT <= 0;  //14 / 73 = 0
    16'b00001110_01001010 : OUT <= 0;  //14 / 74 = 0
    16'b00001110_01001011 : OUT <= 0;  //14 / 75 = 0
    16'b00001110_01001100 : OUT <= 0;  //14 / 76 = 0
    16'b00001110_01001101 : OUT <= 0;  //14 / 77 = 0
    16'b00001110_01001110 : OUT <= 0;  //14 / 78 = 0
    16'b00001110_01001111 : OUT <= 0;  //14 / 79 = 0
    16'b00001110_01010000 : OUT <= 0;  //14 / 80 = 0
    16'b00001110_01010001 : OUT <= 0;  //14 / 81 = 0
    16'b00001110_01010010 : OUT <= 0;  //14 / 82 = 0
    16'b00001110_01010011 : OUT <= 0;  //14 / 83 = 0
    16'b00001110_01010100 : OUT <= 0;  //14 / 84 = 0
    16'b00001110_01010101 : OUT <= 0;  //14 / 85 = 0
    16'b00001110_01010110 : OUT <= 0;  //14 / 86 = 0
    16'b00001110_01010111 : OUT <= 0;  //14 / 87 = 0
    16'b00001110_01011000 : OUT <= 0;  //14 / 88 = 0
    16'b00001110_01011001 : OUT <= 0;  //14 / 89 = 0
    16'b00001110_01011010 : OUT <= 0;  //14 / 90 = 0
    16'b00001110_01011011 : OUT <= 0;  //14 / 91 = 0
    16'b00001110_01011100 : OUT <= 0;  //14 / 92 = 0
    16'b00001110_01011101 : OUT <= 0;  //14 / 93 = 0
    16'b00001110_01011110 : OUT <= 0;  //14 / 94 = 0
    16'b00001110_01011111 : OUT <= 0;  //14 / 95 = 0
    16'b00001110_01100000 : OUT <= 0;  //14 / 96 = 0
    16'b00001110_01100001 : OUT <= 0;  //14 / 97 = 0
    16'b00001110_01100010 : OUT <= 0;  //14 / 98 = 0
    16'b00001110_01100011 : OUT <= 0;  //14 / 99 = 0
    16'b00001110_01100100 : OUT <= 0;  //14 / 100 = 0
    16'b00001110_01100101 : OUT <= 0;  //14 / 101 = 0
    16'b00001110_01100110 : OUT <= 0;  //14 / 102 = 0
    16'b00001110_01100111 : OUT <= 0;  //14 / 103 = 0
    16'b00001110_01101000 : OUT <= 0;  //14 / 104 = 0
    16'b00001110_01101001 : OUT <= 0;  //14 / 105 = 0
    16'b00001110_01101010 : OUT <= 0;  //14 / 106 = 0
    16'b00001110_01101011 : OUT <= 0;  //14 / 107 = 0
    16'b00001110_01101100 : OUT <= 0;  //14 / 108 = 0
    16'b00001110_01101101 : OUT <= 0;  //14 / 109 = 0
    16'b00001110_01101110 : OUT <= 0;  //14 / 110 = 0
    16'b00001110_01101111 : OUT <= 0;  //14 / 111 = 0
    16'b00001110_01110000 : OUT <= 0;  //14 / 112 = 0
    16'b00001110_01110001 : OUT <= 0;  //14 / 113 = 0
    16'b00001110_01110010 : OUT <= 0;  //14 / 114 = 0
    16'b00001110_01110011 : OUT <= 0;  //14 / 115 = 0
    16'b00001110_01110100 : OUT <= 0;  //14 / 116 = 0
    16'b00001110_01110101 : OUT <= 0;  //14 / 117 = 0
    16'b00001110_01110110 : OUT <= 0;  //14 / 118 = 0
    16'b00001110_01110111 : OUT <= 0;  //14 / 119 = 0
    16'b00001110_01111000 : OUT <= 0;  //14 / 120 = 0
    16'b00001110_01111001 : OUT <= 0;  //14 / 121 = 0
    16'b00001110_01111010 : OUT <= 0;  //14 / 122 = 0
    16'b00001110_01111011 : OUT <= 0;  //14 / 123 = 0
    16'b00001110_01111100 : OUT <= 0;  //14 / 124 = 0
    16'b00001110_01111101 : OUT <= 0;  //14 / 125 = 0
    16'b00001110_01111110 : OUT <= 0;  //14 / 126 = 0
    16'b00001110_01111111 : OUT <= 0;  //14 / 127 = 0
    16'b00001110_10000000 : OUT <= 0;  //14 / 128 = 0
    16'b00001110_10000001 : OUT <= 0;  //14 / 129 = 0
    16'b00001110_10000010 : OUT <= 0;  //14 / 130 = 0
    16'b00001110_10000011 : OUT <= 0;  //14 / 131 = 0
    16'b00001110_10000100 : OUT <= 0;  //14 / 132 = 0
    16'b00001110_10000101 : OUT <= 0;  //14 / 133 = 0
    16'b00001110_10000110 : OUT <= 0;  //14 / 134 = 0
    16'b00001110_10000111 : OUT <= 0;  //14 / 135 = 0
    16'b00001110_10001000 : OUT <= 0;  //14 / 136 = 0
    16'b00001110_10001001 : OUT <= 0;  //14 / 137 = 0
    16'b00001110_10001010 : OUT <= 0;  //14 / 138 = 0
    16'b00001110_10001011 : OUT <= 0;  //14 / 139 = 0
    16'b00001110_10001100 : OUT <= 0;  //14 / 140 = 0
    16'b00001110_10001101 : OUT <= 0;  //14 / 141 = 0
    16'b00001110_10001110 : OUT <= 0;  //14 / 142 = 0
    16'b00001110_10001111 : OUT <= 0;  //14 / 143 = 0
    16'b00001110_10010000 : OUT <= 0;  //14 / 144 = 0
    16'b00001110_10010001 : OUT <= 0;  //14 / 145 = 0
    16'b00001110_10010010 : OUT <= 0;  //14 / 146 = 0
    16'b00001110_10010011 : OUT <= 0;  //14 / 147 = 0
    16'b00001110_10010100 : OUT <= 0;  //14 / 148 = 0
    16'b00001110_10010101 : OUT <= 0;  //14 / 149 = 0
    16'b00001110_10010110 : OUT <= 0;  //14 / 150 = 0
    16'b00001110_10010111 : OUT <= 0;  //14 / 151 = 0
    16'b00001110_10011000 : OUT <= 0;  //14 / 152 = 0
    16'b00001110_10011001 : OUT <= 0;  //14 / 153 = 0
    16'b00001110_10011010 : OUT <= 0;  //14 / 154 = 0
    16'b00001110_10011011 : OUT <= 0;  //14 / 155 = 0
    16'b00001110_10011100 : OUT <= 0;  //14 / 156 = 0
    16'b00001110_10011101 : OUT <= 0;  //14 / 157 = 0
    16'b00001110_10011110 : OUT <= 0;  //14 / 158 = 0
    16'b00001110_10011111 : OUT <= 0;  //14 / 159 = 0
    16'b00001110_10100000 : OUT <= 0;  //14 / 160 = 0
    16'b00001110_10100001 : OUT <= 0;  //14 / 161 = 0
    16'b00001110_10100010 : OUT <= 0;  //14 / 162 = 0
    16'b00001110_10100011 : OUT <= 0;  //14 / 163 = 0
    16'b00001110_10100100 : OUT <= 0;  //14 / 164 = 0
    16'b00001110_10100101 : OUT <= 0;  //14 / 165 = 0
    16'b00001110_10100110 : OUT <= 0;  //14 / 166 = 0
    16'b00001110_10100111 : OUT <= 0;  //14 / 167 = 0
    16'b00001110_10101000 : OUT <= 0;  //14 / 168 = 0
    16'b00001110_10101001 : OUT <= 0;  //14 / 169 = 0
    16'b00001110_10101010 : OUT <= 0;  //14 / 170 = 0
    16'b00001110_10101011 : OUT <= 0;  //14 / 171 = 0
    16'b00001110_10101100 : OUT <= 0;  //14 / 172 = 0
    16'b00001110_10101101 : OUT <= 0;  //14 / 173 = 0
    16'b00001110_10101110 : OUT <= 0;  //14 / 174 = 0
    16'b00001110_10101111 : OUT <= 0;  //14 / 175 = 0
    16'b00001110_10110000 : OUT <= 0;  //14 / 176 = 0
    16'b00001110_10110001 : OUT <= 0;  //14 / 177 = 0
    16'b00001110_10110010 : OUT <= 0;  //14 / 178 = 0
    16'b00001110_10110011 : OUT <= 0;  //14 / 179 = 0
    16'b00001110_10110100 : OUT <= 0;  //14 / 180 = 0
    16'b00001110_10110101 : OUT <= 0;  //14 / 181 = 0
    16'b00001110_10110110 : OUT <= 0;  //14 / 182 = 0
    16'b00001110_10110111 : OUT <= 0;  //14 / 183 = 0
    16'b00001110_10111000 : OUT <= 0;  //14 / 184 = 0
    16'b00001110_10111001 : OUT <= 0;  //14 / 185 = 0
    16'b00001110_10111010 : OUT <= 0;  //14 / 186 = 0
    16'b00001110_10111011 : OUT <= 0;  //14 / 187 = 0
    16'b00001110_10111100 : OUT <= 0;  //14 / 188 = 0
    16'b00001110_10111101 : OUT <= 0;  //14 / 189 = 0
    16'b00001110_10111110 : OUT <= 0;  //14 / 190 = 0
    16'b00001110_10111111 : OUT <= 0;  //14 / 191 = 0
    16'b00001110_11000000 : OUT <= 0;  //14 / 192 = 0
    16'b00001110_11000001 : OUT <= 0;  //14 / 193 = 0
    16'b00001110_11000010 : OUT <= 0;  //14 / 194 = 0
    16'b00001110_11000011 : OUT <= 0;  //14 / 195 = 0
    16'b00001110_11000100 : OUT <= 0;  //14 / 196 = 0
    16'b00001110_11000101 : OUT <= 0;  //14 / 197 = 0
    16'b00001110_11000110 : OUT <= 0;  //14 / 198 = 0
    16'b00001110_11000111 : OUT <= 0;  //14 / 199 = 0
    16'b00001110_11001000 : OUT <= 0;  //14 / 200 = 0
    16'b00001110_11001001 : OUT <= 0;  //14 / 201 = 0
    16'b00001110_11001010 : OUT <= 0;  //14 / 202 = 0
    16'b00001110_11001011 : OUT <= 0;  //14 / 203 = 0
    16'b00001110_11001100 : OUT <= 0;  //14 / 204 = 0
    16'b00001110_11001101 : OUT <= 0;  //14 / 205 = 0
    16'b00001110_11001110 : OUT <= 0;  //14 / 206 = 0
    16'b00001110_11001111 : OUT <= 0;  //14 / 207 = 0
    16'b00001110_11010000 : OUT <= 0;  //14 / 208 = 0
    16'b00001110_11010001 : OUT <= 0;  //14 / 209 = 0
    16'b00001110_11010010 : OUT <= 0;  //14 / 210 = 0
    16'b00001110_11010011 : OUT <= 0;  //14 / 211 = 0
    16'b00001110_11010100 : OUT <= 0;  //14 / 212 = 0
    16'b00001110_11010101 : OUT <= 0;  //14 / 213 = 0
    16'b00001110_11010110 : OUT <= 0;  //14 / 214 = 0
    16'b00001110_11010111 : OUT <= 0;  //14 / 215 = 0
    16'b00001110_11011000 : OUT <= 0;  //14 / 216 = 0
    16'b00001110_11011001 : OUT <= 0;  //14 / 217 = 0
    16'b00001110_11011010 : OUT <= 0;  //14 / 218 = 0
    16'b00001110_11011011 : OUT <= 0;  //14 / 219 = 0
    16'b00001110_11011100 : OUT <= 0;  //14 / 220 = 0
    16'b00001110_11011101 : OUT <= 0;  //14 / 221 = 0
    16'b00001110_11011110 : OUT <= 0;  //14 / 222 = 0
    16'b00001110_11011111 : OUT <= 0;  //14 / 223 = 0
    16'b00001110_11100000 : OUT <= 0;  //14 / 224 = 0
    16'b00001110_11100001 : OUT <= 0;  //14 / 225 = 0
    16'b00001110_11100010 : OUT <= 0;  //14 / 226 = 0
    16'b00001110_11100011 : OUT <= 0;  //14 / 227 = 0
    16'b00001110_11100100 : OUT <= 0;  //14 / 228 = 0
    16'b00001110_11100101 : OUT <= 0;  //14 / 229 = 0
    16'b00001110_11100110 : OUT <= 0;  //14 / 230 = 0
    16'b00001110_11100111 : OUT <= 0;  //14 / 231 = 0
    16'b00001110_11101000 : OUT <= 0;  //14 / 232 = 0
    16'b00001110_11101001 : OUT <= 0;  //14 / 233 = 0
    16'b00001110_11101010 : OUT <= 0;  //14 / 234 = 0
    16'b00001110_11101011 : OUT <= 0;  //14 / 235 = 0
    16'b00001110_11101100 : OUT <= 0;  //14 / 236 = 0
    16'b00001110_11101101 : OUT <= 0;  //14 / 237 = 0
    16'b00001110_11101110 : OUT <= 0;  //14 / 238 = 0
    16'b00001110_11101111 : OUT <= 0;  //14 / 239 = 0
    16'b00001110_11110000 : OUT <= 0;  //14 / 240 = 0
    16'b00001110_11110001 : OUT <= 0;  //14 / 241 = 0
    16'b00001110_11110010 : OUT <= 0;  //14 / 242 = 0
    16'b00001110_11110011 : OUT <= 0;  //14 / 243 = 0
    16'b00001110_11110100 : OUT <= 0;  //14 / 244 = 0
    16'b00001110_11110101 : OUT <= 0;  //14 / 245 = 0
    16'b00001110_11110110 : OUT <= 0;  //14 / 246 = 0
    16'b00001110_11110111 : OUT <= 0;  //14 / 247 = 0
    16'b00001110_11111000 : OUT <= 0;  //14 / 248 = 0
    16'b00001110_11111001 : OUT <= 0;  //14 / 249 = 0
    16'b00001110_11111010 : OUT <= 0;  //14 / 250 = 0
    16'b00001110_11111011 : OUT <= 0;  //14 / 251 = 0
    16'b00001110_11111100 : OUT <= 0;  //14 / 252 = 0
    16'b00001110_11111101 : OUT <= 0;  //14 / 253 = 0
    16'b00001110_11111110 : OUT <= 0;  //14 / 254 = 0
    16'b00001110_11111111 : OUT <= 0;  //14 / 255 = 0
    16'b00001111_00000000 : OUT <= 0;  //15 / 0 = 0
    16'b00001111_00000001 : OUT <= 15;  //15 / 1 = 15
    16'b00001111_00000010 : OUT <= 7;  //15 / 2 = 7
    16'b00001111_00000011 : OUT <= 5;  //15 / 3 = 5
    16'b00001111_00000100 : OUT <= 3;  //15 / 4 = 3
    16'b00001111_00000101 : OUT <= 3;  //15 / 5 = 3
    16'b00001111_00000110 : OUT <= 2;  //15 / 6 = 2
    16'b00001111_00000111 : OUT <= 2;  //15 / 7 = 2
    16'b00001111_00001000 : OUT <= 1;  //15 / 8 = 1
    16'b00001111_00001001 : OUT <= 1;  //15 / 9 = 1
    16'b00001111_00001010 : OUT <= 1;  //15 / 10 = 1
    16'b00001111_00001011 : OUT <= 1;  //15 / 11 = 1
    16'b00001111_00001100 : OUT <= 1;  //15 / 12 = 1
    16'b00001111_00001101 : OUT <= 1;  //15 / 13 = 1
    16'b00001111_00001110 : OUT <= 1;  //15 / 14 = 1
    16'b00001111_00001111 : OUT <= 1;  //15 / 15 = 1
    16'b00001111_00010000 : OUT <= 0;  //15 / 16 = 0
    16'b00001111_00010001 : OUT <= 0;  //15 / 17 = 0
    16'b00001111_00010010 : OUT <= 0;  //15 / 18 = 0
    16'b00001111_00010011 : OUT <= 0;  //15 / 19 = 0
    16'b00001111_00010100 : OUT <= 0;  //15 / 20 = 0
    16'b00001111_00010101 : OUT <= 0;  //15 / 21 = 0
    16'b00001111_00010110 : OUT <= 0;  //15 / 22 = 0
    16'b00001111_00010111 : OUT <= 0;  //15 / 23 = 0
    16'b00001111_00011000 : OUT <= 0;  //15 / 24 = 0
    16'b00001111_00011001 : OUT <= 0;  //15 / 25 = 0
    16'b00001111_00011010 : OUT <= 0;  //15 / 26 = 0
    16'b00001111_00011011 : OUT <= 0;  //15 / 27 = 0
    16'b00001111_00011100 : OUT <= 0;  //15 / 28 = 0
    16'b00001111_00011101 : OUT <= 0;  //15 / 29 = 0
    16'b00001111_00011110 : OUT <= 0;  //15 / 30 = 0
    16'b00001111_00011111 : OUT <= 0;  //15 / 31 = 0
    16'b00001111_00100000 : OUT <= 0;  //15 / 32 = 0
    16'b00001111_00100001 : OUT <= 0;  //15 / 33 = 0
    16'b00001111_00100010 : OUT <= 0;  //15 / 34 = 0
    16'b00001111_00100011 : OUT <= 0;  //15 / 35 = 0
    16'b00001111_00100100 : OUT <= 0;  //15 / 36 = 0
    16'b00001111_00100101 : OUT <= 0;  //15 / 37 = 0
    16'b00001111_00100110 : OUT <= 0;  //15 / 38 = 0
    16'b00001111_00100111 : OUT <= 0;  //15 / 39 = 0
    16'b00001111_00101000 : OUT <= 0;  //15 / 40 = 0
    16'b00001111_00101001 : OUT <= 0;  //15 / 41 = 0
    16'b00001111_00101010 : OUT <= 0;  //15 / 42 = 0
    16'b00001111_00101011 : OUT <= 0;  //15 / 43 = 0
    16'b00001111_00101100 : OUT <= 0;  //15 / 44 = 0
    16'b00001111_00101101 : OUT <= 0;  //15 / 45 = 0
    16'b00001111_00101110 : OUT <= 0;  //15 / 46 = 0
    16'b00001111_00101111 : OUT <= 0;  //15 / 47 = 0
    16'b00001111_00110000 : OUT <= 0;  //15 / 48 = 0
    16'b00001111_00110001 : OUT <= 0;  //15 / 49 = 0
    16'b00001111_00110010 : OUT <= 0;  //15 / 50 = 0
    16'b00001111_00110011 : OUT <= 0;  //15 / 51 = 0
    16'b00001111_00110100 : OUT <= 0;  //15 / 52 = 0
    16'b00001111_00110101 : OUT <= 0;  //15 / 53 = 0
    16'b00001111_00110110 : OUT <= 0;  //15 / 54 = 0
    16'b00001111_00110111 : OUT <= 0;  //15 / 55 = 0
    16'b00001111_00111000 : OUT <= 0;  //15 / 56 = 0
    16'b00001111_00111001 : OUT <= 0;  //15 / 57 = 0
    16'b00001111_00111010 : OUT <= 0;  //15 / 58 = 0
    16'b00001111_00111011 : OUT <= 0;  //15 / 59 = 0
    16'b00001111_00111100 : OUT <= 0;  //15 / 60 = 0
    16'b00001111_00111101 : OUT <= 0;  //15 / 61 = 0
    16'b00001111_00111110 : OUT <= 0;  //15 / 62 = 0
    16'b00001111_00111111 : OUT <= 0;  //15 / 63 = 0
    16'b00001111_01000000 : OUT <= 0;  //15 / 64 = 0
    16'b00001111_01000001 : OUT <= 0;  //15 / 65 = 0
    16'b00001111_01000010 : OUT <= 0;  //15 / 66 = 0
    16'b00001111_01000011 : OUT <= 0;  //15 / 67 = 0
    16'b00001111_01000100 : OUT <= 0;  //15 / 68 = 0
    16'b00001111_01000101 : OUT <= 0;  //15 / 69 = 0
    16'b00001111_01000110 : OUT <= 0;  //15 / 70 = 0
    16'b00001111_01000111 : OUT <= 0;  //15 / 71 = 0
    16'b00001111_01001000 : OUT <= 0;  //15 / 72 = 0
    16'b00001111_01001001 : OUT <= 0;  //15 / 73 = 0
    16'b00001111_01001010 : OUT <= 0;  //15 / 74 = 0
    16'b00001111_01001011 : OUT <= 0;  //15 / 75 = 0
    16'b00001111_01001100 : OUT <= 0;  //15 / 76 = 0
    16'b00001111_01001101 : OUT <= 0;  //15 / 77 = 0
    16'b00001111_01001110 : OUT <= 0;  //15 / 78 = 0
    16'b00001111_01001111 : OUT <= 0;  //15 / 79 = 0
    16'b00001111_01010000 : OUT <= 0;  //15 / 80 = 0
    16'b00001111_01010001 : OUT <= 0;  //15 / 81 = 0
    16'b00001111_01010010 : OUT <= 0;  //15 / 82 = 0
    16'b00001111_01010011 : OUT <= 0;  //15 / 83 = 0
    16'b00001111_01010100 : OUT <= 0;  //15 / 84 = 0
    16'b00001111_01010101 : OUT <= 0;  //15 / 85 = 0
    16'b00001111_01010110 : OUT <= 0;  //15 / 86 = 0
    16'b00001111_01010111 : OUT <= 0;  //15 / 87 = 0
    16'b00001111_01011000 : OUT <= 0;  //15 / 88 = 0
    16'b00001111_01011001 : OUT <= 0;  //15 / 89 = 0
    16'b00001111_01011010 : OUT <= 0;  //15 / 90 = 0
    16'b00001111_01011011 : OUT <= 0;  //15 / 91 = 0
    16'b00001111_01011100 : OUT <= 0;  //15 / 92 = 0
    16'b00001111_01011101 : OUT <= 0;  //15 / 93 = 0
    16'b00001111_01011110 : OUT <= 0;  //15 / 94 = 0
    16'b00001111_01011111 : OUT <= 0;  //15 / 95 = 0
    16'b00001111_01100000 : OUT <= 0;  //15 / 96 = 0
    16'b00001111_01100001 : OUT <= 0;  //15 / 97 = 0
    16'b00001111_01100010 : OUT <= 0;  //15 / 98 = 0
    16'b00001111_01100011 : OUT <= 0;  //15 / 99 = 0
    16'b00001111_01100100 : OUT <= 0;  //15 / 100 = 0
    16'b00001111_01100101 : OUT <= 0;  //15 / 101 = 0
    16'b00001111_01100110 : OUT <= 0;  //15 / 102 = 0
    16'b00001111_01100111 : OUT <= 0;  //15 / 103 = 0
    16'b00001111_01101000 : OUT <= 0;  //15 / 104 = 0
    16'b00001111_01101001 : OUT <= 0;  //15 / 105 = 0
    16'b00001111_01101010 : OUT <= 0;  //15 / 106 = 0
    16'b00001111_01101011 : OUT <= 0;  //15 / 107 = 0
    16'b00001111_01101100 : OUT <= 0;  //15 / 108 = 0
    16'b00001111_01101101 : OUT <= 0;  //15 / 109 = 0
    16'b00001111_01101110 : OUT <= 0;  //15 / 110 = 0
    16'b00001111_01101111 : OUT <= 0;  //15 / 111 = 0
    16'b00001111_01110000 : OUT <= 0;  //15 / 112 = 0
    16'b00001111_01110001 : OUT <= 0;  //15 / 113 = 0
    16'b00001111_01110010 : OUT <= 0;  //15 / 114 = 0
    16'b00001111_01110011 : OUT <= 0;  //15 / 115 = 0
    16'b00001111_01110100 : OUT <= 0;  //15 / 116 = 0
    16'b00001111_01110101 : OUT <= 0;  //15 / 117 = 0
    16'b00001111_01110110 : OUT <= 0;  //15 / 118 = 0
    16'b00001111_01110111 : OUT <= 0;  //15 / 119 = 0
    16'b00001111_01111000 : OUT <= 0;  //15 / 120 = 0
    16'b00001111_01111001 : OUT <= 0;  //15 / 121 = 0
    16'b00001111_01111010 : OUT <= 0;  //15 / 122 = 0
    16'b00001111_01111011 : OUT <= 0;  //15 / 123 = 0
    16'b00001111_01111100 : OUT <= 0;  //15 / 124 = 0
    16'b00001111_01111101 : OUT <= 0;  //15 / 125 = 0
    16'b00001111_01111110 : OUT <= 0;  //15 / 126 = 0
    16'b00001111_01111111 : OUT <= 0;  //15 / 127 = 0
    16'b00001111_10000000 : OUT <= 0;  //15 / 128 = 0
    16'b00001111_10000001 : OUT <= 0;  //15 / 129 = 0
    16'b00001111_10000010 : OUT <= 0;  //15 / 130 = 0
    16'b00001111_10000011 : OUT <= 0;  //15 / 131 = 0
    16'b00001111_10000100 : OUT <= 0;  //15 / 132 = 0
    16'b00001111_10000101 : OUT <= 0;  //15 / 133 = 0
    16'b00001111_10000110 : OUT <= 0;  //15 / 134 = 0
    16'b00001111_10000111 : OUT <= 0;  //15 / 135 = 0
    16'b00001111_10001000 : OUT <= 0;  //15 / 136 = 0
    16'b00001111_10001001 : OUT <= 0;  //15 / 137 = 0
    16'b00001111_10001010 : OUT <= 0;  //15 / 138 = 0
    16'b00001111_10001011 : OUT <= 0;  //15 / 139 = 0
    16'b00001111_10001100 : OUT <= 0;  //15 / 140 = 0
    16'b00001111_10001101 : OUT <= 0;  //15 / 141 = 0
    16'b00001111_10001110 : OUT <= 0;  //15 / 142 = 0
    16'b00001111_10001111 : OUT <= 0;  //15 / 143 = 0
    16'b00001111_10010000 : OUT <= 0;  //15 / 144 = 0
    16'b00001111_10010001 : OUT <= 0;  //15 / 145 = 0
    16'b00001111_10010010 : OUT <= 0;  //15 / 146 = 0
    16'b00001111_10010011 : OUT <= 0;  //15 / 147 = 0
    16'b00001111_10010100 : OUT <= 0;  //15 / 148 = 0
    16'b00001111_10010101 : OUT <= 0;  //15 / 149 = 0
    16'b00001111_10010110 : OUT <= 0;  //15 / 150 = 0
    16'b00001111_10010111 : OUT <= 0;  //15 / 151 = 0
    16'b00001111_10011000 : OUT <= 0;  //15 / 152 = 0
    16'b00001111_10011001 : OUT <= 0;  //15 / 153 = 0
    16'b00001111_10011010 : OUT <= 0;  //15 / 154 = 0
    16'b00001111_10011011 : OUT <= 0;  //15 / 155 = 0
    16'b00001111_10011100 : OUT <= 0;  //15 / 156 = 0
    16'b00001111_10011101 : OUT <= 0;  //15 / 157 = 0
    16'b00001111_10011110 : OUT <= 0;  //15 / 158 = 0
    16'b00001111_10011111 : OUT <= 0;  //15 / 159 = 0
    16'b00001111_10100000 : OUT <= 0;  //15 / 160 = 0
    16'b00001111_10100001 : OUT <= 0;  //15 / 161 = 0
    16'b00001111_10100010 : OUT <= 0;  //15 / 162 = 0
    16'b00001111_10100011 : OUT <= 0;  //15 / 163 = 0
    16'b00001111_10100100 : OUT <= 0;  //15 / 164 = 0
    16'b00001111_10100101 : OUT <= 0;  //15 / 165 = 0
    16'b00001111_10100110 : OUT <= 0;  //15 / 166 = 0
    16'b00001111_10100111 : OUT <= 0;  //15 / 167 = 0
    16'b00001111_10101000 : OUT <= 0;  //15 / 168 = 0
    16'b00001111_10101001 : OUT <= 0;  //15 / 169 = 0
    16'b00001111_10101010 : OUT <= 0;  //15 / 170 = 0
    16'b00001111_10101011 : OUT <= 0;  //15 / 171 = 0
    16'b00001111_10101100 : OUT <= 0;  //15 / 172 = 0
    16'b00001111_10101101 : OUT <= 0;  //15 / 173 = 0
    16'b00001111_10101110 : OUT <= 0;  //15 / 174 = 0
    16'b00001111_10101111 : OUT <= 0;  //15 / 175 = 0
    16'b00001111_10110000 : OUT <= 0;  //15 / 176 = 0
    16'b00001111_10110001 : OUT <= 0;  //15 / 177 = 0
    16'b00001111_10110010 : OUT <= 0;  //15 / 178 = 0
    16'b00001111_10110011 : OUT <= 0;  //15 / 179 = 0
    16'b00001111_10110100 : OUT <= 0;  //15 / 180 = 0
    16'b00001111_10110101 : OUT <= 0;  //15 / 181 = 0
    16'b00001111_10110110 : OUT <= 0;  //15 / 182 = 0
    16'b00001111_10110111 : OUT <= 0;  //15 / 183 = 0
    16'b00001111_10111000 : OUT <= 0;  //15 / 184 = 0
    16'b00001111_10111001 : OUT <= 0;  //15 / 185 = 0
    16'b00001111_10111010 : OUT <= 0;  //15 / 186 = 0
    16'b00001111_10111011 : OUT <= 0;  //15 / 187 = 0
    16'b00001111_10111100 : OUT <= 0;  //15 / 188 = 0
    16'b00001111_10111101 : OUT <= 0;  //15 / 189 = 0
    16'b00001111_10111110 : OUT <= 0;  //15 / 190 = 0
    16'b00001111_10111111 : OUT <= 0;  //15 / 191 = 0
    16'b00001111_11000000 : OUT <= 0;  //15 / 192 = 0
    16'b00001111_11000001 : OUT <= 0;  //15 / 193 = 0
    16'b00001111_11000010 : OUT <= 0;  //15 / 194 = 0
    16'b00001111_11000011 : OUT <= 0;  //15 / 195 = 0
    16'b00001111_11000100 : OUT <= 0;  //15 / 196 = 0
    16'b00001111_11000101 : OUT <= 0;  //15 / 197 = 0
    16'b00001111_11000110 : OUT <= 0;  //15 / 198 = 0
    16'b00001111_11000111 : OUT <= 0;  //15 / 199 = 0
    16'b00001111_11001000 : OUT <= 0;  //15 / 200 = 0
    16'b00001111_11001001 : OUT <= 0;  //15 / 201 = 0
    16'b00001111_11001010 : OUT <= 0;  //15 / 202 = 0
    16'b00001111_11001011 : OUT <= 0;  //15 / 203 = 0
    16'b00001111_11001100 : OUT <= 0;  //15 / 204 = 0
    16'b00001111_11001101 : OUT <= 0;  //15 / 205 = 0
    16'b00001111_11001110 : OUT <= 0;  //15 / 206 = 0
    16'b00001111_11001111 : OUT <= 0;  //15 / 207 = 0
    16'b00001111_11010000 : OUT <= 0;  //15 / 208 = 0
    16'b00001111_11010001 : OUT <= 0;  //15 / 209 = 0
    16'b00001111_11010010 : OUT <= 0;  //15 / 210 = 0
    16'b00001111_11010011 : OUT <= 0;  //15 / 211 = 0
    16'b00001111_11010100 : OUT <= 0;  //15 / 212 = 0
    16'b00001111_11010101 : OUT <= 0;  //15 / 213 = 0
    16'b00001111_11010110 : OUT <= 0;  //15 / 214 = 0
    16'b00001111_11010111 : OUT <= 0;  //15 / 215 = 0
    16'b00001111_11011000 : OUT <= 0;  //15 / 216 = 0
    16'b00001111_11011001 : OUT <= 0;  //15 / 217 = 0
    16'b00001111_11011010 : OUT <= 0;  //15 / 218 = 0
    16'b00001111_11011011 : OUT <= 0;  //15 / 219 = 0
    16'b00001111_11011100 : OUT <= 0;  //15 / 220 = 0
    16'b00001111_11011101 : OUT <= 0;  //15 / 221 = 0
    16'b00001111_11011110 : OUT <= 0;  //15 / 222 = 0
    16'b00001111_11011111 : OUT <= 0;  //15 / 223 = 0
    16'b00001111_11100000 : OUT <= 0;  //15 / 224 = 0
    16'b00001111_11100001 : OUT <= 0;  //15 / 225 = 0
    16'b00001111_11100010 : OUT <= 0;  //15 / 226 = 0
    16'b00001111_11100011 : OUT <= 0;  //15 / 227 = 0
    16'b00001111_11100100 : OUT <= 0;  //15 / 228 = 0
    16'b00001111_11100101 : OUT <= 0;  //15 / 229 = 0
    16'b00001111_11100110 : OUT <= 0;  //15 / 230 = 0
    16'b00001111_11100111 : OUT <= 0;  //15 / 231 = 0
    16'b00001111_11101000 : OUT <= 0;  //15 / 232 = 0
    16'b00001111_11101001 : OUT <= 0;  //15 / 233 = 0
    16'b00001111_11101010 : OUT <= 0;  //15 / 234 = 0
    16'b00001111_11101011 : OUT <= 0;  //15 / 235 = 0
    16'b00001111_11101100 : OUT <= 0;  //15 / 236 = 0
    16'b00001111_11101101 : OUT <= 0;  //15 / 237 = 0
    16'b00001111_11101110 : OUT <= 0;  //15 / 238 = 0
    16'b00001111_11101111 : OUT <= 0;  //15 / 239 = 0
    16'b00001111_11110000 : OUT <= 0;  //15 / 240 = 0
    16'b00001111_11110001 : OUT <= 0;  //15 / 241 = 0
    16'b00001111_11110010 : OUT <= 0;  //15 / 242 = 0
    16'b00001111_11110011 : OUT <= 0;  //15 / 243 = 0
    16'b00001111_11110100 : OUT <= 0;  //15 / 244 = 0
    16'b00001111_11110101 : OUT <= 0;  //15 / 245 = 0
    16'b00001111_11110110 : OUT <= 0;  //15 / 246 = 0
    16'b00001111_11110111 : OUT <= 0;  //15 / 247 = 0
    16'b00001111_11111000 : OUT <= 0;  //15 / 248 = 0
    16'b00001111_11111001 : OUT <= 0;  //15 / 249 = 0
    16'b00001111_11111010 : OUT <= 0;  //15 / 250 = 0
    16'b00001111_11111011 : OUT <= 0;  //15 / 251 = 0
    16'b00001111_11111100 : OUT <= 0;  //15 / 252 = 0
    16'b00001111_11111101 : OUT <= 0;  //15 / 253 = 0
    16'b00001111_11111110 : OUT <= 0;  //15 / 254 = 0
    16'b00001111_11111111 : OUT <= 0;  //15 / 255 = 0
    16'b00010000_00000000 : OUT <= 0;  //16 / 0 = 0
    16'b00010000_00000001 : OUT <= 16;  //16 / 1 = 16
    16'b00010000_00000010 : OUT <= 8;  //16 / 2 = 8
    16'b00010000_00000011 : OUT <= 5;  //16 / 3 = 5
    16'b00010000_00000100 : OUT <= 4;  //16 / 4 = 4
    16'b00010000_00000101 : OUT <= 3;  //16 / 5 = 3
    16'b00010000_00000110 : OUT <= 2;  //16 / 6 = 2
    16'b00010000_00000111 : OUT <= 2;  //16 / 7 = 2
    16'b00010000_00001000 : OUT <= 2;  //16 / 8 = 2
    16'b00010000_00001001 : OUT <= 1;  //16 / 9 = 1
    16'b00010000_00001010 : OUT <= 1;  //16 / 10 = 1
    16'b00010000_00001011 : OUT <= 1;  //16 / 11 = 1
    16'b00010000_00001100 : OUT <= 1;  //16 / 12 = 1
    16'b00010000_00001101 : OUT <= 1;  //16 / 13 = 1
    16'b00010000_00001110 : OUT <= 1;  //16 / 14 = 1
    16'b00010000_00001111 : OUT <= 1;  //16 / 15 = 1
    16'b00010000_00010000 : OUT <= 1;  //16 / 16 = 1
    16'b00010000_00010001 : OUT <= 0;  //16 / 17 = 0
    16'b00010000_00010010 : OUT <= 0;  //16 / 18 = 0
    16'b00010000_00010011 : OUT <= 0;  //16 / 19 = 0
    16'b00010000_00010100 : OUT <= 0;  //16 / 20 = 0
    16'b00010000_00010101 : OUT <= 0;  //16 / 21 = 0
    16'b00010000_00010110 : OUT <= 0;  //16 / 22 = 0
    16'b00010000_00010111 : OUT <= 0;  //16 / 23 = 0
    16'b00010000_00011000 : OUT <= 0;  //16 / 24 = 0
    16'b00010000_00011001 : OUT <= 0;  //16 / 25 = 0
    16'b00010000_00011010 : OUT <= 0;  //16 / 26 = 0
    16'b00010000_00011011 : OUT <= 0;  //16 / 27 = 0
    16'b00010000_00011100 : OUT <= 0;  //16 / 28 = 0
    16'b00010000_00011101 : OUT <= 0;  //16 / 29 = 0
    16'b00010000_00011110 : OUT <= 0;  //16 / 30 = 0
    16'b00010000_00011111 : OUT <= 0;  //16 / 31 = 0
    16'b00010000_00100000 : OUT <= 0;  //16 / 32 = 0
    16'b00010000_00100001 : OUT <= 0;  //16 / 33 = 0
    16'b00010000_00100010 : OUT <= 0;  //16 / 34 = 0
    16'b00010000_00100011 : OUT <= 0;  //16 / 35 = 0
    16'b00010000_00100100 : OUT <= 0;  //16 / 36 = 0
    16'b00010000_00100101 : OUT <= 0;  //16 / 37 = 0
    16'b00010000_00100110 : OUT <= 0;  //16 / 38 = 0
    16'b00010000_00100111 : OUT <= 0;  //16 / 39 = 0
    16'b00010000_00101000 : OUT <= 0;  //16 / 40 = 0
    16'b00010000_00101001 : OUT <= 0;  //16 / 41 = 0
    16'b00010000_00101010 : OUT <= 0;  //16 / 42 = 0
    16'b00010000_00101011 : OUT <= 0;  //16 / 43 = 0
    16'b00010000_00101100 : OUT <= 0;  //16 / 44 = 0
    16'b00010000_00101101 : OUT <= 0;  //16 / 45 = 0
    16'b00010000_00101110 : OUT <= 0;  //16 / 46 = 0
    16'b00010000_00101111 : OUT <= 0;  //16 / 47 = 0
    16'b00010000_00110000 : OUT <= 0;  //16 / 48 = 0
    16'b00010000_00110001 : OUT <= 0;  //16 / 49 = 0
    16'b00010000_00110010 : OUT <= 0;  //16 / 50 = 0
    16'b00010000_00110011 : OUT <= 0;  //16 / 51 = 0
    16'b00010000_00110100 : OUT <= 0;  //16 / 52 = 0
    16'b00010000_00110101 : OUT <= 0;  //16 / 53 = 0
    16'b00010000_00110110 : OUT <= 0;  //16 / 54 = 0
    16'b00010000_00110111 : OUT <= 0;  //16 / 55 = 0
    16'b00010000_00111000 : OUT <= 0;  //16 / 56 = 0
    16'b00010000_00111001 : OUT <= 0;  //16 / 57 = 0
    16'b00010000_00111010 : OUT <= 0;  //16 / 58 = 0
    16'b00010000_00111011 : OUT <= 0;  //16 / 59 = 0
    16'b00010000_00111100 : OUT <= 0;  //16 / 60 = 0
    16'b00010000_00111101 : OUT <= 0;  //16 / 61 = 0
    16'b00010000_00111110 : OUT <= 0;  //16 / 62 = 0
    16'b00010000_00111111 : OUT <= 0;  //16 / 63 = 0
    16'b00010000_01000000 : OUT <= 0;  //16 / 64 = 0
    16'b00010000_01000001 : OUT <= 0;  //16 / 65 = 0
    16'b00010000_01000010 : OUT <= 0;  //16 / 66 = 0
    16'b00010000_01000011 : OUT <= 0;  //16 / 67 = 0
    16'b00010000_01000100 : OUT <= 0;  //16 / 68 = 0
    16'b00010000_01000101 : OUT <= 0;  //16 / 69 = 0
    16'b00010000_01000110 : OUT <= 0;  //16 / 70 = 0
    16'b00010000_01000111 : OUT <= 0;  //16 / 71 = 0
    16'b00010000_01001000 : OUT <= 0;  //16 / 72 = 0
    16'b00010000_01001001 : OUT <= 0;  //16 / 73 = 0
    16'b00010000_01001010 : OUT <= 0;  //16 / 74 = 0
    16'b00010000_01001011 : OUT <= 0;  //16 / 75 = 0
    16'b00010000_01001100 : OUT <= 0;  //16 / 76 = 0
    16'b00010000_01001101 : OUT <= 0;  //16 / 77 = 0
    16'b00010000_01001110 : OUT <= 0;  //16 / 78 = 0
    16'b00010000_01001111 : OUT <= 0;  //16 / 79 = 0
    16'b00010000_01010000 : OUT <= 0;  //16 / 80 = 0
    16'b00010000_01010001 : OUT <= 0;  //16 / 81 = 0
    16'b00010000_01010010 : OUT <= 0;  //16 / 82 = 0
    16'b00010000_01010011 : OUT <= 0;  //16 / 83 = 0
    16'b00010000_01010100 : OUT <= 0;  //16 / 84 = 0
    16'b00010000_01010101 : OUT <= 0;  //16 / 85 = 0
    16'b00010000_01010110 : OUT <= 0;  //16 / 86 = 0
    16'b00010000_01010111 : OUT <= 0;  //16 / 87 = 0
    16'b00010000_01011000 : OUT <= 0;  //16 / 88 = 0
    16'b00010000_01011001 : OUT <= 0;  //16 / 89 = 0
    16'b00010000_01011010 : OUT <= 0;  //16 / 90 = 0
    16'b00010000_01011011 : OUT <= 0;  //16 / 91 = 0
    16'b00010000_01011100 : OUT <= 0;  //16 / 92 = 0
    16'b00010000_01011101 : OUT <= 0;  //16 / 93 = 0
    16'b00010000_01011110 : OUT <= 0;  //16 / 94 = 0
    16'b00010000_01011111 : OUT <= 0;  //16 / 95 = 0
    16'b00010000_01100000 : OUT <= 0;  //16 / 96 = 0
    16'b00010000_01100001 : OUT <= 0;  //16 / 97 = 0
    16'b00010000_01100010 : OUT <= 0;  //16 / 98 = 0
    16'b00010000_01100011 : OUT <= 0;  //16 / 99 = 0
    16'b00010000_01100100 : OUT <= 0;  //16 / 100 = 0
    16'b00010000_01100101 : OUT <= 0;  //16 / 101 = 0
    16'b00010000_01100110 : OUT <= 0;  //16 / 102 = 0
    16'b00010000_01100111 : OUT <= 0;  //16 / 103 = 0
    16'b00010000_01101000 : OUT <= 0;  //16 / 104 = 0
    16'b00010000_01101001 : OUT <= 0;  //16 / 105 = 0
    16'b00010000_01101010 : OUT <= 0;  //16 / 106 = 0
    16'b00010000_01101011 : OUT <= 0;  //16 / 107 = 0
    16'b00010000_01101100 : OUT <= 0;  //16 / 108 = 0
    16'b00010000_01101101 : OUT <= 0;  //16 / 109 = 0
    16'b00010000_01101110 : OUT <= 0;  //16 / 110 = 0
    16'b00010000_01101111 : OUT <= 0;  //16 / 111 = 0
    16'b00010000_01110000 : OUT <= 0;  //16 / 112 = 0
    16'b00010000_01110001 : OUT <= 0;  //16 / 113 = 0
    16'b00010000_01110010 : OUT <= 0;  //16 / 114 = 0
    16'b00010000_01110011 : OUT <= 0;  //16 / 115 = 0
    16'b00010000_01110100 : OUT <= 0;  //16 / 116 = 0
    16'b00010000_01110101 : OUT <= 0;  //16 / 117 = 0
    16'b00010000_01110110 : OUT <= 0;  //16 / 118 = 0
    16'b00010000_01110111 : OUT <= 0;  //16 / 119 = 0
    16'b00010000_01111000 : OUT <= 0;  //16 / 120 = 0
    16'b00010000_01111001 : OUT <= 0;  //16 / 121 = 0
    16'b00010000_01111010 : OUT <= 0;  //16 / 122 = 0
    16'b00010000_01111011 : OUT <= 0;  //16 / 123 = 0
    16'b00010000_01111100 : OUT <= 0;  //16 / 124 = 0
    16'b00010000_01111101 : OUT <= 0;  //16 / 125 = 0
    16'b00010000_01111110 : OUT <= 0;  //16 / 126 = 0
    16'b00010000_01111111 : OUT <= 0;  //16 / 127 = 0
    16'b00010000_10000000 : OUT <= 0;  //16 / 128 = 0
    16'b00010000_10000001 : OUT <= 0;  //16 / 129 = 0
    16'b00010000_10000010 : OUT <= 0;  //16 / 130 = 0
    16'b00010000_10000011 : OUT <= 0;  //16 / 131 = 0
    16'b00010000_10000100 : OUT <= 0;  //16 / 132 = 0
    16'b00010000_10000101 : OUT <= 0;  //16 / 133 = 0
    16'b00010000_10000110 : OUT <= 0;  //16 / 134 = 0
    16'b00010000_10000111 : OUT <= 0;  //16 / 135 = 0
    16'b00010000_10001000 : OUT <= 0;  //16 / 136 = 0
    16'b00010000_10001001 : OUT <= 0;  //16 / 137 = 0
    16'b00010000_10001010 : OUT <= 0;  //16 / 138 = 0
    16'b00010000_10001011 : OUT <= 0;  //16 / 139 = 0
    16'b00010000_10001100 : OUT <= 0;  //16 / 140 = 0
    16'b00010000_10001101 : OUT <= 0;  //16 / 141 = 0
    16'b00010000_10001110 : OUT <= 0;  //16 / 142 = 0
    16'b00010000_10001111 : OUT <= 0;  //16 / 143 = 0
    16'b00010000_10010000 : OUT <= 0;  //16 / 144 = 0
    16'b00010000_10010001 : OUT <= 0;  //16 / 145 = 0
    16'b00010000_10010010 : OUT <= 0;  //16 / 146 = 0
    16'b00010000_10010011 : OUT <= 0;  //16 / 147 = 0
    16'b00010000_10010100 : OUT <= 0;  //16 / 148 = 0
    16'b00010000_10010101 : OUT <= 0;  //16 / 149 = 0
    16'b00010000_10010110 : OUT <= 0;  //16 / 150 = 0
    16'b00010000_10010111 : OUT <= 0;  //16 / 151 = 0
    16'b00010000_10011000 : OUT <= 0;  //16 / 152 = 0
    16'b00010000_10011001 : OUT <= 0;  //16 / 153 = 0
    16'b00010000_10011010 : OUT <= 0;  //16 / 154 = 0
    16'b00010000_10011011 : OUT <= 0;  //16 / 155 = 0
    16'b00010000_10011100 : OUT <= 0;  //16 / 156 = 0
    16'b00010000_10011101 : OUT <= 0;  //16 / 157 = 0
    16'b00010000_10011110 : OUT <= 0;  //16 / 158 = 0
    16'b00010000_10011111 : OUT <= 0;  //16 / 159 = 0
    16'b00010000_10100000 : OUT <= 0;  //16 / 160 = 0
    16'b00010000_10100001 : OUT <= 0;  //16 / 161 = 0
    16'b00010000_10100010 : OUT <= 0;  //16 / 162 = 0
    16'b00010000_10100011 : OUT <= 0;  //16 / 163 = 0
    16'b00010000_10100100 : OUT <= 0;  //16 / 164 = 0
    16'b00010000_10100101 : OUT <= 0;  //16 / 165 = 0
    16'b00010000_10100110 : OUT <= 0;  //16 / 166 = 0
    16'b00010000_10100111 : OUT <= 0;  //16 / 167 = 0
    16'b00010000_10101000 : OUT <= 0;  //16 / 168 = 0
    16'b00010000_10101001 : OUT <= 0;  //16 / 169 = 0
    16'b00010000_10101010 : OUT <= 0;  //16 / 170 = 0
    16'b00010000_10101011 : OUT <= 0;  //16 / 171 = 0
    16'b00010000_10101100 : OUT <= 0;  //16 / 172 = 0
    16'b00010000_10101101 : OUT <= 0;  //16 / 173 = 0
    16'b00010000_10101110 : OUT <= 0;  //16 / 174 = 0
    16'b00010000_10101111 : OUT <= 0;  //16 / 175 = 0
    16'b00010000_10110000 : OUT <= 0;  //16 / 176 = 0
    16'b00010000_10110001 : OUT <= 0;  //16 / 177 = 0
    16'b00010000_10110010 : OUT <= 0;  //16 / 178 = 0
    16'b00010000_10110011 : OUT <= 0;  //16 / 179 = 0
    16'b00010000_10110100 : OUT <= 0;  //16 / 180 = 0
    16'b00010000_10110101 : OUT <= 0;  //16 / 181 = 0
    16'b00010000_10110110 : OUT <= 0;  //16 / 182 = 0
    16'b00010000_10110111 : OUT <= 0;  //16 / 183 = 0
    16'b00010000_10111000 : OUT <= 0;  //16 / 184 = 0
    16'b00010000_10111001 : OUT <= 0;  //16 / 185 = 0
    16'b00010000_10111010 : OUT <= 0;  //16 / 186 = 0
    16'b00010000_10111011 : OUT <= 0;  //16 / 187 = 0
    16'b00010000_10111100 : OUT <= 0;  //16 / 188 = 0
    16'b00010000_10111101 : OUT <= 0;  //16 / 189 = 0
    16'b00010000_10111110 : OUT <= 0;  //16 / 190 = 0
    16'b00010000_10111111 : OUT <= 0;  //16 / 191 = 0
    16'b00010000_11000000 : OUT <= 0;  //16 / 192 = 0
    16'b00010000_11000001 : OUT <= 0;  //16 / 193 = 0
    16'b00010000_11000010 : OUT <= 0;  //16 / 194 = 0
    16'b00010000_11000011 : OUT <= 0;  //16 / 195 = 0
    16'b00010000_11000100 : OUT <= 0;  //16 / 196 = 0
    16'b00010000_11000101 : OUT <= 0;  //16 / 197 = 0
    16'b00010000_11000110 : OUT <= 0;  //16 / 198 = 0
    16'b00010000_11000111 : OUT <= 0;  //16 / 199 = 0
    16'b00010000_11001000 : OUT <= 0;  //16 / 200 = 0
    16'b00010000_11001001 : OUT <= 0;  //16 / 201 = 0
    16'b00010000_11001010 : OUT <= 0;  //16 / 202 = 0
    16'b00010000_11001011 : OUT <= 0;  //16 / 203 = 0
    16'b00010000_11001100 : OUT <= 0;  //16 / 204 = 0
    16'b00010000_11001101 : OUT <= 0;  //16 / 205 = 0
    16'b00010000_11001110 : OUT <= 0;  //16 / 206 = 0
    16'b00010000_11001111 : OUT <= 0;  //16 / 207 = 0
    16'b00010000_11010000 : OUT <= 0;  //16 / 208 = 0
    16'b00010000_11010001 : OUT <= 0;  //16 / 209 = 0
    16'b00010000_11010010 : OUT <= 0;  //16 / 210 = 0
    16'b00010000_11010011 : OUT <= 0;  //16 / 211 = 0
    16'b00010000_11010100 : OUT <= 0;  //16 / 212 = 0
    16'b00010000_11010101 : OUT <= 0;  //16 / 213 = 0
    16'b00010000_11010110 : OUT <= 0;  //16 / 214 = 0
    16'b00010000_11010111 : OUT <= 0;  //16 / 215 = 0
    16'b00010000_11011000 : OUT <= 0;  //16 / 216 = 0
    16'b00010000_11011001 : OUT <= 0;  //16 / 217 = 0
    16'b00010000_11011010 : OUT <= 0;  //16 / 218 = 0
    16'b00010000_11011011 : OUT <= 0;  //16 / 219 = 0
    16'b00010000_11011100 : OUT <= 0;  //16 / 220 = 0
    16'b00010000_11011101 : OUT <= 0;  //16 / 221 = 0
    16'b00010000_11011110 : OUT <= 0;  //16 / 222 = 0
    16'b00010000_11011111 : OUT <= 0;  //16 / 223 = 0
    16'b00010000_11100000 : OUT <= 0;  //16 / 224 = 0
    16'b00010000_11100001 : OUT <= 0;  //16 / 225 = 0
    16'b00010000_11100010 : OUT <= 0;  //16 / 226 = 0
    16'b00010000_11100011 : OUT <= 0;  //16 / 227 = 0
    16'b00010000_11100100 : OUT <= 0;  //16 / 228 = 0
    16'b00010000_11100101 : OUT <= 0;  //16 / 229 = 0
    16'b00010000_11100110 : OUT <= 0;  //16 / 230 = 0
    16'b00010000_11100111 : OUT <= 0;  //16 / 231 = 0
    16'b00010000_11101000 : OUT <= 0;  //16 / 232 = 0
    16'b00010000_11101001 : OUT <= 0;  //16 / 233 = 0
    16'b00010000_11101010 : OUT <= 0;  //16 / 234 = 0
    16'b00010000_11101011 : OUT <= 0;  //16 / 235 = 0
    16'b00010000_11101100 : OUT <= 0;  //16 / 236 = 0
    16'b00010000_11101101 : OUT <= 0;  //16 / 237 = 0
    16'b00010000_11101110 : OUT <= 0;  //16 / 238 = 0
    16'b00010000_11101111 : OUT <= 0;  //16 / 239 = 0
    16'b00010000_11110000 : OUT <= 0;  //16 / 240 = 0
    16'b00010000_11110001 : OUT <= 0;  //16 / 241 = 0
    16'b00010000_11110010 : OUT <= 0;  //16 / 242 = 0
    16'b00010000_11110011 : OUT <= 0;  //16 / 243 = 0
    16'b00010000_11110100 : OUT <= 0;  //16 / 244 = 0
    16'b00010000_11110101 : OUT <= 0;  //16 / 245 = 0
    16'b00010000_11110110 : OUT <= 0;  //16 / 246 = 0
    16'b00010000_11110111 : OUT <= 0;  //16 / 247 = 0
    16'b00010000_11111000 : OUT <= 0;  //16 / 248 = 0
    16'b00010000_11111001 : OUT <= 0;  //16 / 249 = 0
    16'b00010000_11111010 : OUT <= 0;  //16 / 250 = 0
    16'b00010000_11111011 : OUT <= 0;  //16 / 251 = 0
    16'b00010000_11111100 : OUT <= 0;  //16 / 252 = 0
    16'b00010000_11111101 : OUT <= 0;  //16 / 253 = 0
    16'b00010000_11111110 : OUT <= 0;  //16 / 254 = 0
    16'b00010000_11111111 : OUT <= 0;  //16 / 255 = 0
    16'b00010001_00000000 : OUT <= 0;  //17 / 0 = 0
    16'b00010001_00000001 : OUT <= 17;  //17 / 1 = 17
    16'b00010001_00000010 : OUT <= 8;  //17 / 2 = 8
    16'b00010001_00000011 : OUT <= 5;  //17 / 3 = 5
    16'b00010001_00000100 : OUT <= 4;  //17 / 4 = 4
    16'b00010001_00000101 : OUT <= 3;  //17 / 5 = 3
    16'b00010001_00000110 : OUT <= 2;  //17 / 6 = 2
    16'b00010001_00000111 : OUT <= 2;  //17 / 7 = 2
    16'b00010001_00001000 : OUT <= 2;  //17 / 8 = 2
    16'b00010001_00001001 : OUT <= 1;  //17 / 9 = 1
    16'b00010001_00001010 : OUT <= 1;  //17 / 10 = 1
    16'b00010001_00001011 : OUT <= 1;  //17 / 11 = 1
    16'b00010001_00001100 : OUT <= 1;  //17 / 12 = 1
    16'b00010001_00001101 : OUT <= 1;  //17 / 13 = 1
    16'b00010001_00001110 : OUT <= 1;  //17 / 14 = 1
    16'b00010001_00001111 : OUT <= 1;  //17 / 15 = 1
    16'b00010001_00010000 : OUT <= 1;  //17 / 16 = 1
    16'b00010001_00010001 : OUT <= 1;  //17 / 17 = 1
    16'b00010001_00010010 : OUT <= 0;  //17 / 18 = 0
    16'b00010001_00010011 : OUT <= 0;  //17 / 19 = 0
    16'b00010001_00010100 : OUT <= 0;  //17 / 20 = 0
    16'b00010001_00010101 : OUT <= 0;  //17 / 21 = 0
    16'b00010001_00010110 : OUT <= 0;  //17 / 22 = 0
    16'b00010001_00010111 : OUT <= 0;  //17 / 23 = 0
    16'b00010001_00011000 : OUT <= 0;  //17 / 24 = 0
    16'b00010001_00011001 : OUT <= 0;  //17 / 25 = 0
    16'b00010001_00011010 : OUT <= 0;  //17 / 26 = 0
    16'b00010001_00011011 : OUT <= 0;  //17 / 27 = 0
    16'b00010001_00011100 : OUT <= 0;  //17 / 28 = 0
    16'b00010001_00011101 : OUT <= 0;  //17 / 29 = 0
    16'b00010001_00011110 : OUT <= 0;  //17 / 30 = 0
    16'b00010001_00011111 : OUT <= 0;  //17 / 31 = 0
    16'b00010001_00100000 : OUT <= 0;  //17 / 32 = 0
    16'b00010001_00100001 : OUT <= 0;  //17 / 33 = 0
    16'b00010001_00100010 : OUT <= 0;  //17 / 34 = 0
    16'b00010001_00100011 : OUT <= 0;  //17 / 35 = 0
    16'b00010001_00100100 : OUT <= 0;  //17 / 36 = 0
    16'b00010001_00100101 : OUT <= 0;  //17 / 37 = 0
    16'b00010001_00100110 : OUT <= 0;  //17 / 38 = 0
    16'b00010001_00100111 : OUT <= 0;  //17 / 39 = 0
    16'b00010001_00101000 : OUT <= 0;  //17 / 40 = 0
    16'b00010001_00101001 : OUT <= 0;  //17 / 41 = 0
    16'b00010001_00101010 : OUT <= 0;  //17 / 42 = 0
    16'b00010001_00101011 : OUT <= 0;  //17 / 43 = 0
    16'b00010001_00101100 : OUT <= 0;  //17 / 44 = 0
    16'b00010001_00101101 : OUT <= 0;  //17 / 45 = 0
    16'b00010001_00101110 : OUT <= 0;  //17 / 46 = 0
    16'b00010001_00101111 : OUT <= 0;  //17 / 47 = 0
    16'b00010001_00110000 : OUT <= 0;  //17 / 48 = 0
    16'b00010001_00110001 : OUT <= 0;  //17 / 49 = 0
    16'b00010001_00110010 : OUT <= 0;  //17 / 50 = 0
    16'b00010001_00110011 : OUT <= 0;  //17 / 51 = 0
    16'b00010001_00110100 : OUT <= 0;  //17 / 52 = 0
    16'b00010001_00110101 : OUT <= 0;  //17 / 53 = 0
    16'b00010001_00110110 : OUT <= 0;  //17 / 54 = 0
    16'b00010001_00110111 : OUT <= 0;  //17 / 55 = 0
    16'b00010001_00111000 : OUT <= 0;  //17 / 56 = 0
    16'b00010001_00111001 : OUT <= 0;  //17 / 57 = 0
    16'b00010001_00111010 : OUT <= 0;  //17 / 58 = 0
    16'b00010001_00111011 : OUT <= 0;  //17 / 59 = 0
    16'b00010001_00111100 : OUT <= 0;  //17 / 60 = 0
    16'b00010001_00111101 : OUT <= 0;  //17 / 61 = 0
    16'b00010001_00111110 : OUT <= 0;  //17 / 62 = 0
    16'b00010001_00111111 : OUT <= 0;  //17 / 63 = 0
    16'b00010001_01000000 : OUT <= 0;  //17 / 64 = 0
    16'b00010001_01000001 : OUT <= 0;  //17 / 65 = 0
    16'b00010001_01000010 : OUT <= 0;  //17 / 66 = 0
    16'b00010001_01000011 : OUT <= 0;  //17 / 67 = 0
    16'b00010001_01000100 : OUT <= 0;  //17 / 68 = 0
    16'b00010001_01000101 : OUT <= 0;  //17 / 69 = 0
    16'b00010001_01000110 : OUT <= 0;  //17 / 70 = 0
    16'b00010001_01000111 : OUT <= 0;  //17 / 71 = 0
    16'b00010001_01001000 : OUT <= 0;  //17 / 72 = 0
    16'b00010001_01001001 : OUT <= 0;  //17 / 73 = 0
    16'b00010001_01001010 : OUT <= 0;  //17 / 74 = 0
    16'b00010001_01001011 : OUT <= 0;  //17 / 75 = 0
    16'b00010001_01001100 : OUT <= 0;  //17 / 76 = 0
    16'b00010001_01001101 : OUT <= 0;  //17 / 77 = 0
    16'b00010001_01001110 : OUT <= 0;  //17 / 78 = 0
    16'b00010001_01001111 : OUT <= 0;  //17 / 79 = 0
    16'b00010001_01010000 : OUT <= 0;  //17 / 80 = 0
    16'b00010001_01010001 : OUT <= 0;  //17 / 81 = 0
    16'b00010001_01010010 : OUT <= 0;  //17 / 82 = 0
    16'b00010001_01010011 : OUT <= 0;  //17 / 83 = 0
    16'b00010001_01010100 : OUT <= 0;  //17 / 84 = 0
    16'b00010001_01010101 : OUT <= 0;  //17 / 85 = 0
    16'b00010001_01010110 : OUT <= 0;  //17 / 86 = 0
    16'b00010001_01010111 : OUT <= 0;  //17 / 87 = 0
    16'b00010001_01011000 : OUT <= 0;  //17 / 88 = 0
    16'b00010001_01011001 : OUT <= 0;  //17 / 89 = 0
    16'b00010001_01011010 : OUT <= 0;  //17 / 90 = 0
    16'b00010001_01011011 : OUT <= 0;  //17 / 91 = 0
    16'b00010001_01011100 : OUT <= 0;  //17 / 92 = 0
    16'b00010001_01011101 : OUT <= 0;  //17 / 93 = 0
    16'b00010001_01011110 : OUT <= 0;  //17 / 94 = 0
    16'b00010001_01011111 : OUT <= 0;  //17 / 95 = 0
    16'b00010001_01100000 : OUT <= 0;  //17 / 96 = 0
    16'b00010001_01100001 : OUT <= 0;  //17 / 97 = 0
    16'b00010001_01100010 : OUT <= 0;  //17 / 98 = 0
    16'b00010001_01100011 : OUT <= 0;  //17 / 99 = 0
    16'b00010001_01100100 : OUT <= 0;  //17 / 100 = 0
    16'b00010001_01100101 : OUT <= 0;  //17 / 101 = 0
    16'b00010001_01100110 : OUT <= 0;  //17 / 102 = 0
    16'b00010001_01100111 : OUT <= 0;  //17 / 103 = 0
    16'b00010001_01101000 : OUT <= 0;  //17 / 104 = 0
    16'b00010001_01101001 : OUT <= 0;  //17 / 105 = 0
    16'b00010001_01101010 : OUT <= 0;  //17 / 106 = 0
    16'b00010001_01101011 : OUT <= 0;  //17 / 107 = 0
    16'b00010001_01101100 : OUT <= 0;  //17 / 108 = 0
    16'b00010001_01101101 : OUT <= 0;  //17 / 109 = 0
    16'b00010001_01101110 : OUT <= 0;  //17 / 110 = 0
    16'b00010001_01101111 : OUT <= 0;  //17 / 111 = 0
    16'b00010001_01110000 : OUT <= 0;  //17 / 112 = 0
    16'b00010001_01110001 : OUT <= 0;  //17 / 113 = 0
    16'b00010001_01110010 : OUT <= 0;  //17 / 114 = 0
    16'b00010001_01110011 : OUT <= 0;  //17 / 115 = 0
    16'b00010001_01110100 : OUT <= 0;  //17 / 116 = 0
    16'b00010001_01110101 : OUT <= 0;  //17 / 117 = 0
    16'b00010001_01110110 : OUT <= 0;  //17 / 118 = 0
    16'b00010001_01110111 : OUT <= 0;  //17 / 119 = 0
    16'b00010001_01111000 : OUT <= 0;  //17 / 120 = 0
    16'b00010001_01111001 : OUT <= 0;  //17 / 121 = 0
    16'b00010001_01111010 : OUT <= 0;  //17 / 122 = 0
    16'b00010001_01111011 : OUT <= 0;  //17 / 123 = 0
    16'b00010001_01111100 : OUT <= 0;  //17 / 124 = 0
    16'b00010001_01111101 : OUT <= 0;  //17 / 125 = 0
    16'b00010001_01111110 : OUT <= 0;  //17 / 126 = 0
    16'b00010001_01111111 : OUT <= 0;  //17 / 127 = 0
    16'b00010001_10000000 : OUT <= 0;  //17 / 128 = 0
    16'b00010001_10000001 : OUT <= 0;  //17 / 129 = 0
    16'b00010001_10000010 : OUT <= 0;  //17 / 130 = 0
    16'b00010001_10000011 : OUT <= 0;  //17 / 131 = 0
    16'b00010001_10000100 : OUT <= 0;  //17 / 132 = 0
    16'b00010001_10000101 : OUT <= 0;  //17 / 133 = 0
    16'b00010001_10000110 : OUT <= 0;  //17 / 134 = 0
    16'b00010001_10000111 : OUT <= 0;  //17 / 135 = 0
    16'b00010001_10001000 : OUT <= 0;  //17 / 136 = 0
    16'b00010001_10001001 : OUT <= 0;  //17 / 137 = 0
    16'b00010001_10001010 : OUT <= 0;  //17 / 138 = 0
    16'b00010001_10001011 : OUT <= 0;  //17 / 139 = 0
    16'b00010001_10001100 : OUT <= 0;  //17 / 140 = 0
    16'b00010001_10001101 : OUT <= 0;  //17 / 141 = 0
    16'b00010001_10001110 : OUT <= 0;  //17 / 142 = 0
    16'b00010001_10001111 : OUT <= 0;  //17 / 143 = 0
    16'b00010001_10010000 : OUT <= 0;  //17 / 144 = 0
    16'b00010001_10010001 : OUT <= 0;  //17 / 145 = 0
    16'b00010001_10010010 : OUT <= 0;  //17 / 146 = 0
    16'b00010001_10010011 : OUT <= 0;  //17 / 147 = 0
    16'b00010001_10010100 : OUT <= 0;  //17 / 148 = 0
    16'b00010001_10010101 : OUT <= 0;  //17 / 149 = 0
    16'b00010001_10010110 : OUT <= 0;  //17 / 150 = 0
    16'b00010001_10010111 : OUT <= 0;  //17 / 151 = 0
    16'b00010001_10011000 : OUT <= 0;  //17 / 152 = 0
    16'b00010001_10011001 : OUT <= 0;  //17 / 153 = 0
    16'b00010001_10011010 : OUT <= 0;  //17 / 154 = 0
    16'b00010001_10011011 : OUT <= 0;  //17 / 155 = 0
    16'b00010001_10011100 : OUT <= 0;  //17 / 156 = 0
    16'b00010001_10011101 : OUT <= 0;  //17 / 157 = 0
    16'b00010001_10011110 : OUT <= 0;  //17 / 158 = 0
    16'b00010001_10011111 : OUT <= 0;  //17 / 159 = 0
    16'b00010001_10100000 : OUT <= 0;  //17 / 160 = 0
    16'b00010001_10100001 : OUT <= 0;  //17 / 161 = 0
    16'b00010001_10100010 : OUT <= 0;  //17 / 162 = 0
    16'b00010001_10100011 : OUT <= 0;  //17 / 163 = 0
    16'b00010001_10100100 : OUT <= 0;  //17 / 164 = 0
    16'b00010001_10100101 : OUT <= 0;  //17 / 165 = 0
    16'b00010001_10100110 : OUT <= 0;  //17 / 166 = 0
    16'b00010001_10100111 : OUT <= 0;  //17 / 167 = 0
    16'b00010001_10101000 : OUT <= 0;  //17 / 168 = 0
    16'b00010001_10101001 : OUT <= 0;  //17 / 169 = 0
    16'b00010001_10101010 : OUT <= 0;  //17 / 170 = 0
    16'b00010001_10101011 : OUT <= 0;  //17 / 171 = 0
    16'b00010001_10101100 : OUT <= 0;  //17 / 172 = 0
    16'b00010001_10101101 : OUT <= 0;  //17 / 173 = 0
    16'b00010001_10101110 : OUT <= 0;  //17 / 174 = 0
    16'b00010001_10101111 : OUT <= 0;  //17 / 175 = 0
    16'b00010001_10110000 : OUT <= 0;  //17 / 176 = 0
    16'b00010001_10110001 : OUT <= 0;  //17 / 177 = 0
    16'b00010001_10110010 : OUT <= 0;  //17 / 178 = 0
    16'b00010001_10110011 : OUT <= 0;  //17 / 179 = 0
    16'b00010001_10110100 : OUT <= 0;  //17 / 180 = 0
    16'b00010001_10110101 : OUT <= 0;  //17 / 181 = 0
    16'b00010001_10110110 : OUT <= 0;  //17 / 182 = 0
    16'b00010001_10110111 : OUT <= 0;  //17 / 183 = 0
    16'b00010001_10111000 : OUT <= 0;  //17 / 184 = 0
    16'b00010001_10111001 : OUT <= 0;  //17 / 185 = 0
    16'b00010001_10111010 : OUT <= 0;  //17 / 186 = 0
    16'b00010001_10111011 : OUT <= 0;  //17 / 187 = 0
    16'b00010001_10111100 : OUT <= 0;  //17 / 188 = 0
    16'b00010001_10111101 : OUT <= 0;  //17 / 189 = 0
    16'b00010001_10111110 : OUT <= 0;  //17 / 190 = 0
    16'b00010001_10111111 : OUT <= 0;  //17 / 191 = 0
    16'b00010001_11000000 : OUT <= 0;  //17 / 192 = 0
    16'b00010001_11000001 : OUT <= 0;  //17 / 193 = 0
    16'b00010001_11000010 : OUT <= 0;  //17 / 194 = 0
    16'b00010001_11000011 : OUT <= 0;  //17 / 195 = 0
    16'b00010001_11000100 : OUT <= 0;  //17 / 196 = 0
    16'b00010001_11000101 : OUT <= 0;  //17 / 197 = 0
    16'b00010001_11000110 : OUT <= 0;  //17 / 198 = 0
    16'b00010001_11000111 : OUT <= 0;  //17 / 199 = 0
    16'b00010001_11001000 : OUT <= 0;  //17 / 200 = 0
    16'b00010001_11001001 : OUT <= 0;  //17 / 201 = 0
    16'b00010001_11001010 : OUT <= 0;  //17 / 202 = 0
    16'b00010001_11001011 : OUT <= 0;  //17 / 203 = 0
    16'b00010001_11001100 : OUT <= 0;  //17 / 204 = 0
    16'b00010001_11001101 : OUT <= 0;  //17 / 205 = 0
    16'b00010001_11001110 : OUT <= 0;  //17 / 206 = 0
    16'b00010001_11001111 : OUT <= 0;  //17 / 207 = 0
    16'b00010001_11010000 : OUT <= 0;  //17 / 208 = 0
    16'b00010001_11010001 : OUT <= 0;  //17 / 209 = 0
    16'b00010001_11010010 : OUT <= 0;  //17 / 210 = 0
    16'b00010001_11010011 : OUT <= 0;  //17 / 211 = 0
    16'b00010001_11010100 : OUT <= 0;  //17 / 212 = 0
    16'b00010001_11010101 : OUT <= 0;  //17 / 213 = 0
    16'b00010001_11010110 : OUT <= 0;  //17 / 214 = 0
    16'b00010001_11010111 : OUT <= 0;  //17 / 215 = 0
    16'b00010001_11011000 : OUT <= 0;  //17 / 216 = 0
    16'b00010001_11011001 : OUT <= 0;  //17 / 217 = 0
    16'b00010001_11011010 : OUT <= 0;  //17 / 218 = 0
    16'b00010001_11011011 : OUT <= 0;  //17 / 219 = 0
    16'b00010001_11011100 : OUT <= 0;  //17 / 220 = 0
    16'b00010001_11011101 : OUT <= 0;  //17 / 221 = 0
    16'b00010001_11011110 : OUT <= 0;  //17 / 222 = 0
    16'b00010001_11011111 : OUT <= 0;  //17 / 223 = 0
    16'b00010001_11100000 : OUT <= 0;  //17 / 224 = 0
    16'b00010001_11100001 : OUT <= 0;  //17 / 225 = 0
    16'b00010001_11100010 : OUT <= 0;  //17 / 226 = 0
    16'b00010001_11100011 : OUT <= 0;  //17 / 227 = 0
    16'b00010001_11100100 : OUT <= 0;  //17 / 228 = 0
    16'b00010001_11100101 : OUT <= 0;  //17 / 229 = 0
    16'b00010001_11100110 : OUT <= 0;  //17 / 230 = 0
    16'b00010001_11100111 : OUT <= 0;  //17 / 231 = 0
    16'b00010001_11101000 : OUT <= 0;  //17 / 232 = 0
    16'b00010001_11101001 : OUT <= 0;  //17 / 233 = 0
    16'b00010001_11101010 : OUT <= 0;  //17 / 234 = 0
    16'b00010001_11101011 : OUT <= 0;  //17 / 235 = 0
    16'b00010001_11101100 : OUT <= 0;  //17 / 236 = 0
    16'b00010001_11101101 : OUT <= 0;  //17 / 237 = 0
    16'b00010001_11101110 : OUT <= 0;  //17 / 238 = 0
    16'b00010001_11101111 : OUT <= 0;  //17 / 239 = 0
    16'b00010001_11110000 : OUT <= 0;  //17 / 240 = 0
    16'b00010001_11110001 : OUT <= 0;  //17 / 241 = 0
    16'b00010001_11110010 : OUT <= 0;  //17 / 242 = 0
    16'b00010001_11110011 : OUT <= 0;  //17 / 243 = 0
    16'b00010001_11110100 : OUT <= 0;  //17 / 244 = 0
    16'b00010001_11110101 : OUT <= 0;  //17 / 245 = 0
    16'b00010001_11110110 : OUT <= 0;  //17 / 246 = 0
    16'b00010001_11110111 : OUT <= 0;  //17 / 247 = 0
    16'b00010001_11111000 : OUT <= 0;  //17 / 248 = 0
    16'b00010001_11111001 : OUT <= 0;  //17 / 249 = 0
    16'b00010001_11111010 : OUT <= 0;  //17 / 250 = 0
    16'b00010001_11111011 : OUT <= 0;  //17 / 251 = 0
    16'b00010001_11111100 : OUT <= 0;  //17 / 252 = 0
    16'b00010001_11111101 : OUT <= 0;  //17 / 253 = 0
    16'b00010001_11111110 : OUT <= 0;  //17 / 254 = 0
    16'b00010001_11111111 : OUT <= 0;  //17 / 255 = 0
    16'b00010010_00000000 : OUT <= 0;  //18 / 0 = 0
    16'b00010010_00000001 : OUT <= 18;  //18 / 1 = 18
    16'b00010010_00000010 : OUT <= 9;  //18 / 2 = 9
    16'b00010010_00000011 : OUT <= 6;  //18 / 3 = 6
    16'b00010010_00000100 : OUT <= 4;  //18 / 4 = 4
    16'b00010010_00000101 : OUT <= 3;  //18 / 5 = 3
    16'b00010010_00000110 : OUT <= 3;  //18 / 6 = 3
    16'b00010010_00000111 : OUT <= 2;  //18 / 7 = 2
    16'b00010010_00001000 : OUT <= 2;  //18 / 8 = 2
    16'b00010010_00001001 : OUT <= 2;  //18 / 9 = 2
    16'b00010010_00001010 : OUT <= 1;  //18 / 10 = 1
    16'b00010010_00001011 : OUT <= 1;  //18 / 11 = 1
    16'b00010010_00001100 : OUT <= 1;  //18 / 12 = 1
    16'b00010010_00001101 : OUT <= 1;  //18 / 13 = 1
    16'b00010010_00001110 : OUT <= 1;  //18 / 14 = 1
    16'b00010010_00001111 : OUT <= 1;  //18 / 15 = 1
    16'b00010010_00010000 : OUT <= 1;  //18 / 16 = 1
    16'b00010010_00010001 : OUT <= 1;  //18 / 17 = 1
    16'b00010010_00010010 : OUT <= 1;  //18 / 18 = 1
    16'b00010010_00010011 : OUT <= 0;  //18 / 19 = 0
    16'b00010010_00010100 : OUT <= 0;  //18 / 20 = 0
    16'b00010010_00010101 : OUT <= 0;  //18 / 21 = 0
    16'b00010010_00010110 : OUT <= 0;  //18 / 22 = 0
    16'b00010010_00010111 : OUT <= 0;  //18 / 23 = 0
    16'b00010010_00011000 : OUT <= 0;  //18 / 24 = 0
    16'b00010010_00011001 : OUT <= 0;  //18 / 25 = 0
    16'b00010010_00011010 : OUT <= 0;  //18 / 26 = 0
    16'b00010010_00011011 : OUT <= 0;  //18 / 27 = 0
    16'b00010010_00011100 : OUT <= 0;  //18 / 28 = 0
    16'b00010010_00011101 : OUT <= 0;  //18 / 29 = 0
    16'b00010010_00011110 : OUT <= 0;  //18 / 30 = 0
    16'b00010010_00011111 : OUT <= 0;  //18 / 31 = 0
    16'b00010010_00100000 : OUT <= 0;  //18 / 32 = 0
    16'b00010010_00100001 : OUT <= 0;  //18 / 33 = 0
    16'b00010010_00100010 : OUT <= 0;  //18 / 34 = 0
    16'b00010010_00100011 : OUT <= 0;  //18 / 35 = 0
    16'b00010010_00100100 : OUT <= 0;  //18 / 36 = 0
    16'b00010010_00100101 : OUT <= 0;  //18 / 37 = 0
    16'b00010010_00100110 : OUT <= 0;  //18 / 38 = 0
    16'b00010010_00100111 : OUT <= 0;  //18 / 39 = 0
    16'b00010010_00101000 : OUT <= 0;  //18 / 40 = 0
    16'b00010010_00101001 : OUT <= 0;  //18 / 41 = 0
    16'b00010010_00101010 : OUT <= 0;  //18 / 42 = 0
    16'b00010010_00101011 : OUT <= 0;  //18 / 43 = 0
    16'b00010010_00101100 : OUT <= 0;  //18 / 44 = 0
    16'b00010010_00101101 : OUT <= 0;  //18 / 45 = 0
    16'b00010010_00101110 : OUT <= 0;  //18 / 46 = 0
    16'b00010010_00101111 : OUT <= 0;  //18 / 47 = 0
    16'b00010010_00110000 : OUT <= 0;  //18 / 48 = 0
    16'b00010010_00110001 : OUT <= 0;  //18 / 49 = 0
    16'b00010010_00110010 : OUT <= 0;  //18 / 50 = 0
    16'b00010010_00110011 : OUT <= 0;  //18 / 51 = 0
    16'b00010010_00110100 : OUT <= 0;  //18 / 52 = 0
    16'b00010010_00110101 : OUT <= 0;  //18 / 53 = 0
    16'b00010010_00110110 : OUT <= 0;  //18 / 54 = 0
    16'b00010010_00110111 : OUT <= 0;  //18 / 55 = 0
    16'b00010010_00111000 : OUT <= 0;  //18 / 56 = 0
    16'b00010010_00111001 : OUT <= 0;  //18 / 57 = 0
    16'b00010010_00111010 : OUT <= 0;  //18 / 58 = 0
    16'b00010010_00111011 : OUT <= 0;  //18 / 59 = 0
    16'b00010010_00111100 : OUT <= 0;  //18 / 60 = 0
    16'b00010010_00111101 : OUT <= 0;  //18 / 61 = 0
    16'b00010010_00111110 : OUT <= 0;  //18 / 62 = 0
    16'b00010010_00111111 : OUT <= 0;  //18 / 63 = 0
    16'b00010010_01000000 : OUT <= 0;  //18 / 64 = 0
    16'b00010010_01000001 : OUT <= 0;  //18 / 65 = 0
    16'b00010010_01000010 : OUT <= 0;  //18 / 66 = 0
    16'b00010010_01000011 : OUT <= 0;  //18 / 67 = 0
    16'b00010010_01000100 : OUT <= 0;  //18 / 68 = 0
    16'b00010010_01000101 : OUT <= 0;  //18 / 69 = 0
    16'b00010010_01000110 : OUT <= 0;  //18 / 70 = 0
    16'b00010010_01000111 : OUT <= 0;  //18 / 71 = 0
    16'b00010010_01001000 : OUT <= 0;  //18 / 72 = 0
    16'b00010010_01001001 : OUT <= 0;  //18 / 73 = 0
    16'b00010010_01001010 : OUT <= 0;  //18 / 74 = 0
    16'b00010010_01001011 : OUT <= 0;  //18 / 75 = 0
    16'b00010010_01001100 : OUT <= 0;  //18 / 76 = 0
    16'b00010010_01001101 : OUT <= 0;  //18 / 77 = 0
    16'b00010010_01001110 : OUT <= 0;  //18 / 78 = 0
    16'b00010010_01001111 : OUT <= 0;  //18 / 79 = 0
    16'b00010010_01010000 : OUT <= 0;  //18 / 80 = 0
    16'b00010010_01010001 : OUT <= 0;  //18 / 81 = 0
    16'b00010010_01010010 : OUT <= 0;  //18 / 82 = 0
    16'b00010010_01010011 : OUT <= 0;  //18 / 83 = 0
    16'b00010010_01010100 : OUT <= 0;  //18 / 84 = 0
    16'b00010010_01010101 : OUT <= 0;  //18 / 85 = 0
    16'b00010010_01010110 : OUT <= 0;  //18 / 86 = 0
    16'b00010010_01010111 : OUT <= 0;  //18 / 87 = 0
    16'b00010010_01011000 : OUT <= 0;  //18 / 88 = 0
    16'b00010010_01011001 : OUT <= 0;  //18 / 89 = 0
    16'b00010010_01011010 : OUT <= 0;  //18 / 90 = 0
    16'b00010010_01011011 : OUT <= 0;  //18 / 91 = 0
    16'b00010010_01011100 : OUT <= 0;  //18 / 92 = 0
    16'b00010010_01011101 : OUT <= 0;  //18 / 93 = 0
    16'b00010010_01011110 : OUT <= 0;  //18 / 94 = 0
    16'b00010010_01011111 : OUT <= 0;  //18 / 95 = 0
    16'b00010010_01100000 : OUT <= 0;  //18 / 96 = 0
    16'b00010010_01100001 : OUT <= 0;  //18 / 97 = 0
    16'b00010010_01100010 : OUT <= 0;  //18 / 98 = 0
    16'b00010010_01100011 : OUT <= 0;  //18 / 99 = 0
    16'b00010010_01100100 : OUT <= 0;  //18 / 100 = 0
    16'b00010010_01100101 : OUT <= 0;  //18 / 101 = 0
    16'b00010010_01100110 : OUT <= 0;  //18 / 102 = 0
    16'b00010010_01100111 : OUT <= 0;  //18 / 103 = 0
    16'b00010010_01101000 : OUT <= 0;  //18 / 104 = 0
    16'b00010010_01101001 : OUT <= 0;  //18 / 105 = 0
    16'b00010010_01101010 : OUT <= 0;  //18 / 106 = 0
    16'b00010010_01101011 : OUT <= 0;  //18 / 107 = 0
    16'b00010010_01101100 : OUT <= 0;  //18 / 108 = 0
    16'b00010010_01101101 : OUT <= 0;  //18 / 109 = 0
    16'b00010010_01101110 : OUT <= 0;  //18 / 110 = 0
    16'b00010010_01101111 : OUT <= 0;  //18 / 111 = 0
    16'b00010010_01110000 : OUT <= 0;  //18 / 112 = 0
    16'b00010010_01110001 : OUT <= 0;  //18 / 113 = 0
    16'b00010010_01110010 : OUT <= 0;  //18 / 114 = 0
    16'b00010010_01110011 : OUT <= 0;  //18 / 115 = 0
    16'b00010010_01110100 : OUT <= 0;  //18 / 116 = 0
    16'b00010010_01110101 : OUT <= 0;  //18 / 117 = 0
    16'b00010010_01110110 : OUT <= 0;  //18 / 118 = 0
    16'b00010010_01110111 : OUT <= 0;  //18 / 119 = 0
    16'b00010010_01111000 : OUT <= 0;  //18 / 120 = 0
    16'b00010010_01111001 : OUT <= 0;  //18 / 121 = 0
    16'b00010010_01111010 : OUT <= 0;  //18 / 122 = 0
    16'b00010010_01111011 : OUT <= 0;  //18 / 123 = 0
    16'b00010010_01111100 : OUT <= 0;  //18 / 124 = 0
    16'b00010010_01111101 : OUT <= 0;  //18 / 125 = 0
    16'b00010010_01111110 : OUT <= 0;  //18 / 126 = 0
    16'b00010010_01111111 : OUT <= 0;  //18 / 127 = 0
    16'b00010010_10000000 : OUT <= 0;  //18 / 128 = 0
    16'b00010010_10000001 : OUT <= 0;  //18 / 129 = 0
    16'b00010010_10000010 : OUT <= 0;  //18 / 130 = 0
    16'b00010010_10000011 : OUT <= 0;  //18 / 131 = 0
    16'b00010010_10000100 : OUT <= 0;  //18 / 132 = 0
    16'b00010010_10000101 : OUT <= 0;  //18 / 133 = 0
    16'b00010010_10000110 : OUT <= 0;  //18 / 134 = 0
    16'b00010010_10000111 : OUT <= 0;  //18 / 135 = 0
    16'b00010010_10001000 : OUT <= 0;  //18 / 136 = 0
    16'b00010010_10001001 : OUT <= 0;  //18 / 137 = 0
    16'b00010010_10001010 : OUT <= 0;  //18 / 138 = 0
    16'b00010010_10001011 : OUT <= 0;  //18 / 139 = 0
    16'b00010010_10001100 : OUT <= 0;  //18 / 140 = 0
    16'b00010010_10001101 : OUT <= 0;  //18 / 141 = 0
    16'b00010010_10001110 : OUT <= 0;  //18 / 142 = 0
    16'b00010010_10001111 : OUT <= 0;  //18 / 143 = 0
    16'b00010010_10010000 : OUT <= 0;  //18 / 144 = 0
    16'b00010010_10010001 : OUT <= 0;  //18 / 145 = 0
    16'b00010010_10010010 : OUT <= 0;  //18 / 146 = 0
    16'b00010010_10010011 : OUT <= 0;  //18 / 147 = 0
    16'b00010010_10010100 : OUT <= 0;  //18 / 148 = 0
    16'b00010010_10010101 : OUT <= 0;  //18 / 149 = 0
    16'b00010010_10010110 : OUT <= 0;  //18 / 150 = 0
    16'b00010010_10010111 : OUT <= 0;  //18 / 151 = 0
    16'b00010010_10011000 : OUT <= 0;  //18 / 152 = 0
    16'b00010010_10011001 : OUT <= 0;  //18 / 153 = 0
    16'b00010010_10011010 : OUT <= 0;  //18 / 154 = 0
    16'b00010010_10011011 : OUT <= 0;  //18 / 155 = 0
    16'b00010010_10011100 : OUT <= 0;  //18 / 156 = 0
    16'b00010010_10011101 : OUT <= 0;  //18 / 157 = 0
    16'b00010010_10011110 : OUT <= 0;  //18 / 158 = 0
    16'b00010010_10011111 : OUT <= 0;  //18 / 159 = 0
    16'b00010010_10100000 : OUT <= 0;  //18 / 160 = 0
    16'b00010010_10100001 : OUT <= 0;  //18 / 161 = 0
    16'b00010010_10100010 : OUT <= 0;  //18 / 162 = 0
    16'b00010010_10100011 : OUT <= 0;  //18 / 163 = 0
    16'b00010010_10100100 : OUT <= 0;  //18 / 164 = 0
    16'b00010010_10100101 : OUT <= 0;  //18 / 165 = 0
    16'b00010010_10100110 : OUT <= 0;  //18 / 166 = 0
    16'b00010010_10100111 : OUT <= 0;  //18 / 167 = 0
    16'b00010010_10101000 : OUT <= 0;  //18 / 168 = 0
    16'b00010010_10101001 : OUT <= 0;  //18 / 169 = 0
    16'b00010010_10101010 : OUT <= 0;  //18 / 170 = 0
    16'b00010010_10101011 : OUT <= 0;  //18 / 171 = 0
    16'b00010010_10101100 : OUT <= 0;  //18 / 172 = 0
    16'b00010010_10101101 : OUT <= 0;  //18 / 173 = 0
    16'b00010010_10101110 : OUT <= 0;  //18 / 174 = 0
    16'b00010010_10101111 : OUT <= 0;  //18 / 175 = 0
    16'b00010010_10110000 : OUT <= 0;  //18 / 176 = 0
    16'b00010010_10110001 : OUT <= 0;  //18 / 177 = 0
    16'b00010010_10110010 : OUT <= 0;  //18 / 178 = 0
    16'b00010010_10110011 : OUT <= 0;  //18 / 179 = 0
    16'b00010010_10110100 : OUT <= 0;  //18 / 180 = 0
    16'b00010010_10110101 : OUT <= 0;  //18 / 181 = 0
    16'b00010010_10110110 : OUT <= 0;  //18 / 182 = 0
    16'b00010010_10110111 : OUT <= 0;  //18 / 183 = 0
    16'b00010010_10111000 : OUT <= 0;  //18 / 184 = 0
    16'b00010010_10111001 : OUT <= 0;  //18 / 185 = 0
    16'b00010010_10111010 : OUT <= 0;  //18 / 186 = 0
    16'b00010010_10111011 : OUT <= 0;  //18 / 187 = 0
    16'b00010010_10111100 : OUT <= 0;  //18 / 188 = 0
    16'b00010010_10111101 : OUT <= 0;  //18 / 189 = 0
    16'b00010010_10111110 : OUT <= 0;  //18 / 190 = 0
    16'b00010010_10111111 : OUT <= 0;  //18 / 191 = 0
    16'b00010010_11000000 : OUT <= 0;  //18 / 192 = 0
    16'b00010010_11000001 : OUT <= 0;  //18 / 193 = 0
    16'b00010010_11000010 : OUT <= 0;  //18 / 194 = 0
    16'b00010010_11000011 : OUT <= 0;  //18 / 195 = 0
    16'b00010010_11000100 : OUT <= 0;  //18 / 196 = 0
    16'b00010010_11000101 : OUT <= 0;  //18 / 197 = 0
    16'b00010010_11000110 : OUT <= 0;  //18 / 198 = 0
    16'b00010010_11000111 : OUT <= 0;  //18 / 199 = 0
    16'b00010010_11001000 : OUT <= 0;  //18 / 200 = 0
    16'b00010010_11001001 : OUT <= 0;  //18 / 201 = 0
    16'b00010010_11001010 : OUT <= 0;  //18 / 202 = 0
    16'b00010010_11001011 : OUT <= 0;  //18 / 203 = 0
    16'b00010010_11001100 : OUT <= 0;  //18 / 204 = 0
    16'b00010010_11001101 : OUT <= 0;  //18 / 205 = 0
    16'b00010010_11001110 : OUT <= 0;  //18 / 206 = 0
    16'b00010010_11001111 : OUT <= 0;  //18 / 207 = 0
    16'b00010010_11010000 : OUT <= 0;  //18 / 208 = 0
    16'b00010010_11010001 : OUT <= 0;  //18 / 209 = 0
    16'b00010010_11010010 : OUT <= 0;  //18 / 210 = 0
    16'b00010010_11010011 : OUT <= 0;  //18 / 211 = 0
    16'b00010010_11010100 : OUT <= 0;  //18 / 212 = 0
    16'b00010010_11010101 : OUT <= 0;  //18 / 213 = 0
    16'b00010010_11010110 : OUT <= 0;  //18 / 214 = 0
    16'b00010010_11010111 : OUT <= 0;  //18 / 215 = 0
    16'b00010010_11011000 : OUT <= 0;  //18 / 216 = 0
    16'b00010010_11011001 : OUT <= 0;  //18 / 217 = 0
    16'b00010010_11011010 : OUT <= 0;  //18 / 218 = 0
    16'b00010010_11011011 : OUT <= 0;  //18 / 219 = 0
    16'b00010010_11011100 : OUT <= 0;  //18 / 220 = 0
    16'b00010010_11011101 : OUT <= 0;  //18 / 221 = 0
    16'b00010010_11011110 : OUT <= 0;  //18 / 222 = 0
    16'b00010010_11011111 : OUT <= 0;  //18 / 223 = 0
    16'b00010010_11100000 : OUT <= 0;  //18 / 224 = 0
    16'b00010010_11100001 : OUT <= 0;  //18 / 225 = 0
    16'b00010010_11100010 : OUT <= 0;  //18 / 226 = 0
    16'b00010010_11100011 : OUT <= 0;  //18 / 227 = 0
    16'b00010010_11100100 : OUT <= 0;  //18 / 228 = 0
    16'b00010010_11100101 : OUT <= 0;  //18 / 229 = 0
    16'b00010010_11100110 : OUT <= 0;  //18 / 230 = 0
    16'b00010010_11100111 : OUT <= 0;  //18 / 231 = 0
    16'b00010010_11101000 : OUT <= 0;  //18 / 232 = 0
    16'b00010010_11101001 : OUT <= 0;  //18 / 233 = 0
    16'b00010010_11101010 : OUT <= 0;  //18 / 234 = 0
    16'b00010010_11101011 : OUT <= 0;  //18 / 235 = 0
    16'b00010010_11101100 : OUT <= 0;  //18 / 236 = 0
    16'b00010010_11101101 : OUT <= 0;  //18 / 237 = 0
    16'b00010010_11101110 : OUT <= 0;  //18 / 238 = 0
    16'b00010010_11101111 : OUT <= 0;  //18 / 239 = 0
    16'b00010010_11110000 : OUT <= 0;  //18 / 240 = 0
    16'b00010010_11110001 : OUT <= 0;  //18 / 241 = 0
    16'b00010010_11110010 : OUT <= 0;  //18 / 242 = 0
    16'b00010010_11110011 : OUT <= 0;  //18 / 243 = 0
    16'b00010010_11110100 : OUT <= 0;  //18 / 244 = 0
    16'b00010010_11110101 : OUT <= 0;  //18 / 245 = 0
    16'b00010010_11110110 : OUT <= 0;  //18 / 246 = 0
    16'b00010010_11110111 : OUT <= 0;  //18 / 247 = 0
    16'b00010010_11111000 : OUT <= 0;  //18 / 248 = 0
    16'b00010010_11111001 : OUT <= 0;  //18 / 249 = 0
    16'b00010010_11111010 : OUT <= 0;  //18 / 250 = 0
    16'b00010010_11111011 : OUT <= 0;  //18 / 251 = 0
    16'b00010010_11111100 : OUT <= 0;  //18 / 252 = 0
    16'b00010010_11111101 : OUT <= 0;  //18 / 253 = 0
    16'b00010010_11111110 : OUT <= 0;  //18 / 254 = 0
    16'b00010010_11111111 : OUT <= 0;  //18 / 255 = 0
    16'b00010011_00000000 : OUT <= 0;  //19 / 0 = 0
    16'b00010011_00000001 : OUT <= 19;  //19 / 1 = 19
    16'b00010011_00000010 : OUT <= 9;  //19 / 2 = 9
    16'b00010011_00000011 : OUT <= 6;  //19 / 3 = 6
    16'b00010011_00000100 : OUT <= 4;  //19 / 4 = 4
    16'b00010011_00000101 : OUT <= 3;  //19 / 5 = 3
    16'b00010011_00000110 : OUT <= 3;  //19 / 6 = 3
    16'b00010011_00000111 : OUT <= 2;  //19 / 7 = 2
    16'b00010011_00001000 : OUT <= 2;  //19 / 8 = 2
    16'b00010011_00001001 : OUT <= 2;  //19 / 9 = 2
    16'b00010011_00001010 : OUT <= 1;  //19 / 10 = 1
    16'b00010011_00001011 : OUT <= 1;  //19 / 11 = 1
    16'b00010011_00001100 : OUT <= 1;  //19 / 12 = 1
    16'b00010011_00001101 : OUT <= 1;  //19 / 13 = 1
    16'b00010011_00001110 : OUT <= 1;  //19 / 14 = 1
    16'b00010011_00001111 : OUT <= 1;  //19 / 15 = 1
    16'b00010011_00010000 : OUT <= 1;  //19 / 16 = 1
    16'b00010011_00010001 : OUT <= 1;  //19 / 17 = 1
    16'b00010011_00010010 : OUT <= 1;  //19 / 18 = 1
    16'b00010011_00010011 : OUT <= 1;  //19 / 19 = 1
    16'b00010011_00010100 : OUT <= 0;  //19 / 20 = 0
    16'b00010011_00010101 : OUT <= 0;  //19 / 21 = 0
    16'b00010011_00010110 : OUT <= 0;  //19 / 22 = 0
    16'b00010011_00010111 : OUT <= 0;  //19 / 23 = 0
    16'b00010011_00011000 : OUT <= 0;  //19 / 24 = 0
    16'b00010011_00011001 : OUT <= 0;  //19 / 25 = 0
    16'b00010011_00011010 : OUT <= 0;  //19 / 26 = 0
    16'b00010011_00011011 : OUT <= 0;  //19 / 27 = 0
    16'b00010011_00011100 : OUT <= 0;  //19 / 28 = 0
    16'b00010011_00011101 : OUT <= 0;  //19 / 29 = 0
    16'b00010011_00011110 : OUT <= 0;  //19 / 30 = 0
    16'b00010011_00011111 : OUT <= 0;  //19 / 31 = 0
    16'b00010011_00100000 : OUT <= 0;  //19 / 32 = 0
    16'b00010011_00100001 : OUT <= 0;  //19 / 33 = 0
    16'b00010011_00100010 : OUT <= 0;  //19 / 34 = 0
    16'b00010011_00100011 : OUT <= 0;  //19 / 35 = 0
    16'b00010011_00100100 : OUT <= 0;  //19 / 36 = 0
    16'b00010011_00100101 : OUT <= 0;  //19 / 37 = 0
    16'b00010011_00100110 : OUT <= 0;  //19 / 38 = 0
    16'b00010011_00100111 : OUT <= 0;  //19 / 39 = 0
    16'b00010011_00101000 : OUT <= 0;  //19 / 40 = 0
    16'b00010011_00101001 : OUT <= 0;  //19 / 41 = 0
    16'b00010011_00101010 : OUT <= 0;  //19 / 42 = 0
    16'b00010011_00101011 : OUT <= 0;  //19 / 43 = 0
    16'b00010011_00101100 : OUT <= 0;  //19 / 44 = 0
    16'b00010011_00101101 : OUT <= 0;  //19 / 45 = 0
    16'b00010011_00101110 : OUT <= 0;  //19 / 46 = 0
    16'b00010011_00101111 : OUT <= 0;  //19 / 47 = 0
    16'b00010011_00110000 : OUT <= 0;  //19 / 48 = 0
    16'b00010011_00110001 : OUT <= 0;  //19 / 49 = 0
    16'b00010011_00110010 : OUT <= 0;  //19 / 50 = 0
    16'b00010011_00110011 : OUT <= 0;  //19 / 51 = 0
    16'b00010011_00110100 : OUT <= 0;  //19 / 52 = 0
    16'b00010011_00110101 : OUT <= 0;  //19 / 53 = 0
    16'b00010011_00110110 : OUT <= 0;  //19 / 54 = 0
    16'b00010011_00110111 : OUT <= 0;  //19 / 55 = 0
    16'b00010011_00111000 : OUT <= 0;  //19 / 56 = 0
    16'b00010011_00111001 : OUT <= 0;  //19 / 57 = 0
    16'b00010011_00111010 : OUT <= 0;  //19 / 58 = 0
    16'b00010011_00111011 : OUT <= 0;  //19 / 59 = 0
    16'b00010011_00111100 : OUT <= 0;  //19 / 60 = 0
    16'b00010011_00111101 : OUT <= 0;  //19 / 61 = 0
    16'b00010011_00111110 : OUT <= 0;  //19 / 62 = 0
    16'b00010011_00111111 : OUT <= 0;  //19 / 63 = 0
    16'b00010011_01000000 : OUT <= 0;  //19 / 64 = 0
    16'b00010011_01000001 : OUT <= 0;  //19 / 65 = 0
    16'b00010011_01000010 : OUT <= 0;  //19 / 66 = 0
    16'b00010011_01000011 : OUT <= 0;  //19 / 67 = 0
    16'b00010011_01000100 : OUT <= 0;  //19 / 68 = 0
    16'b00010011_01000101 : OUT <= 0;  //19 / 69 = 0
    16'b00010011_01000110 : OUT <= 0;  //19 / 70 = 0
    16'b00010011_01000111 : OUT <= 0;  //19 / 71 = 0
    16'b00010011_01001000 : OUT <= 0;  //19 / 72 = 0
    16'b00010011_01001001 : OUT <= 0;  //19 / 73 = 0
    16'b00010011_01001010 : OUT <= 0;  //19 / 74 = 0
    16'b00010011_01001011 : OUT <= 0;  //19 / 75 = 0
    16'b00010011_01001100 : OUT <= 0;  //19 / 76 = 0
    16'b00010011_01001101 : OUT <= 0;  //19 / 77 = 0
    16'b00010011_01001110 : OUT <= 0;  //19 / 78 = 0
    16'b00010011_01001111 : OUT <= 0;  //19 / 79 = 0
    16'b00010011_01010000 : OUT <= 0;  //19 / 80 = 0
    16'b00010011_01010001 : OUT <= 0;  //19 / 81 = 0
    16'b00010011_01010010 : OUT <= 0;  //19 / 82 = 0
    16'b00010011_01010011 : OUT <= 0;  //19 / 83 = 0
    16'b00010011_01010100 : OUT <= 0;  //19 / 84 = 0
    16'b00010011_01010101 : OUT <= 0;  //19 / 85 = 0
    16'b00010011_01010110 : OUT <= 0;  //19 / 86 = 0
    16'b00010011_01010111 : OUT <= 0;  //19 / 87 = 0
    16'b00010011_01011000 : OUT <= 0;  //19 / 88 = 0
    16'b00010011_01011001 : OUT <= 0;  //19 / 89 = 0
    16'b00010011_01011010 : OUT <= 0;  //19 / 90 = 0
    16'b00010011_01011011 : OUT <= 0;  //19 / 91 = 0
    16'b00010011_01011100 : OUT <= 0;  //19 / 92 = 0
    16'b00010011_01011101 : OUT <= 0;  //19 / 93 = 0
    16'b00010011_01011110 : OUT <= 0;  //19 / 94 = 0
    16'b00010011_01011111 : OUT <= 0;  //19 / 95 = 0
    16'b00010011_01100000 : OUT <= 0;  //19 / 96 = 0
    16'b00010011_01100001 : OUT <= 0;  //19 / 97 = 0
    16'b00010011_01100010 : OUT <= 0;  //19 / 98 = 0
    16'b00010011_01100011 : OUT <= 0;  //19 / 99 = 0
    16'b00010011_01100100 : OUT <= 0;  //19 / 100 = 0
    16'b00010011_01100101 : OUT <= 0;  //19 / 101 = 0
    16'b00010011_01100110 : OUT <= 0;  //19 / 102 = 0
    16'b00010011_01100111 : OUT <= 0;  //19 / 103 = 0
    16'b00010011_01101000 : OUT <= 0;  //19 / 104 = 0
    16'b00010011_01101001 : OUT <= 0;  //19 / 105 = 0
    16'b00010011_01101010 : OUT <= 0;  //19 / 106 = 0
    16'b00010011_01101011 : OUT <= 0;  //19 / 107 = 0
    16'b00010011_01101100 : OUT <= 0;  //19 / 108 = 0
    16'b00010011_01101101 : OUT <= 0;  //19 / 109 = 0
    16'b00010011_01101110 : OUT <= 0;  //19 / 110 = 0
    16'b00010011_01101111 : OUT <= 0;  //19 / 111 = 0
    16'b00010011_01110000 : OUT <= 0;  //19 / 112 = 0
    16'b00010011_01110001 : OUT <= 0;  //19 / 113 = 0
    16'b00010011_01110010 : OUT <= 0;  //19 / 114 = 0
    16'b00010011_01110011 : OUT <= 0;  //19 / 115 = 0
    16'b00010011_01110100 : OUT <= 0;  //19 / 116 = 0
    16'b00010011_01110101 : OUT <= 0;  //19 / 117 = 0
    16'b00010011_01110110 : OUT <= 0;  //19 / 118 = 0
    16'b00010011_01110111 : OUT <= 0;  //19 / 119 = 0
    16'b00010011_01111000 : OUT <= 0;  //19 / 120 = 0
    16'b00010011_01111001 : OUT <= 0;  //19 / 121 = 0
    16'b00010011_01111010 : OUT <= 0;  //19 / 122 = 0
    16'b00010011_01111011 : OUT <= 0;  //19 / 123 = 0
    16'b00010011_01111100 : OUT <= 0;  //19 / 124 = 0
    16'b00010011_01111101 : OUT <= 0;  //19 / 125 = 0
    16'b00010011_01111110 : OUT <= 0;  //19 / 126 = 0
    16'b00010011_01111111 : OUT <= 0;  //19 / 127 = 0
    16'b00010011_10000000 : OUT <= 0;  //19 / 128 = 0
    16'b00010011_10000001 : OUT <= 0;  //19 / 129 = 0
    16'b00010011_10000010 : OUT <= 0;  //19 / 130 = 0
    16'b00010011_10000011 : OUT <= 0;  //19 / 131 = 0
    16'b00010011_10000100 : OUT <= 0;  //19 / 132 = 0
    16'b00010011_10000101 : OUT <= 0;  //19 / 133 = 0
    16'b00010011_10000110 : OUT <= 0;  //19 / 134 = 0
    16'b00010011_10000111 : OUT <= 0;  //19 / 135 = 0
    16'b00010011_10001000 : OUT <= 0;  //19 / 136 = 0
    16'b00010011_10001001 : OUT <= 0;  //19 / 137 = 0
    16'b00010011_10001010 : OUT <= 0;  //19 / 138 = 0
    16'b00010011_10001011 : OUT <= 0;  //19 / 139 = 0
    16'b00010011_10001100 : OUT <= 0;  //19 / 140 = 0
    16'b00010011_10001101 : OUT <= 0;  //19 / 141 = 0
    16'b00010011_10001110 : OUT <= 0;  //19 / 142 = 0
    16'b00010011_10001111 : OUT <= 0;  //19 / 143 = 0
    16'b00010011_10010000 : OUT <= 0;  //19 / 144 = 0
    16'b00010011_10010001 : OUT <= 0;  //19 / 145 = 0
    16'b00010011_10010010 : OUT <= 0;  //19 / 146 = 0
    16'b00010011_10010011 : OUT <= 0;  //19 / 147 = 0
    16'b00010011_10010100 : OUT <= 0;  //19 / 148 = 0
    16'b00010011_10010101 : OUT <= 0;  //19 / 149 = 0
    16'b00010011_10010110 : OUT <= 0;  //19 / 150 = 0
    16'b00010011_10010111 : OUT <= 0;  //19 / 151 = 0
    16'b00010011_10011000 : OUT <= 0;  //19 / 152 = 0
    16'b00010011_10011001 : OUT <= 0;  //19 / 153 = 0
    16'b00010011_10011010 : OUT <= 0;  //19 / 154 = 0
    16'b00010011_10011011 : OUT <= 0;  //19 / 155 = 0
    16'b00010011_10011100 : OUT <= 0;  //19 / 156 = 0
    16'b00010011_10011101 : OUT <= 0;  //19 / 157 = 0
    16'b00010011_10011110 : OUT <= 0;  //19 / 158 = 0
    16'b00010011_10011111 : OUT <= 0;  //19 / 159 = 0
    16'b00010011_10100000 : OUT <= 0;  //19 / 160 = 0
    16'b00010011_10100001 : OUT <= 0;  //19 / 161 = 0
    16'b00010011_10100010 : OUT <= 0;  //19 / 162 = 0
    16'b00010011_10100011 : OUT <= 0;  //19 / 163 = 0
    16'b00010011_10100100 : OUT <= 0;  //19 / 164 = 0
    16'b00010011_10100101 : OUT <= 0;  //19 / 165 = 0
    16'b00010011_10100110 : OUT <= 0;  //19 / 166 = 0
    16'b00010011_10100111 : OUT <= 0;  //19 / 167 = 0
    16'b00010011_10101000 : OUT <= 0;  //19 / 168 = 0
    16'b00010011_10101001 : OUT <= 0;  //19 / 169 = 0
    16'b00010011_10101010 : OUT <= 0;  //19 / 170 = 0
    16'b00010011_10101011 : OUT <= 0;  //19 / 171 = 0
    16'b00010011_10101100 : OUT <= 0;  //19 / 172 = 0
    16'b00010011_10101101 : OUT <= 0;  //19 / 173 = 0
    16'b00010011_10101110 : OUT <= 0;  //19 / 174 = 0
    16'b00010011_10101111 : OUT <= 0;  //19 / 175 = 0
    16'b00010011_10110000 : OUT <= 0;  //19 / 176 = 0
    16'b00010011_10110001 : OUT <= 0;  //19 / 177 = 0
    16'b00010011_10110010 : OUT <= 0;  //19 / 178 = 0
    16'b00010011_10110011 : OUT <= 0;  //19 / 179 = 0
    16'b00010011_10110100 : OUT <= 0;  //19 / 180 = 0
    16'b00010011_10110101 : OUT <= 0;  //19 / 181 = 0
    16'b00010011_10110110 : OUT <= 0;  //19 / 182 = 0
    16'b00010011_10110111 : OUT <= 0;  //19 / 183 = 0
    16'b00010011_10111000 : OUT <= 0;  //19 / 184 = 0
    16'b00010011_10111001 : OUT <= 0;  //19 / 185 = 0
    16'b00010011_10111010 : OUT <= 0;  //19 / 186 = 0
    16'b00010011_10111011 : OUT <= 0;  //19 / 187 = 0
    16'b00010011_10111100 : OUT <= 0;  //19 / 188 = 0
    16'b00010011_10111101 : OUT <= 0;  //19 / 189 = 0
    16'b00010011_10111110 : OUT <= 0;  //19 / 190 = 0
    16'b00010011_10111111 : OUT <= 0;  //19 / 191 = 0
    16'b00010011_11000000 : OUT <= 0;  //19 / 192 = 0
    16'b00010011_11000001 : OUT <= 0;  //19 / 193 = 0
    16'b00010011_11000010 : OUT <= 0;  //19 / 194 = 0
    16'b00010011_11000011 : OUT <= 0;  //19 / 195 = 0
    16'b00010011_11000100 : OUT <= 0;  //19 / 196 = 0
    16'b00010011_11000101 : OUT <= 0;  //19 / 197 = 0
    16'b00010011_11000110 : OUT <= 0;  //19 / 198 = 0
    16'b00010011_11000111 : OUT <= 0;  //19 / 199 = 0
    16'b00010011_11001000 : OUT <= 0;  //19 / 200 = 0
    16'b00010011_11001001 : OUT <= 0;  //19 / 201 = 0
    16'b00010011_11001010 : OUT <= 0;  //19 / 202 = 0
    16'b00010011_11001011 : OUT <= 0;  //19 / 203 = 0
    16'b00010011_11001100 : OUT <= 0;  //19 / 204 = 0
    16'b00010011_11001101 : OUT <= 0;  //19 / 205 = 0
    16'b00010011_11001110 : OUT <= 0;  //19 / 206 = 0
    16'b00010011_11001111 : OUT <= 0;  //19 / 207 = 0
    16'b00010011_11010000 : OUT <= 0;  //19 / 208 = 0
    16'b00010011_11010001 : OUT <= 0;  //19 / 209 = 0
    16'b00010011_11010010 : OUT <= 0;  //19 / 210 = 0
    16'b00010011_11010011 : OUT <= 0;  //19 / 211 = 0
    16'b00010011_11010100 : OUT <= 0;  //19 / 212 = 0
    16'b00010011_11010101 : OUT <= 0;  //19 / 213 = 0
    16'b00010011_11010110 : OUT <= 0;  //19 / 214 = 0
    16'b00010011_11010111 : OUT <= 0;  //19 / 215 = 0
    16'b00010011_11011000 : OUT <= 0;  //19 / 216 = 0
    16'b00010011_11011001 : OUT <= 0;  //19 / 217 = 0
    16'b00010011_11011010 : OUT <= 0;  //19 / 218 = 0
    16'b00010011_11011011 : OUT <= 0;  //19 / 219 = 0
    16'b00010011_11011100 : OUT <= 0;  //19 / 220 = 0
    16'b00010011_11011101 : OUT <= 0;  //19 / 221 = 0
    16'b00010011_11011110 : OUT <= 0;  //19 / 222 = 0
    16'b00010011_11011111 : OUT <= 0;  //19 / 223 = 0
    16'b00010011_11100000 : OUT <= 0;  //19 / 224 = 0
    16'b00010011_11100001 : OUT <= 0;  //19 / 225 = 0
    16'b00010011_11100010 : OUT <= 0;  //19 / 226 = 0
    16'b00010011_11100011 : OUT <= 0;  //19 / 227 = 0
    16'b00010011_11100100 : OUT <= 0;  //19 / 228 = 0
    16'b00010011_11100101 : OUT <= 0;  //19 / 229 = 0
    16'b00010011_11100110 : OUT <= 0;  //19 / 230 = 0
    16'b00010011_11100111 : OUT <= 0;  //19 / 231 = 0
    16'b00010011_11101000 : OUT <= 0;  //19 / 232 = 0
    16'b00010011_11101001 : OUT <= 0;  //19 / 233 = 0
    16'b00010011_11101010 : OUT <= 0;  //19 / 234 = 0
    16'b00010011_11101011 : OUT <= 0;  //19 / 235 = 0
    16'b00010011_11101100 : OUT <= 0;  //19 / 236 = 0
    16'b00010011_11101101 : OUT <= 0;  //19 / 237 = 0
    16'b00010011_11101110 : OUT <= 0;  //19 / 238 = 0
    16'b00010011_11101111 : OUT <= 0;  //19 / 239 = 0
    16'b00010011_11110000 : OUT <= 0;  //19 / 240 = 0
    16'b00010011_11110001 : OUT <= 0;  //19 / 241 = 0
    16'b00010011_11110010 : OUT <= 0;  //19 / 242 = 0
    16'b00010011_11110011 : OUT <= 0;  //19 / 243 = 0
    16'b00010011_11110100 : OUT <= 0;  //19 / 244 = 0
    16'b00010011_11110101 : OUT <= 0;  //19 / 245 = 0
    16'b00010011_11110110 : OUT <= 0;  //19 / 246 = 0
    16'b00010011_11110111 : OUT <= 0;  //19 / 247 = 0
    16'b00010011_11111000 : OUT <= 0;  //19 / 248 = 0
    16'b00010011_11111001 : OUT <= 0;  //19 / 249 = 0
    16'b00010011_11111010 : OUT <= 0;  //19 / 250 = 0
    16'b00010011_11111011 : OUT <= 0;  //19 / 251 = 0
    16'b00010011_11111100 : OUT <= 0;  //19 / 252 = 0
    16'b00010011_11111101 : OUT <= 0;  //19 / 253 = 0
    16'b00010011_11111110 : OUT <= 0;  //19 / 254 = 0
    16'b00010011_11111111 : OUT <= 0;  //19 / 255 = 0
    16'b00010100_00000000 : OUT <= 0;  //20 / 0 = 0
    16'b00010100_00000001 : OUT <= 20;  //20 / 1 = 20
    16'b00010100_00000010 : OUT <= 10;  //20 / 2 = 10
    16'b00010100_00000011 : OUT <= 6;  //20 / 3 = 6
    16'b00010100_00000100 : OUT <= 5;  //20 / 4 = 5
    16'b00010100_00000101 : OUT <= 4;  //20 / 5 = 4
    16'b00010100_00000110 : OUT <= 3;  //20 / 6 = 3
    16'b00010100_00000111 : OUT <= 2;  //20 / 7 = 2
    16'b00010100_00001000 : OUT <= 2;  //20 / 8 = 2
    16'b00010100_00001001 : OUT <= 2;  //20 / 9 = 2
    16'b00010100_00001010 : OUT <= 2;  //20 / 10 = 2
    16'b00010100_00001011 : OUT <= 1;  //20 / 11 = 1
    16'b00010100_00001100 : OUT <= 1;  //20 / 12 = 1
    16'b00010100_00001101 : OUT <= 1;  //20 / 13 = 1
    16'b00010100_00001110 : OUT <= 1;  //20 / 14 = 1
    16'b00010100_00001111 : OUT <= 1;  //20 / 15 = 1
    16'b00010100_00010000 : OUT <= 1;  //20 / 16 = 1
    16'b00010100_00010001 : OUT <= 1;  //20 / 17 = 1
    16'b00010100_00010010 : OUT <= 1;  //20 / 18 = 1
    16'b00010100_00010011 : OUT <= 1;  //20 / 19 = 1
    16'b00010100_00010100 : OUT <= 1;  //20 / 20 = 1
    16'b00010100_00010101 : OUT <= 0;  //20 / 21 = 0
    16'b00010100_00010110 : OUT <= 0;  //20 / 22 = 0
    16'b00010100_00010111 : OUT <= 0;  //20 / 23 = 0
    16'b00010100_00011000 : OUT <= 0;  //20 / 24 = 0
    16'b00010100_00011001 : OUT <= 0;  //20 / 25 = 0
    16'b00010100_00011010 : OUT <= 0;  //20 / 26 = 0
    16'b00010100_00011011 : OUT <= 0;  //20 / 27 = 0
    16'b00010100_00011100 : OUT <= 0;  //20 / 28 = 0
    16'b00010100_00011101 : OUT <= 0;  //20 / 29 = 0
    16'b00010100_00011110 : OUT <= 0;  //20 / 30 = 0
    16'b00010100_00011111 : OUT <= 0;  //20 / 31 = 0
    16'b00010100_00100000 : OUT <= 0;  //20 / 32 = 0
    16'b00010100_00100001 : OUT <= 0;  //20 / 33 = 0
    16'b00010100_00100010 : OUT <= 0;  //20 / 34 = 0
    16'b00010100_00100011 : OUT <= 0;  //20 / 35 = 0
    16'b00010100_00100100 : OUT <= 0;  //20 / 36 = 0
    16'b00010100_00100101 : OUT <= 0;  //20 / 37 = 0
    16'b00010100_00100110 : OUT <= 0;  //20 / 38 = 0
    16'b00010100_00100111 : OUT <= 0;  //20 / 39 = 0
    16'b00010100_00101000 : OUT <= 0;  //20 / 40 = 0
    16'b00010100_00101001 : OUT <= 0;  //20 / 41 = 0
    16'b00010100_00101010 : OUT <= 0;  //20 / 42 = 0
    16'b00010100_00101011 : OUT <= 0;  //20 / 43 = 0
    16'b00010100_00101100 : OUT <= 0;  //20 / 44 = 0
    16'b00010100_00101101 : OUT <= 0;  //20 / 45 = 0
    16'b00010100_00101110 : OUT <= 0;  //20 / 46 = 0
    16'b00010100_00101111 : OUT <= 0;  //20 / 47 = 0
    16'b00010100_00110000 : OUT <= 0;  //20 / 48 = 0
    16'b00010100_00110001 : OUT <= 0;  //20 / 49 = 0
    16'b00010100_00110010 : OUT <= 0;  //20 / 50 = 0
    16'b00010100_00110011 : OUT <= 0;  //20 / 51 = 0
    16'b00010100_00110100 : OUT <= 0;  //20 / 52 = 0
    16'b00010100_00110101 : OUT <= 0;  //20 / 53 = 0
    16'b00010100_00110110 : OUT <= 0;  //20 / 54 = 0
    16'b00010100_00110111 : OUT <= 0;  //20 / 55 = 0
    16'b00010100_00111000 : OUT <= 0;  //20 / 56 = 0
    16'b00010100_00111001 : OUT <= 0;  //20 / 57 = 0
    16'b00010100_00111010 : OUT <= 0;  //20 / 58 = 0
    16'b00010100_00111011 : OUT <= 0;  //20 / 59 = 0
    16'b00010100_00111100 : OUT <= 0;  //20 / 60 = 0
    16'b00010100_00111101 : OUT <= 0;  //20 / 61 = 0
    16'b00010100_00111110 : OUT <= 0;  //20 / 62 = 0
    16'b00010100_00111111 : OUT <= 0;  //20 / 63 = 0
    16'b00010100_01000000 : OUT <= 0;  //20 / 64 = 0
    16'b00010100_01000001 : OUT <= 0;  //20 / 65 = 0
    16'b00010100_01000010 : OUT <= 0;  //20 / 66 = 0
    16'b00010100_01000011 : OUT <= 0;  //20 / 67 = 0
    16'b00010100_01000100 : OUT <= 0;  //20 / 68 = 0
    16'b00010100_01000101 : OUT <= 0;  //20 / 69 = 0
    16'b00010100_01000110 : OUT <= 0;  //20 / 70 = 0
    16'b00010100_01000111 : OUT <= 0;  //20 / 71 = 0
    16'b00010100_01001000 : OUT <= 0;  //20 / 72 = 0
    16'b00010100_01001001 : OUT <= 0;  //20 / 73 = 0
    16'b00010100_01001010 : OUT <= 0;  //20 / 74 = 0
    16'b00010100_01001011 : OUT <= 0;  //20 / 75 = 0
    16'b00010100_01001100 : OUT <= 0;  //20 / 76 = 0
    16'b00010100_01001101 : OUT <= 0;  //20 / 77 = 0
    16'b00010100_01001110 : OUT <= 0;  //20 / 78 = 0
    16'b00010100_01001111 : OUT <= 0;  //20 / 79 = 0
    16'b00010100_01010000 : OUT <= 0;  //20 / 80 = 0
    16'b00010100_01010001 : OUT <= 0;  //20 / 81 = 0
    16'b00010100_01010010 : OUT <= 0;  //20 / 82 = 0
    16'b00010100_01010011 : OUT <= 0;  //20 / 83 = 0
    16'b00010100_01010100 : OUT <= 0;  //20 / 84 = 0
    16'b00010100_01010101 : OUT <= 0;  //20 / 85 = 0
    16'b00010100_01010110 : OUT <= 0;  //20 / 86 = 0
    16'b00010100_01010111 : OUT <= 0;  //20 / 87 = 0
    16'b00010100_01011000 : OUT <= 0;  //20 / 88 = 0
    16'b00010100_01011001 : OUT <= 0;  //20 / 89 = 0
    16'b00010100_01011010 : OUT <= 0;  //20 / 90 = 0
    16'b00010100_01011011 : OUT <= 0;  //20 / 91 = 0
    16'b00010100_01011100 : OUT <= 0;  //20 / 92 = 0
    16'b00010100_01011101 : OUT <= 0;  //20 / 93 = 0
    16'b00010100_01011110 : OUT <= 0;  //20 / 94 = 0
    16'b00010100_01011111 : OUT <= 0;  //20 / 95 = 0
    16'b00010100_01100000 : OUT <= 0;  //20 / 96 = 0
    16'b00010100_01100001 : OUT <= 0;  //20 / 97 = 0
    16'b00010100_01100010 : OUT <= 0;  //20 / 98 = 0
    16'b00010100_01100011 : OUT <= 0;  //20 / 99 = 0
    16'b00010100_01100100 : OUT <= 0;  //20 / 100 = 0
    16'b00010100_01100101 : OUT <= 0;  //20 / 101 = 0
    16'b00010100_01100110 : OUT <= 0;  //20 / 102 = 0
    16'b00010100_01100111 : OUT <= 0;  //20 / 103 = 0
    16'b00010100_01101000 : OUT <= 0;  //20 / 104 = 0
    16'b00010100_01101001 : OUT <= 0;  //20 / 105 = 0
    16'b00010100_01101010 : OUT <= 0;  //20 / 106 = 0
    16'b00010100_01101011 : OUT <= 0;  //20 / 107 = 0
    16'b00010100_01101100 : OUT <= 0;  //20 / 108 = 0
    16'b00010100_01101101 : OUT <= 0;  //20 / 109 = 0
    16'b00010100_01101110 : OUT <= 0;  //20 / 110 = 0
    16'b00010100_01101111 : OUT <= 0;  //20 / 111 = 0
    16'b00010100_01110000 : OUT <= 0;  //20 / 112 = 0
    16'b00010100_01110001 : OUT <= 0;  //20 / 113 = 0
    16'b00010100_01110010 : OUT <= 0;  //20 / 114 = 0
    16'b00010100_01110011 : OUT <= 0;  //20 / 115 = 0
    16'b00010100_01110100 : OUT <= 0;  //20 / 116 = 0
    16'b00010100_01110101 : OUT <= 0;  //20 / 117 = 0
    16'b00010100_01110110 : OUT <= 0;  //20 / 118 = 0
    16'b00010100_01110111 : OUT <= 0;  //20 / 119 = 0
    16'b00010100_01111000 : OUT <= 0;  //20 / 120 = 0
    16'b00010100_01111001 : OUT <= 0;  //20 / 121 = 0
    16'b00010100_01111010 : OUT <= 0;  //20 / 122 = 0
    16'b00010100_01111011 : OUT <= 0;  //20 / 123 = 0
    16'b00010100_01111100 : OUT <= 0;  //20 / 124 = 0
    16'b00010100_01111101 : OUT <= 0;  //20 / 125 = 0
    16'b00010100_01111110 : OUT <= 0;  //20 / 126 = 0
    16'b00010100_01111111 : OUT <= 0;  //20 / 127 = 0
    16'b00010100_10000000 : OUT <= 0;  //20 / 128 = 0
    16'b00010100_10000001 : OUT <= 0;  //20 / 129 = 0
    16'b00010100_10000010 : OUT <= 0;  //20 / 130 = 0
    16'b00010100_10000011 : OUT <= 0;  //20 / 131 = 0
    16'b00010100_10000100 : OUT <= 0;  //20 / 132 = 0
    16'b00010100_10000101 : OUT <= 0;  //20 / 133 = 0
    16'b00010100_10000110 : OUT <= 0;  //20 / 134 = 0
    16'b00010100_10000111 : OUT <= 0;  //20 / 135 = 0
    16'b00010100_10001000 : OUT <= 0;  //20 / 136 = 0
    16'b00010100_10001001 : OUT <= 0;  //20 / 137 = 0
    16'b00010100_10001010 : OUT <= 0;  //20 / 138 = 0
    16'b00010100_10001011 : OUT <= 0;  //20 / 139 = 0
    16'b00010100_10001100 : OUT <= 0;  //20 / 140 = 0
    16'b00010100_10001101 : OUT <= 0;  //20 / 141 = 0
    16'b00010100_10001110 : OUT <= 0;  //20 / 142 = 0
    16'b00010100_10001111 : OUT <= 0;  //20 / 143 = 0
    16'b00010100_10010000 : OUT <= 0;  //20 / 144 = 0
    16'b00010100_10010001 : OUT <= 0;  //20 / 145 = 0
    16'b00010100_10010010 : OUT <= 0;  //20 / 146 = 0
    16'b00010100_10010011 : OUT <= 0;  //20 / 147 = 0
    16'b00010100_10010100 : OUT <= 0;  //20 / 148 = 0
    16'b00010100_10010101 : OUT <= 0;  //20 / 149 = 0
    16'b00010100_10010110 : OUT <= 0;  //20 / 150 = 0
    16'b00010100_10010111 : OUT <= 0;  //20 / 151 = 0
    16'b00010100_10011000 : OUT <= 0;  //20 / 152 = 0
    16'b00010100_10011001 : OUT <= 0;  //20 / 153 = 0
    16'b00010100_10011010 : OUT <= 0;  //20 / 154 = 0
    16'b00010100_10011011 : OUT <= 0;  //20 / 155 = 0
    16'b00010100_10011100 : OUT <= 0;  //20 / 156 = 0
    16'b00010100_10011101 : OUT <= 0;  //20 / 157 = 0
    16'b00010100_10011110 : OUT <= 0;  //20 / 158 = 0
    16'b00010100_10011111 : OUT <= 0;  //20 / 159 = 0
    16'b00010100_10100000 : OUT <= 0;  //20 / 160 = 0
    16'b00010100_10100001 : OUT <= 0;  //20 / 161 = 0
    16'b00010100_10100010 : OUT <= 0;  //20 / 162 = 0
    16'b00010100_10100011 : OUT <= 0;  //20 / 163 = 0
    16'b00010100_10100100 : OUT <= 0;  //20 / 164 = 0
    16'b00010100_10100101 : OUT <= 0;  //20 / 165 = 0
    16'b00010100_10100110 : OUT <= 0;  //20 / 166 = 0
    16'b00010100_10100111 : OUT <= 0;  //20 / 167 = 0
    16'b00010100_10101000 : OUT <= 0;  //20 / 168 = 0
    16'b00010100_10101001 : OUT <= 0;  //20 / 169 = 0
    16'b00010100_10101010 : OUT <= 0;  //20 / 170 = 0
    16'b00010100_10101011 : OUT <= 0;  //20 / 171 = 0
    16'b00010100_10101100 : OUT <= 0;  //20 / 172 = 0
    16'b00010100_10101101 : OUT <= 0;  //20 / 173 = 0
    16'b00010100_10101110 : OUT <= 0;  //20 / 174 = 0
    16'b00010100_10101111 : OUT <= 0;  //20 / 175 = 0
    16'b00010100_10110000 : OUT <= 0;  //20 / 176 = 0
    16'b00010100_10110001 : OUT <= 0;  //20 / 177 = 0
    16'b00010100_10110010 : OUT <= 0;  //20 / 178 = 0
    16'b00010100_10110011 : OUT <= 0;  //20 / 179 = 0
    16'b00010100_10110100 : OUT <= 0;  //20 / 180 = 0
    16'b00010100_10110101 : OUT <= 0;  //20 / 181 = 0
    16'b00010100_10110110 : OUT <= 0;  //20 / 182 = 0
    16'b00010100_10110111 : OUT <= 0;  //20 / 183 = 0
    16'b00010100_10111000 : OUT <= 0;  //20 / 184 = 0
    16'b00010100_10111001 : OUT <= 0;  //20 / 185 = 0
    16'b00010100_10111010 : OUT <= 0;  //20 / 186 = 0
    16'b00010100_10111011 : OUT <= 0;  //20 / 187 = 0
    16'b00010100_10111100 : OUT <= 0;  //20 / 188 = 0
    16'b00010100_10111101 : OUT <= 0;  //20 / 189 = 0
    16'b00010100_10111110 : OUT <= 0;  //20 / 190 = 0
    16'b00010100_10111111 : OUT <= 0;  //20 / 191 = 0
    16'b00010100_11000000 : OUT <= 0;  //20 / 192 = 0
    16'b00010100_11000001 : OUT <= 0;  //20 / 193 = 0
    16'b00010100_11000010 : OUT <= 0;  //20 / 194 = 0
    16'b00010100_11000011 : OUT <= 0;  //20 / 195 = 0
    16'b00010100_11000100 : OUT <= 0;  //20 / 196 = 0
    16'b00010100_11000101 : OUT <= 0;  //20 / 197 = 0
    16'b00010100_11000110 : OUT <= 0;  //20 / 198 = 0
    16'b00010100_11000111 : OUT <= 0;  //20 / 199 = 0
    16'b00010100_11001000 : OUT <= 0;  //20 / 200 = 0
    16'b00010100_11001001 : OUT <= 0;  //20 / 201 = 0
    16'b00010100_11001010 : OUT <= 0;  //20 / 202 = 0
    16'b00010100_11001011 : OUT <= 0;  //20 / 203 = 0
    16'b00010100_11001100 : OUT <= 0;  //20 / 204 = 0
    16'b00010100_11001101 : OUT <= 0;  //20 / 205 = 0
    16'b00010100_11001110 : OUT <= 0;  //20 / 206 = 0
    16'b00010100_11001111 : OUT <= 0;  //20 / 207 = 0
    16'b00010100_11010000 : OUT <= 0;  //20 / 208 = 0
    16'b00010100_11010001 : OUT <= 0;  //20 / 209 = 0
    16'b00010100_11010010 : OUT <= 0;  //20 / 210 = 0
    16'b00010100_11010011 : OUT <= 0;  //20 / 211 = 0
    16'b00010100_11010100 : OUT <= 0;  //20 / 212 = 0
    16'b00010100_11010101 : OUT <= 0;  //20 / 213 = 0
    16'b00010100_11010110 : OUT <= 0;  //20 / 214 = 0
    16'b00010100_11010111 : OUT <= 0;  //20 / 215 = 0
    16'b00010100_11011000 : OUT <= 0;  //20 / 216 = 0
    16'b00010100_11011001 : OUT <= 0;  //20 / 217 = 0
    16'b00010100_11011010 : OUT <= 0;  //20 / 218 = 0
    16'b00010100_11011011 : OUT <= 0;  //20 / 219 = 0
    16'b00010100_11011100 : OUT <= 0;  //20 / 220 = 0
    16'b00010100_11011101 : OUT <= 0;  //20 / 221 = 0
    16'b00010100_11011110 : OUT <= 0;  //20 / 222 = 0
    16'b00010100_11011111 : OUT <= 0;  //20 / 223 = 0
    16'b00010100_11100000 : OUT <= 0;  //20 / 224 = 0
    16'b00010100_11100001 : OUT <= 0;  //20 / 225 = 0
    16'b00010100_11100010 : OUT <= 0;  //20 / 226 = 0
    16'b00010100_11100011 : OUT <= 0;  //20 / 227 = 0
    16'b00010100_11100100 : OUT <= 0;  //20 / 228 = 0
    16'b00010100_11100101 : OUT <= 0;  //20 / 229 = 0
    16'b00010100_11100110 : OUT <= 0;  //20 / 230 = 0
    16'b00010100_11100111 : OUT <= 0;  //20 / 231 = 0
    16'b00010100_11101000 : OUT <= 0;  //20 / 232 = 0
    16'b00010100_11101001 : OUT <= 0;  //20 / 233 = 0
    16'b00010100_11101010 : OUT <= 0;  //20 / 234 = 0
    16'b00010100_11101011 : OUT <= 0;  //20 / 235 = 0
    16'b00010100_11101100 : OUT <= 0;  //20 / 236 = 0
    16'b00010100_11101101 : OUT <= 0;  //20 / 237 = 0
    16'b00010100_11101110 : OUT <= 0;  //20 / 238 = 0
    16'b00010100_11101111 : OUT <= 0;  //20 / 239 = 0
    16'b00010100_11110000 : OUT <= 0;  //20 / 240 = 0
    16'b00010100_11110001 : OUT <= 0;  //20 / 241 = 0
    16'b00010100_11110010 : OUT <= 0;  //20 / 242 = 0
    16'b00010100_11110011 : OUT <= 0;  //20 / 243 = 0
    16'b00010100_11110100 : OUT <= 0;  //20 / 244 = 0
    16'b00010100_11110101 : OUT <= 0;  //20 / 245 = 0
    16'b00010100_11110110 : OUT <= 0;  //20 / 246 = 0
    16'b00010100_11110111 : OUT <= 0;  //20 / 247 = 0
    16'b00010100_11111000 : OUT <= 0;  //20 / 248 = 0
    16'b00010100_11111001 : OUT <= 0;  //20 / 249 = 0
    16'b00010100_11111010 : OUT <= 0;  //20 / 250 = 0
    16'b00010100_11111011 : OUT <= 0;  //20 / 251 = 0
    16'b00010100_11111100 : OUT <= 0;  //20 / 252 = 0
    16'b00010100_11111101 : OUT <= 0;  //20 / 253 = 0
    16'b00010100_11111110 : OUT <= 0;  //20 / 254 = 0
    16'b00010100_11111111 : OUT <= 0;  //20 / 255 = 0
    16'b00010101_00000000 : OUT <= 0;  //21 / 0 = 0
    16'b00010101_00000001 : OUT <= 21;  //21 / 1 = 21
    16'b00010101_00000010 : OUT <= 10;  //21 / 2 = 10
    16'b00010101_00000011 : OUT <= 7;  //21 / 3 = 7
    16'b00010101_00000100 : OUT <= 5;  //21 / 4 = 5
    16'b00010101_00000101 : OUT <= 4;  //21 / 5 = 4
    16'b00010101_00000110 : OUT <= 3;  //21 / 6 = 3
    16'b00010101_00000111 : OUT <= 3;  //21 / 7 = 3
    16'b00010101_00001000 : OUT <= 2;  //21 / 8 = 2
    16'b00010101_00001001 : OUT <= 2;  //21 / 9 = 2
    16'b00010101_00001010 : OUT <= 2;  //21 / 10 = 2
    16'b00010101_00001011 : OUT <= 1;  //21 / 11 = 1
    16'b00010101_00001100 : OUT <= 1;  //21 / 12 = 1
    16'b00010101_00001101 : OUT <= 1;  //21 / 13 = 1
    16'b00010101_00001110 : OUT <= 1;  //21 / 14 = 1
    16'b00010101_00001111 : OUT <= 1;  //21 / 15 = 1
    16'b00010101_00010000 : OUT <= 1;  //21 / 16 = 1
    16'b00010101_00010001 : OUT <= 1;  //21 / 17 = 1
    16'b00010101_00010010 : OUT <= 1;  //21 / 18 = 1
    16'b00010101_00010011 : OUT <= 1;  //21 / 19 = 1
    16'b00010101_00010100 : OUT <= 1;  //21 / 20 = 1
    16'b00010101_00010101 : OUT <= 1;  //21 / 21 = 1
    16'b00010101_00010110 : OUT <= 0;  //21 / 22 = 0
    16'b00010101_00010111 : OUT <= 0;  //21 / 23 = 0
    16'b00010101_00011000 : OUT <= 0;  //21 / 24 = 0
    16'b00010101_00011001 : OUT <= 0;  //21 / 25 = 0
    16'b00010101_00011010 : OUT <= 0;  //21 / 26 = 0
    16'b00010101_00011011 : OUT <= 0;  //21 / 27 = 0
    16'b00010101_00011100 : OUT <= 0;  //21 / 28 = 0
    16'b00010101_00011101 : OUT <= 0;  //21 / 29 = 0
    16'b00010101_00011110 : OUT <= 0;  //21 / 30 = 0
    16'b00010101_00011111 : OUT <= 0;  //21 / 31 = 0
    16'b00010101_00100000 : OUT <= 0;  //21 / 32 = 0
    16'b00010101_00100001 : OUT <= 0;  //21 / 33 = 0
    16'b00010101_00100010 : OUT <= 0;  //21 / 34 = 0
    16'b00010101_00100011 : OUT <= 0;  //21 / 35 = 0
    16'b00010101_00100100 : OUT <= 0;  //21 / 36 = 0
    16'b00010101_00100101 : OUT <= 0;  //21 / 37 = 0
    16'b00010101_00100110 : OUT <= 0;  //21 / 38 = 0
    16'b00010101_00100111 : OUT <= 0;  //21 / 39 = 0
    16'b00010101_00101000 : OUT <= 0;  //21 / 40 = 0
    16'b00010101_00101001 : OUT <= 0;  //21 / 41 = 0
    16'b00010101_00101010 : OUT <= 0;  //21 / 42 = 0
    16'b00010101_00101011 : OUT <= 0;  //21 / 43 = 0
    16'b00010101_00101100 : OUT <= 0;  //21 / 44 = 0
    16'b00010101_00101101 : OUT <= 0;  //21 / 45 = 0
    16'b00010101_00101110 : OUT <= 0;  //21 / 46 = 0
    16'b00010101_00101111 : OUT <= 0;  //21 / 47 = 0
    16'b00010101_00110000 : OUT <= 0;  //21 / 48 = 0
    16'b00010101_00110001 : OUT <= 0;  //21 / 49 = 0
    16'b00010101_00110010 : OUT <= 0;  //21 / 50 = 0
    16'b00010101_00110011 : OUT <= 0;  //21 / 51 = 0
    16'b00010101_00110100 : OUT <= 0;  //21 / 52 = 0
    16'b00010101_00110101 : OUT <= 0;  //21 / 53 = 0
    16'b00010101_00110110 : OUT <= 0;  //21 / 54 = 0
    16'b00010101_00110111 : OUT <= 0;  //21 / 55 = 0
    16'b00010101_00111000 : OUT <= 0;  //21 / 56 = 0
    16'b00010101_00111001 : OUT <= 0;  //21 / 57 = 0
    16'b00010101_00111010 : OUT <= 0;  //21 / 58 = 0
    16'b00010101_00111011 : OUT <= 0;  //21 / 59 = 0
    16'b00010101_00111100 : OUT <= 0;  //21 / 60 = 0
    16'b00010101_00111101 : OUT <= 0;  //21 / 61 = 0
    16'b00010101_00111110 : OUT <= 0;  //21 / 62 = 0
    16'b00010101_00111111 : OUT <= 0;  //21 / 63 = 0
    16'b00010101_01000000 : OUT <= 0;  //21 / 64 = 0
    16'b00010101_01000001 : OUT <= 0;  //21 / 65 = 0
    16'b00010101_01000010 : OUT <= 0;  //21 / 66 = 0
    16'b00010101_01000011 : OUT <= 0;  //21 / 67 = 0
    16'b00010101_01000100 : OUT <= 0;  //21 / 68 = 0
    16'b00010101_01000101 : OUT <= 0;  //21 / 69 = 0
    16'b00010101_01000110 : OUT <= 0;  //21 / 70 = 0
    16'b00010101_01000111 : OUT <= 0;  //21 / 71 = 0
    16'b00010101_01001000 : OUT <= 0;  //21 / 72 = 0
    16'b00010101_01001001 : OUT <= 0;  //21 / 73 = 0
    16'b00010101_01001010 : OUT <= 0;  //21 / 74 = 0
    16'b00010101_01001011 : OUT <= 0;  //21 / 75 = 0
    16'b00010101_01001100 : OUT <= 0;  //21 / 76 = 0
    16'b00010101_01001101 : OUT <= 0;  //21 / 77 = 0
    16'b00010101_01001110 : OUT <= 0;  //21 / 78 = 0
    16'b00010101_01001111 : OUT <= 0;  //21 / 79 = 0
    16'b00010101_01010000 : OUT <= 0;  //21 / 80 = 0
    16'b00010101_01010001 : OUT <= 0;  //21 / 81 = 0
    16'b00010101_01010010 : OUT <= 0;  //21 / 82 = 0
    16'b00010101_01010011 : OUT <= 0;  //21 / 83 = 0
    16'b00010101_01010100 : OUT <= 0;  //21 / 84 = 0
    16'b00010101_01010101 : OUT <= 0;  //21 / 85 = 0
    16'b00010101_01010110 : OUT <= 0;  //21 / 86 = 0
    16'b00010101_01010111 : OUT <= 0;  //21 / 87 = 0
    16'b00010101_01011000 : OUT <= 0;  //21 / 88 = 0
    16'b00010101_01011001 : OUT <= 0;  //21 / 89 = 0
    16'b00010101_01011010 : OUT <= 0;  //21 / 90 = 0
    16'b00010101_01011011 : OUT <= 0;  //21 / 91 = 0
    16'b00010101_01011100 : OUT <= 0;  //21 / 92 = 0
    16'b00010101_01011101 : OUT <= 0;  //21 / 93 = 0
    16'b00010101_01011110 : OUT <= 0;  //21 / 94 = 0
    16'b00010101_01011111 : OUT <= 0;  //21 / 95 = 0
    16'b00010101_01100000 : OUT <= 0;  //21 / 96 = 0
    16'b00010101_01100001 : OUT <= 0;  //21 / 97 = 0
    16'b00010101_01100010 : OUT <= 0;  //21 / 98 = 0
    16'b00010101_01100011 : OUT <= 0;  //21 / 99 = 0
    16'b00010101_01100100 : OUT <= 0;  //21 / 100 = 0
    16'b00010101_01100101 : OUT <= 0;  //21 / 101 = 0
    16'b00010101_01100110 : OUT <= 0;  //21 / 102 = 0
    16'b00010101_01100111 : OUT <= 0;  //21 / 103 = 0
    16'b00010101_01101000 : OUT <= 0;  //21 / 104 = 0
    16'b00010101_01101001 : OUT <= 0;  //21 / 105 = 0
    16'b00010101_01101010 : OUT <= 0;  //21 / 106 = 0
    16'b00010101_01101011 : OUT <= 0;  //21 / 107 = 0
    16'b00010101_01101100 : OUT <= 0;  //21 / 108 = 0
    16'b00010101_01101101 : OUT <= 0;  //21 / 109 = 0
    16'b00010101_01101110 : OUT <= 0;  //21 / 110 = 0
    16'b00010101_01101111 : OUT <= 0;  //21 / 111 = 0
    16'b00010101_01110000 : OUT <= 0;  //21 / 112 = 0
    16'b00010101_01110001 : OUT <= 0;  //21 / 113 = 0
    16'b00010101_01110010 : OUT <= 0;  //21 / 114 = 0
    16'b00010101_01110011 : OUT <= 0;  //21 / 115 = 0
    16'b00010101_01110100 : OUT <= 0;  //21 / 116 = 0
    16'b00010101_01110101 : OUT <= 0;  //21 / 117 = 0
    16'b00010101_01110110 : OUT <= 0;  //21 / 118 = 0
    16'b00010101_01110111 : OUT <= 0;  //21 / 119 = 0
    16'b00010101_01111000 : OUT <= 0;  //21 / 120 = 0
    16'b00010101_01111001 : OUT <= 0;  //21 / 121 = 0
    16'b00010101_01111010 : OUT <= 0;  //21 / 122 = 0
    16'b00010101_01111011 : OUT <= 0;  //21 / 123 = 0
    16'b00010101_01111100 : OUT <= 0;  //21 / 124 = 0
    16'b00010101_01111101 : OUT <= 0;  //21 / 125 = 0
    16'b00010101_01111110 : OUT <= 0;  //21 / 126 = 0
    16'b00010101_01111111 : OUT <= 0;  //21 / 127 = 0
    16'b00010101_10000000 : OUT <= 0;  //21 / 128 = 0
    16'b00010101_10000001 : OUT <= 0;  //21 / 129 = 0
    16'b00010101_10000010 : OUT <= 0;  //21 / 130 = 0
    16'b00010101_10000011 : OUT <= 0;  //21 / 131 = 0
    16'b00010101_10000100 : OUT <= 0;  //21 / 132 = 0
    16'b00010101_10000101 : OUT <= 0;  //21 / 133 = 0
    16'b00010101_10000110 : OUT <= 0;  //21 / 134 = 0
    16'b00010101_10000111 : OUT <= 0;  //21 / 135 = 0
    16'b00010101_10001000 : OUT <= 0;  //21 / 136 = 0
    16'b00010101_10001001 : OUT <= 0;  //21 / 137 = 0
    16'b00010101_10001010 : OUT <= 0;  //21 / 138 = 0
    16'b00010101_10001011 : OUT <= 0;  //21 / 139 = 0
    16'b00010101_10001100 : OUT <= 0;  //21 / 140 = 0
    16'b00010101_10001101 : OUT <= 0;  //21 / 141 = 0
    16'b00010101_10001110 : OUT <= 0;  //21 / 142 = 0
    16'b00010101_10001111 : OUT <= 0;  //21 / 143 = 0
    16'b00010101_10010000 : OUT <= 0;  //21 / 144 = 0
    16'b00010101_10010001 : OUT <= 0;  //21 / 145 = 0
    16'b00010101_10010010 : OUT <= 0;  //21 / 146 = 0
    16'b00010101_10010011 : OUT <= 0;  //21 / 147 = 0
    16'b00010101_10010100 : OUT <= 0;  //21 / 148 = 0
    16'b00010101_10010101 : OUT <= 0;  //21 / 149 = 0
    16'b00010101_10010110 : OUT <= 0;  //21 / 150 = 0
    16'b00010101_10010111 : OUT <= 0;  //21 / 151 = 0
    16'b00010101_10011000 : OUT <= 0;  //21 / 152 = 0
    16'b00010101_10011001 : OUT <= 0;  //21 / 153 = 0
    16'b00010101_10011010 : OUT <= 0;  //21 / 154 = 0
    16'b00010101_10011011 : OUT <= 0;  //21 / 155 = 0
    16'b00010101_10011100 : OUT <= 0;  //21 / 156 = 0
    16'b00010101_10011101 : OUT <= 0;  //21 / 157 = 0
    16'b00010101_10011110 : OUT <= 0;  //21 / 158 = 0
    16'b00010101_10011111 : OUT <= 0;  //21 / 159 = 0
    16'b00010101_10100000 : OUT <= 0;  //21 / 160 = 0
    16'b00010101_10100001 : OUT <= 0;  //21 / 161 = 0
    16'b00010101_10100010 : OUT <= 0;  //21 / 162 = 0
    16'b00010101_10100011 : OUT <= 0;  //21 / 163 = 0
    16'b00010101_10100100 : OUT <= 0;  //21 / 164 = 0
    16'b00010101_10100101 : OUT <= 0;  //21 / 165 = 0
    16'b00010101_10100110 : OUT <= 0;  //21 / 166 = 0
    16'b00010101_10100111 : OUT <= 0;  //21 / 167 = 0
    16'b00010101_10101000 : OUT <= 0;  //21 / 168 = 0
    16'b00010101_10101001 : OUT <= 0;  //21 / 169 = 0
    16'b00010101_10101010 : OUT <= 0;  //21 / 170 = 0
    16'b00010101_10101011 : OUT <= 0;  //21 / 171 = 0
    16'b00010101_10101100 : OUT <= 0;  //21 / 172 = 0
    16'b00010101_10101101 : OUT <= 0;  //21 / 173 = 0
    16'b00010101_10101110 : OUT <= 0;  //21 / 174 = 0
    16'b00010101_10101111 : OUT <= 0;  //21 / 175 = 0
    16'b00010101_10110000 : OUT <= 0;  //21 / 176 = 0
    16'b00010101_10110001 : OUT <= 0;  //21 / 177 = 0
    16'b00010101_10110010 : OUT <= 0;  //21 / 178 = 0
    16'b00010101_10110011 : OUT <= 0;  //21 / 179 = 0
    16'b00010101_10110100 : OUT <= 0;  //21 / 180 = 0
    16'b00010101_10110101 : OUT <= 0;  //21 / 181 = 0
    16'b00010101_10110110 : OUT <= 0;  //21 / 182 = 0
    16'b00010101_10110111 : OUT <= 0;  //21 / 183 = 0
    16'b00010101_10111000 : OUT <= 0;  //21 / 184 = 0
    16'b00010101_10111001 : OUT <= 0;  //21 / 185 = 0
    16'b00010101_10111010 : OUT <= 0;  //21 / 186 = 0
    16'b00010101_10111011 : OUT <= 0;  //21 / 187 = 0
    16'b00010101_10111100 : OUT <= 0;  //21 / 188 = 0
    16'b00010101_10111101 : OUT <= 0;  //21 / 189 = 0
    16'b00010101_10111110 : OUT <= 0;  //21 / 190 = 0
    16'b00010101_10111111 : OUT <= 0;  //21 / 191 = 0
    16'b00010101_11000000 : OUT <= 0;  //21 / 192 = 0
    16'b00010101_11000001 : OUT <= 0;  //21 / 193 = 0
    16'b00010101_11000010 : OUT <= 0;  //21 / 194 = 0
    16'b00010101_11000011 : OUT <= 0;  //21 / 195 = 0
    16'b00010101_11000100 : OUT <= 0;  //21 / 196 = 0
    16'b00010101_11000101 : OUT <= 0;  //21 / 197 = 0
    16'b00010101_11000110 : OUT <= 0;  //21 / 198 = 0
    16'b00010101_11000111 : OUT <= 0;  //21 / 199 = 0
    16'b00010101_11001000 : OUT <= 0;  //21 / 200 = 0
    16'b00010101_11001001 : OUT <= 0;  //21 / 201 = 0
    16'b00010101_11001010 : OUT <= 0;  //21 / 202 = 0
    16'b00010101_11001011 : OUT <= 0;  //21 / 203 = 0
    16'b00010101_11001100 : OUT <= 0;  //21 / 204 = 0
    16'b00010101_11001101 : OUT <= 0;  //21 / 205 = 0
    16'b00010101_11001110 : OUT <= 0;  //21 / 206 = 0
    16'b00010101_11001111 : OUT <= 0;  //21 / 207 = 0
    16'b00010101_11010000 : OUT <= 0;  //21 / 208 = 0
    16'b00010101_11010001 : OUT <= 0;  //21 / 209 = 0
    16'b00010101_11010010 : OUT <= 0;  //21 / 210 = 0
    16'b00010101_11010011 : OUT <= 0;  //21 / 211 = 0
    16'b00010101_11010100 : OUT <= 0;  //21 / 212 = 0
    16'b00010101_11010101 : OUT <= 0;  //21 / 213 = 0
    16'b00010101_11010110 : OUT <= 0;  //21 / 214 = 0
    16'b00010101_11010111 : OUT <= 0;  //21 / 215 = 0
    16'b00010101_11011000 : OUT <= 0;  //21 / 216 = 0
    16'b00010101_11011001 : OUT <= 0;  //21 / 217 = 0
    16'b00010101_11011010 : OUT <= 0;  //21 / 218 = 0
    16'b00010101_11011011 : OUT <= 0;  //21 / 219 = 0
    16'b00010101_11011100 : OUT <= 0;  //21 / 220 = 0
    16'b00010101_11011101 : OUT <= 0;  //21 / 221 = 0
    16'b00010101_11011110 : OUT <= 0;  //21 / 222 = 0
    16'b00010101_11011111 : OUT <= 0;  //21 / 223 = 0
    16'b00010101_11100000 : OUT <= 0;  //21 / 224 = 0
    16'b00010101_11100001 : OUT <= 0;  //21 / 225 = 0
    16'b00010101_11100010 : OUT <= 0;  //21 / 226 = 0
    16'b00010101_11100011 : OUT <= 0;  //21 / 227 = 0
    16'b00010101_11100100 : OUT <= 0;  //21 / 228 = 0
    16'b00010101_11100101 : OUT <= 0;  //21 / 229 = 0
    16'b00010101_11100110 : OUT <= 0;  //21 / 230 = 0
    16'b00010101_11100111 : OUT <= 0;  //21 / 231 = 0
    16'b00010101_11101000 : OUT <= 0;  //21 / 232 = 0
    16'b00010101_11101001 : OUT <= 0;  //21 / 233 = 0
    16'b00010101_11101010 : OUT <= 0;  //21 / 234 = 0
    16'b00010101_11101011 : OUT <= 0;  //21 / 235 = 0
    16'b00010101_11101100 : OUT <= 0;  //21 / 236 = 0
    16'b00010101_11101101 : OUT <= 0;  //21 / 237 = 0
    16'b00010101_11101110 : OUT <= 0;  //21 / 238 = 0
    16'b00010101_11101111 : OUT <= 0;  //21 / 239 = 0
    16'b00010101_11110000 : OUT <= 0;  //21 / 240 = 0
    16'b00010101_11110001 : OUT <= 0;  //21 / 241 = 0
    16'b00010101_11110010 : OUT <= 0;  //21 / 242 = 0
    16'b00010101_11110011 : OUT <= 0;  //21 / 243 = 0
    16'b00010101_11110100 : OUT <= 0;  //21 / 244 = 0
    16'b00010101_11110101 : OUT <= 0;  //21 / 245 = 0
    16'b00010101_11110110 : OUT <= 0;  //21 / 246 = 0
    16'b00010101_11110111 : OUT <= 0;  //21 / 247 = 0
    16'b00010101_11111000 : OUT <= 0;  //21 / 248 = 0
    16'b00010101_11111001 : OUT <= 0;  //21 / 249 = 0
    16'b00010101_11111010 : OUT <= 0;  //21 / 250 = 0
    16'b00010101_11111011 : OUT <= 0;  //21 / 251 = 0
    16'b00010101_11111100 : OUT <= 0;  //21 / 252 = 0
    16'b00010101_11111101 : OUT <= 0;  //21 / 253 = 0
    16'b00010101_11111110 : OUT <= 0;  //21 / 254 = 0
    16'b00010101_11111111 : OUT <= 0;  //21 / 255 = 0
    16'b00010110_00000000 : OUT <= 0;  //22 / 0 = 0
    16'b00010110_00000001 : OUT <= 22;  //22 / 1 = 22
    16'b00010110_00000010 : OUT <= 11;  //22 / 2 = 11
    16'b00010110_00000011 : OUT <= 7;  //22 / 3 = 7
    16'b00010110_00000100 : OUT <= 5;  //22 / 4 = 5
    16'b00010110_00000101 : OUT <= 4;  //22 / 5 = 4
    16'b00010110_00000110 : OUT <= 3;  //22 / 6 = 3
    16'b00010110_00000111 : OUT <= 3;  //22 / 7 = 3
    16'b00010110_00001000 : OUT <= 2;  //22 / 8 = 2
    16'b00010110_00001001 : OUT <= 2;  //22 / 9 = 2
    16'b00010110_00001010 : OUT <= 2;  //22 / 10 = 2
    16'b00010110_00001011 : OUT <= 2;  //22 / 11 = 2
    16'b00010110_00001100 : OUT <= 1;  //22 / 12 = 1
    16'b00010110_00001101 : OUT <= 1;  //22 / 13 = 1
    16'b00010110_00001110 : OUT <= 1;  //22 / 14 = 1
    16'b00010110_00001111 : OUT <= 1;  //22 / 15 = 1
    16'b00010110_00010000 : OUT <= 1;  //22 / 16 = 1
    16'b00010110_00010001 : OUT <= 1;  //22 / 17 = 1
    16'b00010110_00010010 : OUT <= 1;  //22 / 18 = 1
    16'b00010110_00010011 : OUT <= 1;  //22 / 19 = 1
    16'b00010110_00010100 : OUT <= 1;  //22 / 20 = 1
    16'b00010110_00010101 : OUT <= 1;  //22 / 21 = 1
    16'b00010110_00010110 : OUT <= 1;  //22 / 22 = 1
    16'b00010110_00010111 : OUT <= 0;  //22 / 23 = 0
    16'b00010110_00011000 : OUT <= 0;  //22 / 24 = 0
    16'b00010110_00011001 : OUT <= 0;  //22 / 25 = 0
    16'b00010110_00011010 : OUT <= 0;  //22 / 26 = 0
    16'b00010110_00011011 : OUT <= 0;  //22 / 27 = 0
    16'b00010110_00011100 : OUT <= 0;  //22 / 28 = 0
    16'b00010110_00011101 : OUT <= 0;  //22 / 29 = 0
    16'b00010110_00011110 : OUT <= 0;  //22 / 30 = 0
    16'b00010110_00011111 : OUT <= 0;  //22 / 31 = 0
    16'b00010110_00100000 : OUT <= 0;  //22 / 32 = 0
    16'b00010110_00100001 : OUT <= 0;  //22 / 33 = 0
    16'b00010110_00100010 : OUT <= 0;  //22 / 34 = 0
    16'b00010110_00100011 : OUT <= 0;  //22 / 35 = 0
    16'b00010110_00100100 : OUT <= 0;  //22 / 36 = 0
    16'b00010110_00100101 : OUT <= 0;  //22 / 37 = 0
    16'b00010110_00100110 : OUT <= 0;  //22 / 38 = 0
    16'b00010110_00100111 : OUT <= 0;  //22 / 39 = 0
    16'b00010110_00101000 : OUT <= 0;  //22 / 40 = 0
    16'b00010110_00101001 : OUT <= 0;  //22 / 41 = 0
    16'b00010110_00101010 : OUT <= 0;  //22 / 42 = 0
    16'b00010110_00101011 : OUT <= 0;  //22 / 43 = 0
    16'b00010110_00101100 : OUT <= 0;  //22 / 44 = 0
    16'b00010110_00101101 : OUT <= 0;  //22 / 45 = 0
    16'b00010110_00101110 : OUT <= 0;  //22 / 46 = 0
    16'b00010110_00101111 : OUT <= 0;  //22 / 47 = 0
    16'b00010110_00110000 : OUT <= 0;  //22 / 48 = 0
    16'b00010110_00110001 : OUT <= 0;  //22 / 49 = 0
    16'b00010110_00110010 : OUT <= 0;  //22 / 50 = 0
    16'b00010110_00110011 : OUT <= 0;  //22 / 51 = 0
    16'b00010110_00110100 : OUT <= 0;  //22 / 52 = 0
    16'b00010110_00110101 : OUT <= 0;  //22 / 53 = 0
    16'b00010110_00110110 : OUT <= 0;  //22 / 54 = 0
    16'b00010110_00110111 : OUT <= 0;  //22 / 55 = 0
    16'b00010110_00111000 : OUT <= 0;  //22 / 56 = 0
    16'b00010110_00111001 : OUT <= 0;  //22 / 57 = 0
    16'b00010110_00111010 : OUT <= 0;  //22 / 58 = 0
    16'b00010110_00111011 : OUT <= 0;  //22 / 59 = 0
    16'b00010110_00111100 : OUT <= 0;  //22 / 60 = 0
    16'b00010110_00111101 : OUT <= 0;  //22 / 61 = 0
    16'b00010110_00111110 : OUT <= 0;  //22 / 62 = 0
    16'b00010110_00111111 : OUT <= 0;  //22 / 63 = 0
    16'b00010110_01000000 : OUT <= 0;  //22 / 64 = 0
    16'b00010110_01000001 : OUT <= 0;  //22 / 65 = 0
    16'b00010110_01000010 : OUT <= 0;  //22 / 66 = 0
    16'b00010110_01000011 : OUT <= 0;  //22 / 67 = 0
    16'b00010110_01000100 : OUT <= 0;  //22 / 68 = 0
    16'b00010110_01000101 : OUT <= 0;  //22 / 69 = 0
    16'b00010110_01000110 : OUT <= 0;  //22 / 70 = 0
    16'b00010110_01000111 : OUT <= 0;  //22 / 71 = 0
    16'b00010110_01001000 : OUT <= 0;  //22 / 72 = 0
    16'b00010110_01001001 : OUT <= 0;  //22 / 73 = 0
    16'b00010110_01001010 : OUT <= 0;  //22 / 74 = 0
    16'b00010110_01001011 : OUT <= 0;  //22 / 75 = 0
    16'b00010110_01001100 : OUT <= 0;  //22 / 76 = 0
    16'b00010110_01001101 : OUT <= 0;  //22 / 77 = 0
    16'b00010110_01001110 : OUT <= 0;  //22 / 78 = 0
    16'b00010110_01001111 : OUT <= 0;  //22 / 79 = 0
    16'b00010110_01010000 : OUT <= 0;  //22 / 80 = 0
    16'b00010110_01010001 : OUT <= 0;  //22 / 81 = 0
    16'b00010110_01010010 : OUT <= 0;  //22 / 82 = 0
    16'b00010110_01010011 : OUT <= 0;  //22 / 83 = 0
    16'b00010110_01010100 : OUT <= 0;  //22 / 84 = 0
    16'b00010110_01010101 : OUT <= 0;  //22 / 85 = 0
    16'b00010110_01010110 : OUT <= 0;  //22 / 86 = 0
    16'b00010110_01010111 : OUT <= 0;  //22 / 87 = 0
    16'b00010110_01011000 : OUT <= 0;  //22 / 88 = 0
    16'b00010110_01011001 : OUT <= 0;  //22 / 89 = 0
    16'b00010110_01011010 : OUT <= 0;  //22 / 90 = 0
    16'b00010110_01011011 : OUT <= 0;  //22 / 91 = 0
    16'b00010110_01011100 : OUT <= 0;  //22 / 92 = 0
    16'b00010110_01011101 : OUT <= 0;  //22 / 93 = 0
    16'b00010110_01011110 : OUT <= 0;  //22 / 94 = 0
    16'b00010110_01011111 : OUT <= 0;  //22 / 95 = 0
    16'b00010110_01100000 : OUT <= 0;  //22 / 96 = 0
    16'b00010110_01100001 : OUT <= 0;  //22 / 97 = 0
    16'b00010110_01100010 : OUT <= 0;  //22 / 98 = 0
    16'b00010110_01100011 : OUT <= 0;  //22 / 99 = 0
    16'b00010110_01100100 : OUT <= 0;  //22 / 100 = 0
    16'b00010110_01100101 : OUT <= 0;  //22 / 101 = 0
    16'b00010110_01100110 : OUT <= 0;  //22 / 102 = 0
    16'b00010110_01100111 : OUT <= 0;  //22 / 103 = 0
    16'b00010110_01101000 : OUT <= 0;  //22 / 104 = 0
    16'b00010110_01101001 : OUT <= 0;  //22 / 105 = 0
    16'b00010110_01101010 : OUT <= 0;  //22 / 106 = 0
    16'b00010110_01101011 : OUT <= 0;  //22 / 107 = 0
    16'b00010110_01101100 : OUT <= 0;  //22 / 108 = 0
    16'b00010110_01101101 : OUT <= 0;  //22 / 109 = 0
    16'b00010110_01101110 : OUT <= 0;  //22 / 110 = 0
    16'b00010110_01101111 : OUT <= 0;  //22 / 111 = 0
    16'b00010110_01110000 : OUT <= 0;  //22 / 112 = 0
    16'b00010110_01110001 : OUT <= 0;  //22 / 113 = 0
    16'b00010110_01110010 : OUT <= 0;  //22 / 114 = 0
    16'b00010110_01110011 : OUT <= 0;  //22 / 115 = 0
    16'b00010110_01110100 : OUT <= 0;  //22 / 116 = 0
    16'b00010110_01110101 : OUT <= 0;  //22 / 117 = 0
    16'b00010110_01110110 : OUT <= 0;  //22 / 118 = 0
    16'b00010110_01110111 : OUT <= 0;  //22 / 119 = 0
    16'b00010110_01111000 : OUT <= 0;  //22 / 120 = 0
    16'b00010110_01111001 : OUT <= 0;  //22 / 121 = 0
    16'b00010110_01111010 : OUT <= 0;  //22 / 122 = 0
    16'b00010110_01111011 : OUT <= 0;  //22 / 123 = 0
    16'b00010110_01111100 : OUT <= 0;  //22 / 124 = 0
    16'b00010110_01111101 : OUT <= 0;  //22 / 125 = 0
    16'b00010110_01111110 : OUT <= 0;  //22 / 126 = 0
    16'b00010110_01111111 : OUT <= 0;  //22 / 127 = 0
    16'b00010110_10000000 : OUT <= 0;  //22 / 128 = 0
    16'b00010110_10000001 : OUT <= 0;  //22 / 129 = 0
    16'b00010110_10000010 : OUT <= 0;  //22 / 130 = 0
    16'b00010110_10000011 : OUT <= 0;  //22 / 131 = 0
    16'b00010110_10000100 : OUT <= 0;  //22 / 132 = 0
    16'b00010110_10000101 : OUT <= 0;  //22 / 133 = 0
    16'b00010110_10000110 : OUT <= 0;  //22 / 134 = 0
    16'b00010110_10000111 : OUT <= 0;  //22 / 135 = 0
    16'b00010110_10001000 : OUT <= 0;  //22 / 136 = 0
    16'b00010110_10001001 : OUT <= 0;  //22 / 137 = 0
    16'b00010110_10001010 : OUT <= 0;  //22 / 138 = 0
    16'b00010110_10001011 : OUT <= 0;  //22 / 139 = 0
    16'b00010110_10001100 : OUT <= 0;  //22 / 140 = 0
    16'b00010110_10001101 : OUT <= 0;  //22 / 141 = 0
    16'b00010110_10001110 : OUT <= 0;  //22 / 142 = 0
    16'b00010110_10001111 : OUT <= 0;  //22 / 143 = 0
    16'b00010110_10010000 : OUT <= 0;  //22 / 144 = 0
    16'b00010110_10010001 : OUT <= 0;  //22 / 145 = 0
    16'b00010110_10010010 : OUT <= 0;  //22 / 146 = 0
    16'b00010110_10010011 : OUT <= 0;  //22 / 147 = 0
    16'b00010110_10010100 : OUT <= 0;  //22 / 148 = 0
    16'b00010110_10010101 : OUT <= 0;  //22 / 149 = 0
    16'b00010110_10010110 : OUT <= 0;  //22 / 150 = 0
    16'b00010110_10010111 : OUT <= 0;  //22 / 151 = 0
    16'b00010110_10011000 : OUT <= 0;  //22 / 152 = 0
    16'b00010110_10011001 : OUT <= 0;  //22 / 153 = 0
    16'b00010110_10011010 : OUT <= 0;  //22 / 154 = 0
    16'b00010110_10011011 : OUT <= 0;  //22 / 155 = 0
    16'b00010110_10011100 : OUT <= 0;  //22 / 156 = 0
    16'b00010110_10011101 : OUT <= 0;  //22 / 157 = 0
    16'b00010110_10011110 : OUT <= 0;  //22 / 158 = 0
    16'b00010110_10011111 : OUT <= 0;  //22 / 159 = 0
    16'b00010110_10100000 : OUT <= 0;  //22 / 160 = 0
    16'b00010110_10100001 : OUT <= 0;  //22 / 161 = 0
    16'b00010110_10100010 : OUT <= 0;  //22 / 162 = 0
    16'b00010110_10100011 : OUT <= 0;  //22 / 163 = 0
    16'b00010110_10100100 : OUT <= 0;  //22 / 164 = 0
    16'b00010110_10100101 : OUT <= 0;  //22 / 165 = 0
    16'b00010110_10100110 : OUT <= 0;  //22 / 166 = 0
    16'b00010110_10100111 : OUT <= 0;  //22 / 167 = 0
    16'b00010110_10101000 : OUT <= 0;  //22 / 168 = 0
    16'b00010110_10101001 : OUT <= 0;  //22 / 169 = 0
    16'b00010110_10101010 : OUT <= 0;  //22 / 170 = 0
    16'b00010110_10101011 : OUT <= 0;  //22 / 171 = 0
    16'b00010110_10101100 : OUT <= 0;  //22 / 172 = 0
    16'b00010110_10101101 : OUT <= 0;  //22 / 173 = 0
    16'b00010110_10101110 : OUT <= 0;  //22 / 174 = 0
    16'b00010110_10101111 : OUT <= 0;  //22 / 175 = 0
    16'b00010110_10110000 : OUT <= 0;  //22 / 176 = 0
    16'b00010110_10110001 : OUT <= 0;  //22 / 177 = 0
    16'b00010110_10110010 : OUT <= 0;  //22 / 178 = 0
    16'b00010110_10110011 : OUT <= 0;  //22 / 179 = 0
    16'b00010110_10110100 : OUT <= 0;  //22 / 180 = 0
    16'b00010110_10110101 : OUT <= 0;  //22 / 181 = 0
    16'b00010110_10110110 : OUT <= 0;  //22 / 182 = 0
    16'b00010110_10110111 : OUT <= 0;  //22 / 183 = 0
    16'b00010110_10111000 : OUT <= 0;  //22 / 184 = 0
    16'b00010110_10111001 : OUT <= 0;  //22 / 185 = 0
    16'b00010110_10111010 : OUT <= 0;  //22 / 186 = 0
    16'b00010110_10111011 : OUT <= 0;  //22 / 187 = 0
    16'b00010110_10111100 : OUT <= 0;  //22 / 188 = 0
    16'b00010110_10111101 : OUT <= 0;  //22 / 189 = 0
    16'b00010110_10111110 : OUT <= 0;  //22 / 190 = 0
    16'b00010110_10111111 : OUT <= 0;  //22 / 191 = 0
    16'b00010110_11000000 : OUT <= 0;  //22 / 192 = 0
    16'b00010110_11000001 : OUT <= 0;  //22 / 193 = 0
    16'b00010110_11000010 : OUT <= 0;  //22 / 194 = 0
    16'b00010110_11000011 : OUT <= 0;  //22 / 195 = 0
    16'b00010110_11000100 : OUT <= 0;  //22 / 196 = 0
    16'b00010110_11000101 : OUT <= 0;  //22 / 197 = 0
    16'b00010110_11000110 : OUT <= 0;  //22 / 198 = 0
    16'b00010110_11000111 : OUT <= 0;  //22 / 199 = 0
    16'b00010110_11001000 : OUT <= 0;  //22 / 200 = 0
    16'b00010110_11001001 : OUT <= 0;  //22 / 201 = 0
    16'b00010110_11001010 : OUT <= 0;  //22 / 202 = 0
    16'b00010110_11001011 : OUT <= 0;  //22 / 203 = 0
    16'b00010110_11001100 : OUT <= 0;  //22 / 204 = 0
    16'b00010110_11001101 : OUT <= 0;  //22 / 205 = 0
    16'b00010110_11001110 : OUT <= 0;  //22 / 206 = 0
    16'b00010110_11001111 : OUT <= 0;  //22 / 207 = 0
    16'b00010110_11010000 : OUT <= 0;  //22 / 208 = 0
    16'b00010110_11010001 : OUT <= 0;  //22 / 209 = 0
    16'b00010110_11010010 : OUT <= 0;  //22 / 210 = 0
    16'b00010110_11010011 : OUT <= 0;  //22 / 211 = 0
    16'b00010110_11010100 : OUT <= 0;  //22 / 212 = 0
    16'b00010110_11010101 : OUT <= 0;  //22 / 213 = 0
    16'b00010110_11010110 : OUT <= 0;  //22 / 214 = 0
    16'b00010110_11010111 : OUT <= 0;  //22 / 215 = 0
    16'b00010110_11011000 : OUT <= 0;  //22 / 216 = 0
    16'b00010110_11011001 : OUT <= 0;  //22 / 217 = 0
    16'b00010110_11011010 : OUT <= 0;  //22 / 218 = 0
    16'b00010110_11011011 : OUT <= 0;  //22 / 219 = 0
    16'b00010110_11011100 : OUT <= 0;  //22 / 220 = 0
    16'b00010110_11011101 : OUT <= 0;  //22 / 221 = 0
    16'b00010110_11011110 : OUT <= 0;  //22 / 222 = 0
    16'b00010110_11011111 : OUT <= 0;  //22 / 223 = 0
    16'b00010110_11100000 : OUT <= 0;  //22 / 224 = 0
    16'b00010110_11100001 : OUT <= 0;  //22 / 225 = 0
    16'b00010110_11100010 : OUT <= 0;  //22 / 226 = 0
    16'b00010110_11100011 : OUT <= 0;  //22 / 227 = 0
    16'b00010110_11100100 : OUT <= 0;  //22 / 228 = 0
    16'b00010110_11100101 : OUT <= 0;  //22 / 229 = 0
    16'b00010110_11100110 : OUT <= 0;  //22 / 230 = 0
    16'b00010110_11100111 : OUT <= 0;  //22 / 231 = 0
    16'b00010110_11101000 : OUT <= 0;  //22 / 232 = 0
    16'b00010110_11101001 : OUT <= 0;  //22 / 233 = 0
    16'b00010110_11101010 : OUT <= 0;  //22 / 234 = 0
    16'b00010110_11101011 : OUT <= 0;  //22 / 235 = 0
    16'b00010110_11101100 : OUT <= 0;  //22 / 236 = 0
    16'b00010110_11101101 : OUT <= 0;  //22 / 237 = 0
    16'b00010110_11101110 : OUT <= 0;  //22 / 238 = 0
    16'b00010110_11101111 : OUT <= 0;  //22 / 239 = 0
    16'b00010110_11110000 : OUT <= 0;  //22 / 240 = 0
    16'b00010110_11110001 : OUT <= 0;  //22 / 241 = 0
    16'b00010110_11110010 : OUT <= 0;  //22 / 242 = 0
    16'b00010110_11110011 : OUT <= 0;  //22 / 243 = 0
    16'b00010110_11110100 : OUT <= 0;  //22 / 244 = 0
    16'b00010110_11110101 : OUT <= 0;  //22 / 245 = 0
    16'b00010110_11110110 : OUT <= 0;  //22 / 246 = 0
    16'b00010110_11110111 : OUT <= 0;  //22 / 247 = 0
    16'b00010110_11111000 : OUT <= 0;  //22 / 248 = 0
    16'b00010110_11111001 : OUT <= 0;  //22 / 249 = 0
    16'b00010110_11111010 : OUT <= 0;  //22 / 250 = 0
    16'b00010110_11111011 : OUT <= 0;  //22 / 251 = 0
    16'b00010110_11111100 : OUT <= 0;  //22 / 252 = 0
    16'b00010110_11111101 : OUT <= 0;  //22 / 253 = 0
    16'b00010110_11111110 : OUT <= 0;  //22 / 254 = 0
    16'b00010110_11111111 : OUT <= 0;  //22 / 255 = 0
    16'b00010111_00000000 : OUT <= 0;  //23 / 0 = 0
    16'b00010111_00000001 : OUT <= 23;  //23 / 1 = 23
    16'b00010111_00000010 : OUT <= 11;  //23 / 2 = 11
    16'b00010111_00000011 : OUT <= 7;  //23 / 3 = 7
    16'b00010111_00000100 : OUT <= 5;  //23 / 4 = 5
    16'b00010111_00000101 : OUT <= 4;  //23 / 5 = 4
    16'b00010111_00000110 : OUT <= 3;  //23 / 6 = 3
    16'b00010111_00000111 : OUT <= 3;  //23 / 7 = 3
    16'b00010111_00001000 : OUT <= 2;  //23 / 8 = 2
    16'b00010111_00001001 : OUT <= 2;  //23 / 9 = 2
    16'b00010111_00001010 : OUT <= 2;  //23 / 10 = 2
    16'b00010111_00001011 : OUT <= 2;  //23 / 11 = 2
    16'b00010111_00001100 : OUT <= 1;  //23 / 12 = 1
    16'b00010111_00001101 : OUT <= 1;  //23 / 13 = 1
    16'b00010111_00001110 : OUT <= 1;  //23 / 14 = 1
    16'b00010111_00001111 : OUT <= 1;  //23 / 15 = 1
    16'b00010111_00010000 : OUT <= 1;  //23 / 16 = 1
    16'b00010111_00010001 : OUT <= 1;  //23 / 17 = 1
    16'b00010111_00010010 : OUT <= 1;  //23 / 18 = 1
    16'b00010111_00010011 : OUT <= 1;  //23 / 19 = 1
    16'b00010111_00010100 : OUT <= 1;  //23 / 20 = 1
    16'b00010111_00010101 : OUT <= 1;  //23 / 21 = 1
    16'b00010111_00010110 : OUT <= 1;  //23 / 22 = 1
    16'b00010111_00010111 : OUT <= 1;  //23 / 23 = 1
    16'b00010111_00011000 : OUT <= 0;  //23 / 24 = 0
    16'b00010111_00011001 : OUT <= 0;  //23 / 25 = 0
    16'b00010111_00011010 : OUT <= 0;  //23 / 26 = 0
    16'b00010111_00011011 : OUT <= 0;  //23 / 27 = 0
    16'b00010111_00011100 : OUT <= 0;  //23 / 28 = 0
    16'b00010111_00011101 : OUT <= 0;  //23 / 29 = 0
    16'b00010111_00011110 : OUT <= 0;  //23 / 30 = 0
    16'b00010111_00011111 : OUT <= 0;  //23 / 31 = 0
    16'b00010111_00100000 : OUT <= 0;  //23 / 32 = 0
    16'b00010111_00100001 : OUT <= 0;  //23 / 33 = 0
    16'b00010111_00100010 : OUT <= 0;  //23 / 34 = 0
    16'b00010111_00100011 : OUT <= 0;  //23 / 35 = 0
    16'b00010111_00100100 : OUT <= 0;  //23 / 36 = 0
    16'b00010111_00100101 : OUT <= 0;  //23 / 37 = 0
    16'b00010111_00100110 : OUT <= 0;  //23 / 38 = 0
    16'b00010111_00100111 : OUT <= 0;  //23 / 39 = 0
    16'b00010111_00101000 : OUT <= 0;  //23 / 40 = 0
    16'b00010111_00101001 : OUT <= 0;  //23 / 41 = 0
    16'b00010111_00101010 : OUT <= 0;  //23 / 42 = 0
    16'b00010111_00101011 : OUT <= 0;  //23 / 43 = 0
    16'b00010111_00101100 : OUT <= 0;  //23 / 44 = 0
    16'b00010111_00101101 : OUT <= 0;  //23 / 45 = 0
    16'b00010111_00101110 : OUT <= 0;  //23 / 46 = 0
    16'b00010111_00101111 : OUT <= 0;  //23 / 47 = 0
    16'b00010111_00110000 : OUT <= 0;  //23 / 48 = 0
    16'b00010111_00110001 : OUT <= 0;  //23 / 49 = 0
    16'b00010111_00110010 : OUT <= 0;  //23 / 50 = 0
    16'b00010111_00110011 : OUT <= 0;  //23 / 51 = 0
    16'b00010111_00110100 : OUT <= 0;  //23 / 52 = 0
    16'b00010111_00110101 : OUT <= 0;  //23 / 53 = 0
    16'b00010111_00110110 : OUT <= 0;  //23 / 54 = 0
    16'b00010111_00110111 : OUT <= 0;  //23 / 55 = 0
    16'b00010111_00111000 : OUT <= 0;  //23 / 56 = 0
    16'b00010111_00111001 : OUT <= 0;  //23 / 57 = 0
    16'b00010111_00111010 : OUT <= 0;  //23 / 58 = 0
    16'b00010111_00111011 : OUT <= 0;  //23 / 59 = 0
    16'b00010111_00111100 : OUT <= 0;  //23 / 60 = 0
    16'b00010111_00111101 : OUT <= 0;  //23 / 61 = 0
    16'b00010111_00111110 : OUT <= 0;  //23 / 62 = 0
    16'b00010111_00111111 : OUT <= 0;  //23 / 63 = 0
    16'b00010111_01000000 : OUT <= 0;  //23 / 64 = 0
    16'b00010111_01000001 : OUT <= 0;  //23 / 65 = 0
    16'b00010111_01000010 : OUT <= 0;  //23 / 66 = 0
    16'b00010111_01000011 : OUT <= 0;  //23 / 67 = 0
    16'b00010111_01000100 : OUT <= 0;  //23 / 68 = 0
    16'b00010111_01000101 : OUT <= 0;  //23 / 69 = 0
    16'b00010111_01000110 : OUT <= 0;  //23 / 70 = 0
    16'b00010111_01000111 : OUT <= 0;  //23 / 71 = 0
    16'b00010111_01001000 : OUT <= 0;  //23 / 72 = 0
    16'b00010111_01001001 : OUT <= 0;  //23 / 73 = 0
    16'b00010111_01001010 : OUT <= 0;  //23 / 74 = 0
    16'b00010111_01001011 : OUT <= 0;  //23 / 75 = 0
    16'b00010111_01001100 : OUT <= 0;  //23 / 76 = 0
    16'b00010111_01001101 : OUT <= 0;  //23 / 77 = 0
    16'b00010111_01001110 : OUT <= 0;  //23 / 78 = 0
    16'b00010111_01001111 : OUT <= 0;  //23 / 79 = 0
    16'b00010111_01010000 : OUT <= 0;  //23 / 80 = 0
    16'b00010111_01010001 : OUT <= 0;  //23 / 81 = 0
    16'b00010111_01010010 : OUT <= 0;  //23 / 82 = 0
    16'b00010111_01010011 : OUT <= 0;  //23 / 83 = 0
    16'b00010111_01010100 : OUT <= 0;  //23 / 84 = 0
    16'b00010111_01010101 : OUT <= 0;  //23 / 85 = 0
    16'b00010111_01010110 : OUT <= 0;  //23 / 86 = 0
    16'b00010111_01010111 : OUT <= 0;  //23 / 87 = 0
    16'b00010111_01011000 : OUT <= 0;  //23 / 88 = 0
    16'b00010111_01011001 : OUT <= 0;  //23 / 89 = 0
    16'b00010111_01011010 : OUT <= 0;  //23 / 90 = 0
    16'b00010111_01011011 : OUT <= 0;  //23 / 91 = 0
    16'b00010111_01011100 : OUT <= 0;  //23 / 92 = 0
    16'b00010111_01011101 : OUT <= 0;  //23 / 93 = 0
    16'b00010111_01011110 : OUT <= 0;  //23 / 94 = 0
    16'b00010111_01011111 : OUT <= 0;  //23 / 95 = 0
    16'b00010111_01100000 : OUT <= 0;  //23 / 96 = 0
    16'b00010111_01100001 : OUT <= 0;  //23 / 97 = 0
    16'b00010111_01100010 : OUT <= 0;  //23 / 98 = 0
    16'b00010111_01100011 : OUT <= 0;  //23 / 99 = 0
    16'b00010111_01100100 : OUT <= 0;  //23 / 100 = 0
    16'b00010111_01100101 : OUT <= 0;  //23 / 101 = 0
    16'b00010111_01100110 : OUT <= 0;  //23 / 102 = 0
    16'b00010111_01100111 : OUT <= 0;  //23 / 103 = 0
    16'b00010111_01101000 : OUT <= 0;  //23 / 104 = 0
    16'b00010111_01101001 : OUT <= 0;  //23 / 105 = 0
    16'b00010111_01101010 : OUT <= 0;  //23 / 106 = 0
    16'b00010111_01101011 : OUT <= 0;  //23 / 107 = 0
    16'b00010111_01101100 : OUT <= 0;  //23 / 108 = 0
    16'b00010111_01101101 : OUT <= 0;  //23 / 109 = 0
    16'b00010111_01101110 : OUT <= 0;  //23 / 110 = 0
    16'b00010111_01101111 : OUT <= 0;  //23 / 111 = 0
    16'b00010111_01110000 : OUT <= 0;  //23 / 112 = 0
    16'b00010111_01110001 : OUT <= 0;  //23 / 113 = 0
    16'b00010111_01110010 : OUT <= 0;  //23 / 114 = 0
    16'b00010111_01110011 : OUT <= 0;  //23 / 115 = 0
    16'b00010111_01110100 : OUT <= 0;  //23 / 116 = 0
    16'b00010111_01110101 : OUT <= 0;  //23 / 117 = 0
    16'b00010111_01110110 : OUT <= 0;  //23 / 118 = 0
    16'b00010111_01110111 : OUT <= 0;  //23 / 119 = 0
    16'b00010111_01111000 : OUT <= 0;  //23 / 120 = 0
    16'b00010111_01111001 : OUT <= 0;  //23 / 121 = 0
    16'b00010111_01111010 : OUT <= 0;  //23 / 122 = 0
    16'b00010111_01111011 : OUT <= 0;  //23 / 123 = 0
    16'b00010111_01111100 : OUT <= 0;  //23 / 124 = 0
    16'b00010111_01111101 : OUT <= 0;  //23 / 125 = 0
    16'b00010111_01111110 : OUT <= 0;  //23 / 126 = 0
    16'b00010111_01111111 : OUT <= 0;  //23 / 127 = 0
    16'b00010111_10000000 : OUT <= 0;  //23 / 128 = 0
    16'b00010111_10000001 : OUT <= 0;  //23 / 129 = 0
    16'b00010111_10000010 : OUT <= 0;  //23 / 130 = 0
    16'b00010111_10000011 : OUT <= 0;  //23 / 131 = 0
    16'b00010111_10000100 : OUT <= 0;  //23 / 132 = 0
    16'b00010111_10000101 : OUT <= 0;  //23 / 133 = 0
    16'b00010111_10000110 : OUT <= 0;  //23 / 134 = 0
    16'b00010111_10000111 : OUT <= 0;  //23 / 135 = 0
    16'b00010111_10001000 : OUT <= 0;  //23 / 136 = 0
    16'b00010111_10001001 : OUT <= 0;  //23 / 137 = 0
    16'b00010111_10001010 : OUT <= 0;  //23 / 138 = 0
    16'b00010111_10001011 : OUT <= 0;  //23 / 139 = 0
    16'b00010111_10001100 : OUT <= 0;  //23 / 140 = 0
    16'b00010111_10001101 : OUT <= 0;  //23 / 141 = 0
    16'b00010111_10001110 : OUT <= 0;  //23 / 142 = 0
    16'b00010111_10001111 : OUT <= 0;  //23 / 143 = 0
    16'b00010111_10010000 : OUT <= 0;  //23 / 144 = 0
    16'b00010111_10010001 : OUT <= 0;  //23 / 145 = 0
    16'b00010111_10010010 : OUT <= 0;  //23 / 146 = 0
    16'b00010111_10010011 : OUT <= 0;  //23 / 147 = 0
    16'b00010111_10010100 : OUT <= 0;  //23 / 148 = 0
    16'b00010111_10010101 : OUT <= 0;  //23 / 149 = 0
    16'b00010111_10010110 : OUT <= 0;  //23 / 150 = 0
    16'b00010111_10010111 : OUT <= 0;  //23 / 151 = 0
    16'b00010111_10011000 : OUT <= 0;  //23 / 152 = 0
    16'b00010111_10011001 : OUT <= 0;  //23 / 153 = 0
    16'b00010111_10011010 : OUT <= 0;  //23 / 154 = 0
    16'b00010111_10011011 : OUT <= 0;  //23 / 155 = 0
    16'b00010111_10011100 : OUT <= 0;  //23 / 156 = 0
    16'b00010111_10011101 : OUT <= 0;  //23 / 157 = 0
    16'b00010111_10011110 : OUT <= 0;  //23 / 158 = 0
    16'b00010111_10011111 : OUT <= 0;  //23 / 159 = 0
    16'b00010111_10100000 : OUT <= 0;  //23 / 160 = 0
    16'b00010111_10100001 : OUT <= 0;  //23 / 161 = 0
    16'b00010111_10100010 : OUT <= 0;  //23 / 162 = 0
    16'b00010111_10100011 : OUT <= 0;  //23 / 163 = 0
    16'b00010111_10100100 : OUT <= 0;  //23 / 164 = 0
    16'b00010111_10100101 : OUT <= 0;  //23 / 165 = 0
    16'b00010111_10100110 : OUT <= 0;  //23 / 166 = 0
    16'b00010111_10100111 : OUT <= 0;  //23 / 167 = 0
    16'b00010111_10101000 : OUT <= 0;  //23 / 168 = 0
    16'b00010111_10101001 : OUT <= 0;  //23 / 169 = 0
    16'b00010111_10101010 : OUT <= 0;  //23 / 170 = 0
    16'b00010111_10101011 : OUT <= 0;  //23 / 171 = 0
    16'b00010111_10101100 : OUT <= 0;  //23 / 172 = 0
    16'b00010111_10101101 : OUT <= 0;  //23 / 173 = 0
    16'b00010111_10101110 : OUT <= 0;  //23 / 174 = 0
    16'b00010111_10101111 : OUT <= 0;  //23 / 175 = 0
    16'b00010111_10110000 : OUT <= 0;  //23 / 176 = 0
    16'b00010111_10110001 : OUT <= 0;  //23 / 177 = 0
    16'b00010111_10110010 : OUT <= 0;  //23 / 178 = 0
    16'b00010111_10110011 : OUT <= 0;  //23 / 179 = 0
    16'b00010111_10110100 : OUT <= 0;  //23 / 180 = 0
    16'b00010111_10110101 : OUT <= 0;  //23 / 181 = 0
    16'b00010111_10110110 : OUT <= 0;  //23 / 182 = 0
    16'b00010111_10110111 : OUT <= 0;  //23 / 183 = 0
    16'b00010111_10111000 : OUT <= 0;  //23 / 184 = 0
    16'b00010111_10111001 : OUT <= 0;  //23 / 185 = 0
    16'b00010111_10111010 : OUT <= 0;  //23 / 186 = 0
    16'b00010111_10111011 : OUT <= 0;  //23 / 187 = 0
    16'b00010111_10111100 : OUT <= 0;  //23 / 188 = 0
    16'b00010111_10111101 : OUT <= 0;  //23 / 189 = 0
    16'b00010111_10111110 : OUT <= 0;  //23 / 190 = 0
    16'b00010111_10111111 : OUT <= 0;  //23 / 191 = 0
    16'b00010111_11000000 : OUT <= 0;  //23 / 192 = 0
    16'b00010111_11000001 : OUT <= 0;  //23 / 193 = 0
    16'b00010111_11000010 : OUT <= 0;  //23 / 194 = 0
    16'b00010111_11000011 : OUT <= 0;  //23 / 195 = 0
    16'b00010111_11000100 : OUT <= 0;  //23 / 196 = 0
    16'b00010111_11000101 : OUT <= 0;  //23 / 197 = 0
    16'b00010111_11000110 : OUT <= 0;  //23 / 198 = 0
    16'b00010111_11000111 : OUT <= 0;  //23 / 199 = 0
    16'b00010111_11001000 : OUT <= 0;  //23 / 200 = 0
    16'b00010111_11001001 : OUT <= 0;  //23 / 201 = 0
    16'b00010111_11001010 : OUT <= 0;  //23 / 202 = 0
    16'b00010111_11001011 : OUT <= 0;  //23 / 203 = 0
    16'b00010111_11001100 : OUT <= 0;  //23 / 204 = 0
    16'b00010111_11001101 : OUT <= 0;  //23 / 205 = 0
    16'b00010111_11001110 : OUT <= 0;  //23 / 206 = 0
    16'b00010111_11001111 : OUT <= 0;  //23 / 207 = 0
    16'b00010111_11010000 : OUT <= 0;  //23 / 208 = 0
    16'b00010111_11010001 : OUT <= 0;  //23 / 209 = 0
    16'b00010111_11010010 : OUT <= 0;  //23 / 210 = 0
    16'b00010111_11010011 : OUT <= 0;  //23 / 211 = 0
    16'b00010111_11010100 : OUT <= 0;  //23 / 212 = 0
    16'b00010111_11010101 : OUT <= 0;  //23 / 213 = 0
    16'b00010111_11010110 : OUT <= 0;  //23 / 214 = 0
    16'b00010111_11010111 : OUT <= 0;  //23 / 215 = 0
    16'b00010111_11011000 : OUT <= 0;  //23 / 216 = 0
    16'b00010111_11011001 : OUT <= 0;  //23 / 217 = 0
    16'b00010111_11011010 : OUT <= 0;  //23 / 218 = 0
    16'b00010111_11011011 : OUT <= 0;  //23 / 219 = 0
    16'b00010111_11011100 : OUT <= 0;  //23 / 220 = 0
    16'b00010111_11011101 : OUT <= 0;  //23 / 221 = 0
    16'b00010111_11011110 : OUT <= 0;  //23 / 222 = 0
    16'b00010111_11011111 : OUT <= 0;  //23 / 223 = 0
    16'b00010111_11100000 : OUT <= 0;  //23 / 224 = 0
    16'b00010111_11100001 : OUT <= 0;  //23 / 225 = 0
    16'b00010111_11100010 : OUT <= 0;  //23 / 226 = 0
    16'b00010111_11100011 : OUT <= 0;  //23 / 227 = 0
    16'b00010111_11100100 : OUT <= 0;  //23 / 228 = 0
    16'b00010111_11100101 : OUT <= 0;  //23 / 229 = 0
    16'b00010111_11100110 : OUT <= 0;  //23 / 230 = 0
    16'b00010111_11100111 : OUT <= 0;  //23 / 231 = 0
    16'b00010111_11101000 : OUT <= 0;  //23 / 232 = 0
    16'b00010111_11101001 : OUT <= 0;  //23 / 233 = 0
    16'b00010111_11101010 : OUT <= 0;  //23 / 234 = 0
    16'b00010111_11101011 : OUT <= 0;  //23 / 235 = 0
    16'b00010111_11101100 : OUT <= 0;  //23 / 236 = 0
    16'b00010111_11101101 : OUT <= 0;  //23 / 237 = 0
    16'b00010111_11101110 : OUT <= 0;  //23 / 238 = 0
    16'b00010111_11101111 : OUT <= 0;  //23 / 239 = 0
    16'b00010111_11110000 : OUT <= 0;  //23 / 240 = 0
    16'b00010111_11110001 : OUT <= 0;  //23 / 241 = 0
    16'b00010111_11110010 : OUT <= 0;  //23 / 242 = 0
    16'b00010111_11110011 : OUT <= 0;  //23 / 243 = 0
    16'b00010111_11110100 : OUT <= 0;  //23 / 244 = 0
    16'b00010111_11110101 : OUT <= 0;  //23 / 245 = 0
    16'b00010111_11110110 : OUT <= 0;  //23 / 246 = 0
    16'b00010111_11110111 : OUT <= 0;  //23 / 247 = 0
    16'b00010111_11111000 : OUT <= 0;  //23 / 248 = 0
    16'b00010111_11111001 : OUT <= 0;  //23 / 249 = 0
    16'b00010111_11111010 : OUT <= 0;  //23 / 250 = 0
    16'b00010111_11111011 : OUT <= 0;  //23 / 251 = 0
    16'b00010111_11111100 : OUT <= 0;  //23 / 252 = 0
    16'b00010111_11111101 : OUT <= 0;  //23 / 253 = 0
    16'b00010111_11111110 : OUT <= 0;  //23 / 254 = 0
    16'b00010111_11111111 : OUT <= 0;  //23 / 255 = 0
    16'b00011000_00000000 : OUT <= 0;  //24 / 0 = 0
    16'b00011000_00000001 : OUT <= 24;  //24 / 1 = 24
    16'b00011000_00000010 : OUT <= 12;  //24 / 2 = 12
    16'b00011000_00000011 : OUT <= 8;  //24 / 3 = 8
    16'b00011000_00000100 : OUT <= 6;  //24 / 4 = 6
    16'b00011000_00000101 : OUT <= 4;  //24 / 5 = 4
    16'b00011000_00000110 : OUT <= 4;  //24 / 6 = 4
    16'b00011000_00000111 : OUT <= 3;  //24 / 7 = 3
    16'b00011000_00001000 : OUT <= 3;  //24 / 8 = 3
    16'b00011000_00001001 : OUT <= 2;  //24 / 9 = 2
    16'b00011000_00001010 : OUT <= 2;  //24 / 10 = 2
    16'b00011000_00001011 : OUT <= 2;  //24 / 11 = 2
    16'b00011000_00001100 : OUT <= 2;  //24 / 12 = 2
    16'b00011000_00001101 : OUT <= 1;  //24 / 13 = 1
    16'b00011000_00001110 : OUT <= 1;  //24 / 14 = 1
    16'b00011000_00001111 : OUT <= 1;  //24 / 15 = 1
    16'b00011000_00010000 : OUT <= 1;  //24 / 16 = 1
    16'b00011000_00010001 : OUT <= 1;  //24 / 17 = 1
    16'b00011000_00010010 : OUT <= 1;  //24 / 18 = 1
    16'b00011000_00010011 : OUT <= 1;  //24 / 19 = 1
    16'b00011000_00010100 : OUT <= 1;  //24 / 20 = 1
    16'b00011000_00010101 : OUT <= 1;  //24 / 21 = 1
    16'b00011000_00010110 : OUT <= 1;  //24 / 22 = 1
    16'b00011000_00010111 : OUT <= 1;  //24 / 23 = 1
    16'b00011000_00011000 : OUT <= 1;  //24 / 24 = 1
    16'b00011000_00011001 : OUT <= 0;  //24 / 25 = 0
    16'b00011000_00011010 : OUT <= 0;  //24 / 26 = 0
    16'b00011000_00011011 : OUT <= 0;  //24 / 27 = 0
    16'b00011000_00011100 : OUT <= 0;  //24 / 28 = 0
    16'b00011000_00011101 : OUT <= 0;  //24 / 29 = 0
    16'b00011000_00011110 : OUT <= 0;  //24 / 30 = 0
    16'b00011000_00011111 : OUT <= 0;  //24 / 31 = 0
    16'b00011000_00100000 : OUT <= 0;  //24 / 32 = 0
    16'b00011000_00100001 : OUT <= 0;  //24 / 33 = 0
    16'b00011000_00100010 : OUT <= 0;  //24 / 34 = 0
    16'b00011000_00100011 : OUT <= 0;  //24 / 35 = 0
    16'b00011000_00100100 : OUT <= 0;  //24 / 36 = 0
    16'b00011000_00100101 : OUT <= 0;  //24 / 37 = 0
    16'b00011000_00100110 : OUT <= 0;  //24 / 38 = 0
    16'b00011000_00100111 : OUT <= 0;  //24 / 39 = 0
    16'b00011000_00101000 : OUT <= 0;  //24 / 40 = 0
    16'b00011000_00101001 : OUT <= 0;  //24 / 41 = 0
    16'b00011000_00101010 : OUT <= 0;  //24 / 42 = 0
    16'b00011000_00101011 : OUT <= 0;  //24 / 43 = 0
    16'b00011000_00101100 : OUT <= 0;  //24 / 44 = 0
    16'b00011000_00101101 : OUT <= 0;  //24 / 45 = 0
    16'b00011000_00101110 : OUT <= 0;  //24 / 46 = 0
    16'b00011000_00101111 : OUT <= 0;  //24 / 47 = 0
    16'b00011000_00110000 : OUT <= 0;  //24 / 48 = 0
    16'b00011000_00110001 : OUT <= 0;  //24 / 49 = 0
    16'b00011000_00110010 : OUT <= 0;  //24 / 50 = 0
    16'b00011000_00110011 : OUT <= 0;  //24 / 51 = 0
    16'b00011000_00110100 : OUT <= 0;  //24 / 52 = 0
    16'b00011000_00110101 : OUT <= 0;  //24 / 53 = 0
    16'b00011000_00110110 : OUT <= 0;  //24 / 54 = 0
    16'b00011000_00110111 : OUT <= 0;  //24 / 55 = 0
    16'b00011000_00111000 : OUT <= 0;  //24 / 56 = 0
    16'b00011000_00111001 : OUT <= 0;  //24 / 57 = 0
    16'b00011000_00111010 : OUT <= 0;  //24 / 58 = 0
    16'b00011000_00111011 : OUT <= 0;  //24 / 59 = 0
    16'b00011000_00111100 : OUT <= 0;  //24 / 60 = 0
    16'b00011000_00111101 : OUT <= 0;  //24 / 61 = 0
    16'b00011000_00111110 : OUT <= 0;  //24 / 62 = 0
    16'b00011000_00111111 : OUT <= 0;  //24 / 63 = 0
    16'b00011000_01000000 : OUT <= 0;  //24 / 64 = 0
    16'b00011000_01000001 : OUT <= 0;  //24 / 65 = 0
    16'b00011000_01000010 : OUT <= 0;  //24 / 66 = 0
    16'b00011000_01000011 : OUT <= 0;  //24 / 67 = 0
    16'b00011000_01000100 : OUT <= 0;  //24 / 68 = 0
    16'b00011000_01000101 : OUT <= 0;  //24 / 69 = 0
    16'b00011000_01000110 : OUT <= 0;  //24 / 70 = 0
    16'b00011000_01000111 : OUT <= 0;  //24 / 71 = 0
    16'b00011000_01001000 : OUT <= 0;  //24 / 72 = 0
    16'b00011000_01001001 : OUT <= 0;  //24 / 73 = 0
    16'b00011000_01001010 : OUT <= 0;  //24 / 74 = 0
    16'b00011000_01001011 : OUT <= 0;  //24 / 75 = 0
    16'b00011000_01001100 : OUT <= 0;  //24 / 76 = 0
    16'b00011000_01001101 : OUT <= 0;  //24 / 77 = 0
    16'b00011000_01001110 : OUT <= 0;  //24 / 78 = 0
    16'b00011000_01001111 : OUT <= 0;  //24 / 79 = 0
    16'b00011000_01010000 : OUT <= 0;  //24 / 80 = 0
    16'b00011000_01010001 : OUT <= 0;  //24 / 81 = 0
    16'b00011000_01010010 : OUT <= 0;  //24 / 82 = 0
    16'b00011000_01010011 : OUT <= 0;  //24 / 83 = 0
    16'b00011000_01010100 : OUT <= 0;  //24 / 84 = 0
    16'b00011000_01010101 : OUT <= 0;  //24 / 85 = 0
    16'b00011000_01010110 : OUT <= 0;  //24 / 86 = 0
    16'b00011000_01010111 : OUT <= 0;  //24 / 87 = 0
    16'b00011000_01011000 : OUT <= 0;  //24 / 88 = 0
    16'b00011000_01011001 : OUT <= 0;  //24 / 89 = 0
    16'b00011000_01011010 : OUT <= 0;  //24 / 90 = 0
    16'b00011000_01011011 : OUT <= 0;  //24 / 91 = 0
    16'b00011000_01011100 : OUT <= 0;  //24 / 92 = 0
    16'b00011000_01011101 : OUT <= 0;  //24 / 93 = 0
    16'b00011000_01011110 : OUT <= 0;  //24 / 94 = 0
    16'b00011000_01011111 : OUT <= 0;  //24 / 95 = 0
    16'b00011000_01100000 : OUT <= 0;  //24 / 96 = 0
    16'b00011000_01100001 : OUT <= 0;  //24 / 97 = 0
    16'b00011000_01100010 : OUT <= 0;  //24 / 98 = 0
    16'b00011000_01100011 : OUT <= 0;  //24 / 99 = 0
    16'b00011000_01100100 : OUT <= 0;  //24 / 100 = 0
    16'b00011000_01100101 : OUT <= 0;  //24 / 101 = 0
    16'b00011000_01100110 : OUT <= 0;  //24 / 102 = 0
    16'b00011000_01100111 : OUT <= 0;  //24 / 103 = 0
    16'b00011000_01101000 : OUT <= 0;  //24 / 104 = 0
    16'b00011000_01101001 : OUT <= 0;  //24 / 105 = 0
    16'b00011000_01101010 : OUT <= 0;  //24 / 106 = 0
    16'b00011000_01101011 : OUT <= 0;  //24 / 107 = 0
    16'b00011000_01101100 : OUT <= 0;  //24 / 108 = 0
    16'b00011000_01101101 : OUT <= 0;  //24 / 109 = 0
    16'b00011000_01101110 : OUT <= 0;  //24 / 110 = 0
    16'b00011000_01101111 : OUT <= 0;  //24 / 111 = 0
    16'b00011000_01110000 : OUT <= 0;  //24 / 112 = 0
    16'b00011000_01110001 : OUT <= 0;  //24 / 113 = 0
    16'b00011000_01110010 : OUT <= 0;  //24 / 114 = 0
    16'b00011000_01110011 : OUT <= 0;  //24 / 115 = 0
    16'b00011000_01110100 : OUT <= 0;  //24 / 116 = 0
    16'b00011000_01110101 : OUT <= 0;  //24 / 117 = 0
    16'b00011000_01110110 : OUT <= 0;  //24 / 118 = 0
    16'b00011000_01110111 : OUT <= 0;  //24 / 119 = 0
    16'b00011000_01111000 : OUT <= 0;  //24 / 120 = 0
    16'b00011000_01111001 : OUT <= 0;  //24 / 121 = 0
    16'b00011000_01111010 : OUT <= 0;  //24 / 122 = 0
    16'b00011000_01111011 : OUT <= 0;  //24 / 123 = 0
    16'b00011000_01111100 : OUT <= 0;  //24 / 124 = 0
    16'b00011000_01111101 : OUT <= 0;  //24 / 125 = 0
    16'b00011000_01111110 : OUT <= 0;  //24 / 126 = 0
    16'b00011000_01111111 : OUT <= 0;  //24 / 127 = 0
    16'b00011000_10000000 : OUT <= 0;  //24 / 128 = 0
    16'b00011000_10000001 : OUT <= 0;  //24 / 129 = 0
    16'b00011000_10000010 : OUT <= 0;  //24 / 130 = 0
    16'b00011000_10000011 : OUT <= 0;  //24 / 131 = 0
    16'b00011000_10000100 : OUT <= 0;  //24 / 132 = 0
    16'b00011000_10000101 : OUT <= 0;  //24 / 133 = 0
    16'b00011000_10000110 : OUT <= 0;  //24 / 134 = 0
    16'b00011000_10000111 : OUT <= 0;  //24 / 135 = 0
    16'b00011000_10001000 : OUT <= 0;  //24 / 136 = 0
    16'b00011000_10001001 : OUT <= 0;  //24 / 137 = 0
    16'b00011000_10001010 : OUT <= 0;  //24 / 138 = 0
    16'b00011000_10001011 : OUT <= 0;  //24 / 139 = 0
    16'b00011000_10001100 : OUT <= 0;  //24 / 140 = 0
    16'b00011000_10001101 : OUT <= 0;  //24 / 141 = 0
    16'b00011000_10001110 : OUT <= 0;  //24 / 142 = 0
    16'b00011000_10001111 : OUT <= 0;  //24 / 143 = 0
    16'b00011000_10010000 : OUT <= 0;  //24 / 144 = 0
    16'b00011000_10010001 : OUT <= 0;  //24 / 145 = 0
    16'b00011000_10010010 : OUT <= 0;  //24 / 146 = 0
    16'b00011000_10010011 : OUT <= 0;  //24 / 147 = 0
    16'b00011000_10010100 : OUT <= 0;  //24 / 148 = 0
    16'b00011000_10010101 : OUT <= 0;  //24 / 149 = 0
    16'b00011000_10010110 : OUT <= 0;  //24 / 150 = 0
    16'b00011000_10010111 : OUT <= 0;  //24 / 151 = 0
    16'b00011000_10011000 : OUT <= 0;  //24 / 152 = 0
    16'b00011000_10011001 : OUT <= 0;  //24 / 153 = 0
    16'b00011000_10011010 : OUT <= 0;  //24 / 154 = 0
    16'b00011000_10011011 : OUT <= 0;  //24 / 155 = 0
    16'b00011000_10011100 : OUT <= 0;  //24 / 156 = 0
    16'b00011000_10011101 : OUT <= 0;  //24 / 157 = 0
    16'b00011000_10011110 : OUT <= 0;  //24 / 158 = 0
    16'b00011000_10011111 : OUT <= 0;  //24 / 159 = 0
    16'b00011000_10100000 : OUT <= 0;  //24 / 160 = 0
    16'b00011000_10100001 : OUT <= 0;  //24 / 161 = 0
    16'b00011000_10100010 : OUT <= 0;  //24 / 162 = 0
    16'b00011000_10100011 : OUT <= 0;  //24 / 163 = 0
    16'b00011000_10100100 : OUT <= 0;  //24 / 164 = 0
    16'b00011000_10100101 : OUT <= 0;  //24 / 165 = 0
    16'b00011000_10100110 : OUT <= 0;  //24 / 166 = 0
    16'b00011000_10100111 : OUT <= 0;  //24 / 167 = 0
    16'b00011000_10101000 : OUT <= 0;  //24 / 168 = 0
    16'b00011000_10101001 : OUT <= 0;  //24 / 169 = 0
    16'b00011000_10101010 : OUT <= 0;  //24 / 170 = 0
    16'b00011000_10101011 : OUT <= 0;  //24 / 171 = 0
    16'b00011000_10101100 : OUT <= 0;  //24 / 172 = 0
    16'b00011000_10101101 : OUT <= 0;  //24 / 173 = 0
    16'b00011000_10101110 : OUT <= 0;  //24 / 174 = 0
    16'b00011000_10101111 : OUT <= 0;  //24 / 175 = 0
    16'b00011000_10110000 : OUT <= 0;  //24 / 176 = 0
    16'b00011000_10110001 : OUT <= 0;  //24 / 177 = 0
    16'b00011000_10110010 : OUT <= 0;  //24 / 178 = 0
    16'b00011000_10110011 : OUT <= 0;  //24 / 179 = 0
    16'b00011000_10110100 : OUT <= 0;  //24 / 180 = 0
    16'b00011000_10110101 : OUT <= 0;  //24 / 181 = 0
    16'b00011000_10110110 : OUT <= 0;  //24 / 182 = 0
    16'b00011000_10110111 : OUT <= 0;  //24 / 183 = 0
    16'b00011000_10111000 : OUT <= 0;  //24 / 184 = 0
    16'b00011000_10111001 : OUT <= 0;  //24 / 185 = 0
    16'b00011000_10111010 : OUT <= 0;  //24 / 186 = 0
    16'b00011000_10111011 : OUT <= 0;  //24 / 187 = 0
    16'b00011000_10111100 : OUT <= 0;  //24 / 188 = 0
    16'b00011000_10111101 : OUT <= 0;  //24 / 189 = 0
    16'b00011000_10111110 : OUT <= 0;  //24 / 190 = 0
    16'b00011000_10111111 : OUT <= 0;  //24 / 191 = 0
    16'b00011000_11000000 : OUT <= 0;  //24 / 192 = 0
    16'b00011000_11000001 : OUT <= 0;  //24 / 193 = 0
    16'b00011000_11000010 : OUT <= 0;  //24 / 194 = 0
    16'b00011000_11000011 : OUT <= 0;  //24 / 195 = 0
    16'b00011000_11000100 : OUT <= 0;  //24 / 196 = 0
    16'b00011000_11000101 : OUT <= 0;  //24 / 197 = 0
    16'b00011000_11000110 : OUT <= 0;  //24 / 198 = 0
    16'b00011000_11000111 : OUT <= 0;  //24 / 199 = 0
    16'b00011000_11001000 : OUT <= 0;  //24 / 200 = 0
    16'b00011000_11001001 : OUT <= 0;  //24 / 201 = 0
    16'b00011000_11001010 : OUT <= 0;  //24 / 202 = 0
    16'b00011000_11001011 : OUT <= 0;  //24 / 203 = 0
    16'b00011000_11001100 : OUT <= 0;  //24 / 204 = 0
    16'b00011000_11001101 : OUT <= 0;  //24 / 205 = 0
    16'b00011000_11001110 : OUT <= 0;  //24 / 206 = 0
    16'b00011000_11001111 : OUT <= 0;  //24 / 207 = 0
    16'b00011000_11010000 : OUT <= 0;  //24 / 208 = 0
    16'b00011000_11010001 : OUT <= 0;  //24 / 209 = 0
    16'b00011000_11010010 : OUT <= 0;  //24 / 210 = 0
    16'b00011000_11010011 : OUT <= 0;  //24 / 211 = 0
    16'b00011000_11010100 : OUT <= 0;  //24 / 212 = 0
    16'b00011000_11010101 : OUT <= 0;  //24 / 213 = 0
    16'b00011000_11010110 : OUT <= 0;  //24 / 214 = 0
    16'b00011000_11010111 : OUT <= 0;  //24 / 215 = 0
    16'b00011000_11011000 : OUT <= 0;  //24 / 216 = 0
    16'b00011000_11011001 : OUT <= 0;  //24 / 217 = 0
    16'b00011000_11011010 : OUT <= 0;  //24 / 218 = 0
    16'b00011000_11011011 : OUT <= 0;  //24 / 219 = 0
    16'b00011000_11011100 : OUT <= 0;  //24 / 220 = 0
    16'b00011000_11011101 : OUT <= 0;  //24 / 221 = 0
    16'b00011000_11011110 : OUT <= 0;  //24 / 222 = 0
    16'b00011000_11011111 : OUT <= 0;  //24 / 223 = 0
    16'b00011000_11100000 : OUT <= 0;  //24 / 224 = 0
    16'b00011000_11100001 : OUT <= 0;  //24 / 225 = 0
    16'b00011000_11100010 : OUT <= 0;  //24 / 226 = 0
    16'b00011000_11100011 : OUT <= 0;  //24 / 227 = 0
    16'b00011000_11100100 : OUT <= 0;  //24 / 228 = 0
    16'b00011000_11100101 : OUT <= 0;  //24 / 229 = 0
    16'b00011000_11100110 : OUT <= 0;  //24 / 230 = 0
    16'b00011000_11100111 : OUT <= 0;  //24 / 231 = 0
    16'b00011000_11101000 : OUT <= 0;  //24 / 232 = 0
    16'b00011000_11101001 : OUT <= 0;  //24 / 233 = 0
    16'b00011000_11101010 : OUT <= 0;  //24 / 234 = 0
    16'b00011000_11101011 : OUT <= 0;  //24 / 235 = 0
    16'b00011000_11101100 : OUT <= 0;  //24 / 236 = 0
    16'b00011000_11101101 : OUT <= 0;  //24 / 237 = 0
    16'b00011000_11101110 : OUT <= 0;  //24 / 238 = 0
    16'b00011000_11101111 : OUT <= 0;  //24 / 239 = 0
    16'b00011000_11110000 : OUT <= 0;  //24 / 240 = 0
    16'b00011000_11110001 : OUT <= 0;  //24 / 241 = 0
    16'b00011000_11110010 : OUT <= 0;  //24 / 242 = 0
    16'b00011000_11110011 : OUT <= 0;  //24 / 243 = 0
    16'b00011000_11110100 : OUT <= 0;  //24 / 244 = 0
    16'b00011000_11110101 : OUT <= 0;  //24 / 245 = 0
    16'b00011000_11110110 : OUT <= 0;  //24 / 246 = 0
    16'b00011000_11110111 : OUT <= 0;  //24 / 247 = 0
    16'b00011000_11111000 : OUT <= 0;  //24 / 248 = 0
    16'b00011000_11111001 : OUT <= 0;  //24 / 249 = 0
    16'b00011000_11111010 : OUT <= 0;  //24 / 250 = 0
    16'b00011000_11111011 : OUT <= 0;  //24 / 251 = 0
    16'b00011000_11111100 : OUT <= 0;  //24 / 252 = 0
    16'b00011000_11111101 : OUT <= 0;  //24 / 253 = 0
    16'b00011000_11111110 : OUT <= 0;  //24 / 254 = 0
    16'b00011000_11111111 : OUT <= 0;  //24 / 255 = 0
    16'b00011001_00000000 : OUT <= 0;  //25 / 0 = 0
    16'b00011001_00000001 : OUT <= 25;  //25 / 1 = 25
    16'b00011001_00000010 : OUT <= 12;  //25 / 2 = 12
    16'b00011001_00000011 : OUT <= 8;  //25 / 3 = 8
    16'b00011001_00000100 : OUT <= 6;  //25 / 4 = 6
    16'b00011001_00000101 : OUT <= 5;  //25 / 5 = 5
    16'b00011001_00000110 : OUT <= 4;  //25 / 6 = 4
    16'b00011001_00000111 : OUT <= 3;  //25 / 7 = 3
    16'b00011001_00001000 : OUT <= 3;  //25 / 8 = 3
    16'b00011001_00001001 : OUT <= 2;  //25 / 9 = 2
    16'b00011001_00001010 : OUT <= 2;  //25 / 10 = 2
    16'b00011001_00001011 : OUT <= 2;  //25 / 11 = 2
    16'b00011001_00001100 : OUT <= 2;  //25 / 12 = 2
    16'b00011001_00001101 : OUT <= 1;  //25 / 13 = 1
    16'b00011001_00001110 : OUT <= 1;  //25 / 14 = 1
    16'b00011001_00001111 : OUT <= 1;  //25 / 15 = 1
    16'b00011001_00010000 : OUT <= 1;  //25 / 16 = 1
    16'b00011001_00010001 : OUT <= 1;  //25 / 17 = 1
    16'b00011001_00010010 : OUT <= 1;  //25 / 18 = 1
    16'b00011001_00010011 : OUT <= 1;  //25 / 19 = 1
    16'b00011001_00010100 : OUT <= 1;  //25 / 20 = 1
    16'b00011001_00010101 : OUT <= 1;  //25 / 21 = 1
    16'b00011001_00010110 : OUT <= 1;  //25 / 22 = 1
    16'b00011001_00010111 : OUT <= 1;  //25 / 23 = 1
    16'b00011001_00011000 : OUT <= 1;  //25 / 24 = 1
    16'b00011001_00011001 : OUT <= 1;  //25 / 25 = 1
    16'b00011001_00011010 : OUT <= 0;  //25 / 26 = 0
    16'b00011001_00011011 : OUT <= 0;  //25 / 27 = 0
    16'b00011001_00011100 : OUT <= 0;  //25 / 28 = 0
    16'b00011001_00011101 : OUT <= 0;  //25 / 29 = 0
    16'b00011001_00011110 : OUT <= 0;  //25 / 30 = 0
    16'b00011001_00011111 : OUT <= 0;  //25 / 31 = 0
    16'b00011001_00100000 : OUT <= 0;  //25 / 32 = 0
    16'b00011001_00100001 : OUT <= 0;  //25 / 33 = 0
    16'b00011001_00100010 : OUT <= 0;  //25 / 34 = 0
    16'b00011001_00100011 : OUT <= 0;  //25 / 35 = 0
    16'b00011001_00100100 : OUT <= 0;  //25 / 36 = 0
    16'b00011001_00100101 : OUT <= 0;  //25 / 37 = 0
    16'b00011001_00100110 : OUT <= 0;  //25 / 38 = 0
    16'b00011001_00100111 : OUT <= 0;  //25 / 39 = 0
    16'b00011001_00101000 : OUT <= 0;  //25 / 40 = 0
    16'b00011001_00101001 : OUT <= 0;  //25 / 41 = 0
    16'b00011001_00101010 : OUT <= 0;  //25 / 42 = 0
    16'b00011001_00101011 : OUT <= 0;  //25 / 43 = 0
    16'b00011001_00101100 : OUT <= 0;  //25 / 44 = 0
    16'b00011001_00101101 : OUT <= 0;  //25 / 45 = 0
    16'b00011001_00101110 : OUT <= 0;  //25 / 46 = 0
    16'b00011001_00101111 : OUT <= 0;  //25 / 47 = 0
    16'b00011001_00110000 : OUT <= 0;  //25 / 48 = 0
    16'b00011001_00110001 : OUT <= 0;  //25 / 49 = 0
    16'b00011001_00110010 : OUT <= 0;  //25 / 50 = 0
    16'b00011001_00110011 : OUT <= 0;  //25 / 51 = 0
    16'b00011001_00110100 : OUT <= 0;  //25 / 52 = 0
    16'b00011001_00110101 : OUT <= 0;  //25 / 53 = 0
    16'b00011001_00110110 : OUT <= 0;  //25 / 54 = 0
    16'b00011001_00110111 : OUT <= 0;  //25 / 55 = 0
    16'b00011001_00111000 : OUT <= 0;  //25 / 56 = 0
    16'b00011001_00111001 : OUT <= 0;  //25 / 57 = 0
    16'b00011001_00111010 : OUT <= 0;  //25 / 58 = 0
    16'b00011001_00111011 : OUT <= 0;  //25 / 59 = 0
    16'b00011001_00111100 : OUT <= 0;  //25 / 60 = 0
    16'b00011001_00111101 : OUT <= 0;  //25 / 61 = 0
    16'b00011001_00111110 : OUT <= 0;  //25 / 62 = 0
    16'b00011001_00111111 : OUT <= 0;  //25 / 63 = 0
    16'b00011001_01000000 : OUT <= 0;  //25 / 64 = 0
    16'b00011001_01000001 : OUT <= 0;  //25 / 65 = 0
    16'b00011001_01000010 : OUT <= 0;  //25 / 66 = 0
    16'b00011001_01000011 : OUT <= 0;  //25 / 67 = 0
    16'b00011001_01000100 : OUT <= 0;  //25 / 68 = 0
    16'b00011001_01000101 : OUT <= 0;  //25 / 69 = 0
    16'b00011001_01000110 : OUT <= 0;  //25 / 70 = 0
    16'b00011001_01000111 : OUT <= 0;  //25 / 71 = 0
    16'b00011001_01001000 : OUT <= 0;  //25 / 72 = 0
    16'b00011001_01001001 : OUT <= 0;  //25 / 73 = 0
    16'b00011001_01001010 : OUT <= 0;  //25 / 74 = 0
    16'b00011001_01001011 : OUT <= 0;  //25 / 75 = 0
    16'b00011001_01001100 : OUT <= 0;  //25 / 76 = 0
    16'b00011001_01001101 : OUT <= 0;  //25 / 77 = 0
    16'b00011001_01001110 : OUT <= 0;  //25 / 78 = 0
    16'b00011001_01001111 : OUT <= 0;  //25 / 79 = 0
    16'b00011001_01010000 : OUT <= 0;  //25 / 80 = 0
    16'b00011001_01010001 : OUT <= 0;  //25 / 81 = 0
    16'b00011001_01010010 : OUT <= 0;  //25 / 82 = 0
    16'b00011001_01010011 : OUT <= 0;  //25 / 83 = 0
    16'b00011001_01010100 : OUT <= 0;  //25 / 84 = 0
    16'b00011001_01010101 : OUT <= 0;  //25 / 85 = 0
    16'b00011001_01010110 : OUT <= 0;  //25 / 86 = 0
    16'b00011001_01010111 : OUT <= 0;  //25 / 87 = 0
    16'b00011001_01011000 : OUT <= 0;  //25 / 88 = 0
    16'b00011001_01011001 : OUT <= 0;  //25 / 89 = 0
    16'b00011001_01011010 : OUT <= 0;  //25 / 90 = 0
    16'b00011001_01011011 : OUT <= 0;  //25 / 91 = 0
    16'b00011001_01011100 : OUT <= 0;  //25 / 92 = 0
    16'b00011001_01011101 : OUT <= 0;  //25 / 93 = 0
    16'b00011001_01011110 : OUT <= 0;  //25 / 94 = 0
    16'b00011001_01011111 : OUT <= 0;  //25 / 95 = 0
    16'b00011001_01100000 : OUT <= 0;  //25 / 96 = 0
    16'b00011001_01100001 : OUT <= 0;  //25 / 97 = 0
    16'b00011001_01100010 : OUT <= 0;  //25 / 98 = 0
    16'b00011001_01100011 : OUT <= 0;  //25 / 99 = 0
    16'b00011001_01100100 : OUT <= 0;  //25 / 100 = 0
    16'b00011001_01100101 : OUT <= 0;  //25 / 101 = 0
    16'b00011001_01100110 : OUT <= 0;  //25 / 102 = 0
    16'b00011001_01100111 : OUT <= 0;  //25 / 103 = 0
    16'b00011001_01101000 : OUT <= 0;  //25 / 104 = 0
    16'b00011001_01101001 : OUT <= 0;  //25 / 105 = 0
    16'b00011001_01101010 : OUT <= 0;  //25 / 106 = 0
    16'b00011001_01101011 : OUT <= 0;  //25 / 107 = 0
    16'b00011001_01101100 : OUT <= 0;  //25 / 108 = 0
    16'b00011001_01101101 : OUT <= 0;  //25 / 109 = 0
    16'b00011001_01101110 : OUT <= 0;  //25 / 110 = 0
    16'b00011001_01101111 : OUT <= 0;  //25 / 111 = 0
    16'b00011001_01110000 : OUT <= 0;  //25 / 112 = 0
    16'b00011001_01110001 : OUT <= 0;  //25 / 113 = 0
    16'b00011001_01110010 : OUT <= 0;  //25 / 114 = 0
    16'b00011001_01110011 : OUT <= 0;  //25 / 115 = 0
    16'b00011001_01110100 : OUT <= 0;  //25 / 116 = 0
    16'b00011001_01110101 : OUT <= 0;  //25 / 117 = 0
    16'b00011001_01110110 : OUT <= 0;  //25 / 118 = 0
    16'b00011001_01110111 : OUT <= 0;  //25 / 119 = 0
    16'b00011001_01111000 : OUT <= 0;  //25 / 120 = 0
    16'b00011001_01111001 : OUT <= 0;  //25 / 121 = 0
    16'b00011001_01111010 : OUT <= 0;  //25 / 122 = 0
    16'b00011001_01111011 : OUT <= 0;  //25 / 123 = 0
    16'b00011001_01111100 : OUT <= 0;  //25 / 124 = 0
    16'b00011001_01111101 : OUT <= 0;  //25 / 125 = 0
    16'b00011001_01111110 : OUT <= 0;  //25 / 126 = 0
    16'b00011001_01111111 : OUT <= 0;  //25 / 127 = 0
    16'b00011001_10000000 : OUT <= 0;  //25 / 128 = 0
    16'b00011001_10000001 : OUT <= 0;  //25 / 129 = 0
    16'b00011001_10000010 : OUT <= 0;  //25 / 130 = 0
    16'b00011001_10000011 : OUT <= 0;  //25 / 131 = 0
    16'b00011001_10000100 : OUT <= 0;  //25 / 132 = 0
    16'b00011001_10000101 : OUT <= 0;  //25 / 133 = 0
    16'b00011001_10000110 : OUT <= 0;  //25 / 134 = 0
    16'b00011001_10000111 : OUT <= 0;  //25 / 135 = 0
    16'b00011001_10001000 : OUT <= 0;  //25 / 136 = 0
    16'b00011001_10001001 : OUT <= 0;  //25 / 137 = 0
    16'b00011001_10001010 : OUT <= 0;  //25 / 138 = 0
    16'b00011001_10001011 : OUT <= 0;  //25 / 139 = 0
    16'b00011001_10001100 : OUT <= 0;  //25 / 140 = 0
    16'b00011001_10001101 : OUT <= 0;  //25 / 141 = 0
    16'b00011001_10001110 : OUT <= 0;  //25 / 142 = 0
    16'b00011001_10001111 : OUT <= 0;  //25 / 143 = 0
    16'b00011001_10010000 : OUT <= 0;  //25 / 144 = 0
    16'b00011001_10010001 : OUT <= 0;  //25 / 145 = 0
    16'b00011001_10010010 : OUT <= 0;  //25 / 146 = 0
    16'b00011001_10010011 : OUT <= 0;  //25 / 147 = 0
    16'b00011001_10010100 : OUT <= 0;  //25 / 148 = 0
    16'b00011001_10010101 : OUT <= 0;  //25 / 149 = 0
    16'b00011001_10010110 : OUT <= 0;  //25 / 150 = 0
    16'b00011001_10010111 : OUT <= 0;  //25 / 151 = 0
    16'b00011001_10011000 : OUT <= 0;  //25 / 152 = 0
    16'b00011001_10011001 : OUT <= 0;  //25 / 153 = 0
    16'b00011001_10011010 : OUT <= 0;  //25 / 154 = 0
    16'b00011001_10011011 : OUT <= 0;  //25 / 155 = 0
    16'b00011001_10011100 : OUT <= 0;  //25 / 156 = 0
    16'b00011001_10011101 : OUT <= 0;  //25 / 157 = 0
    16'b00011001_10011110 : OUT <= 0;  //25 / 158 = 0
    16'b00011001_10011111 : OUT <= 0;  //25 / 159 = 0
    16'b00011001_10100000 : OUT <= 0;  //25 / 160 = 0
    16'b00011001_10100001 : OUT <= 0;  //25 / 161 = 0
    16'b00011001_10100010 : OUT <= 0;  //25 / 162 = 0
    16'b00011001_10100011 : OUT <= 0;  //25 / 163 = 0
    16'b00011001_10100100 : OUT <= 0;  //25 / 164 = 0
    16'b00011001_10100101 : OUT <= 0;  //25 / 165 = 0
    16'b00011001_10100110 : OUT <= 0;  //25 / 166 = 0
    16'b00011001_10100111 : OUT <= 0;  //25 / 167 = 0
    16'b00011001_10101000 : OUT <= 0;  //25 / 168 = 0
    16'b00011001_10101001 : OUT <= 0;  //25 / 169 = 0
    16'b00011001_10101010 : OUT <= 0;  //25 / 170 = 0
    16'b00011001_10101011 : OUT <= 0;  //25 / 171 = 0
    16'b00011001_10101100 : OUT <= 0;  //25 / 172 = 0
    16'b00011001_10101101 : OUT <= 0;  //25 / 173 = 0
    16'b00011001_10101110 : OUT <= 0;  //25 / 174 = 0
    16'b00011001_10101111 : OUT <= 0;  //25 / 175 = 0
    16'b00011001_10110000 : OUT <= 0;  //25 / 176 = 0
    16'b00011001_10110001 : OUT <= 0;  //25 / 177 = 0
    16'b00011001_10110010 : OUT <= 0;  //25 / 178 = 0
    16'b00011001_10110011 : OUT <= 0;  //25 / 179 = 0
    16'b00011001_10110100 : OUT <= 0;  //25 / 180 = 0
    16'b00011001_10110101 : OUT <= 0;  //25 / 181 = 0
    16'b00011001_10110110 : OUT <= 0;  //25 / 182 = 0
    16'b00011001_10110111 : OUT <= 0;  //25 / 183 = 0
    16'b00011001_10111000 : OUT <= 0;  //25 / 184 = 0
    16'b00011001_10111001 : OUT <= 0;  //25 / 185 = 0
    16'b00011001_10111010 : OUT <= 0;  //25 / 186 = 0
    16'b00011001_10111011 : OUT <= 0;  //25 / 187 = 0
    16'b00011001_10111100 : OUT <= 0;  //25 / 188 = 0
    16'b00011001_10111101 : OUT <= 0;  //25 / 189 = 0
    16'b00011001_10111110 : OUT <= 0;  //25 / 190 = 0
    16'b00011001_10111111 : OUT <= 0;  //25 / 191 = 0
    16'b00011001_11000000 : OUT <= 0;  //25 / 192 = 0
    16'b00011001_11000001 : OUT <= 0;  //25 / 193 = 0
    16'b00011001_11000010 : OUT <= 0;  //25 / 194 = 0
    16'b00011001_11000011 : OUT <= 0;  //25 / 195 = 0
    16'b00011001_11000100 : OUT <= 0;  //25 / 196 = 0
    16'b00011001_11000101 : OUT <= 0;  //25 / 197 = 0
    16'b00011001_11000110 : OUT <= 0;  //25 / 198 = 0
    16'b00011001_11000111 : OUT <= 0;  //25 / 199 = 0
    16'b00011001_11001000 : OUT <= 0;  //25 / 200 = 0
    16'b00011001_11001001 : OUT <= 0;  //25 / 201 = 0
    16'b00011001_11001010 : OUT <= 0;  //25 / 202 = 0
    16'b00011001_11001011 : OUT <= 0;  //25 / 203 = 0
    16'b00011001_11001100 : OUT <= 0;  //25 / 204 = 0
    16'b00011001_11001101 : OUT <= 0;  //25 / 205 = 0
    16'b00011001_11001110 : OUT <= 0;  //25 / 206 = 0
    16'b00011001_11001111 : OUT <= 0;  //25 / 207 = 0
    16'b00011001_11010000 : OUT <= 0;  //25 / 208 = 0
    16'b00011001_11010001 : OUT <= 0;  //25 / 209 = 0
    16'b00011001_11010010 : OUT <= 0;  //25 / 210 = 0
    16'b00011001_11010011 : OUT <= 0;  //25 / 211 = 0
    16'b00011001_11010100 : OUT <= 0;  //25 / 212 = 0
    16'b00011001_11010101 : OUT <= 0;  //25 / 213 = 0
    16'b00011001_11010110 : OUT <= 0;  //25 / 214 = 0
    16'b00011001_11010111 : OUT <= 0;  //25 / 215 = 0
    16'b00011001_11011000 : OUT <= 0;  //25 / 216 = 0
    16'b00011001_11011001 : OUT <= 0;  //25 / 217 = 0
    16'b00011001_11011010 : OUT <= 0;  //25 / 218 = 0
    16'b00011001_11011011 : OUT <= 0;  //25 / 219 = 0
    16'b00011001_11011100 : OUT <= 0;  //25 / 220 = 0
    16'b00011001_11011101 : OUT <= 0;  //25 / 221 = 0
    16'b00011001_11011110 : OUT <= 0;  //25 / 222 = 0
    16'b00011001_11011111 : OUT <= 0;  //25 / 223 = 0
    16'b00011001_11100000 : OUT <= 0;  //25 / 224 = 0
    16'b00011001_11100001 : OUT <= 0;  //25 / 225 = 0
    16'b00011001_11100010 : OUT <= 0;  //25 / 226 = 0
    16'b00011001_11100011 : OUT <= 0;  //25 / 227 = 0
    16'b00011001_11100100 : OUT <= 0;  //25 / 228 = 0
    16'b00011001_11100101 : OUT <= 0;  //25 / 229 = 0
    16'b00011001_11100110 : OUT <= 0;  //25 / 230 = 0
    16'b00011001_11100111 : OUT <= 0;  //25 / 231 = 0
    16'b00011001_11101000 : OUT <= 0;  //25 / 232 = 0
    16'b00011001_11101001 : OUT <= 0;  //25 / 233 = 0
    16'b00011001_11101010 : OUT <= 0;  //25 / 234 = 0
    16'b00011001_11101011 : OUT <= 0;  //25 / 235 = 0
    16'b00011001_11101100 : OUT <= 0;  //25 / 236 = 0
    16'b00011001_11101101 : OUT <= 0;  //25 / 237 = 0
    16'b00011001_11101110 : OUT <= 0;  //25 / 238 = 0
    16'b00011001_11101111 : OUT <= 0;  //25 / 239 = 0
    16'b00011001_11110000 : OUT <= 0;  //25 / 240 = 0
    16'b00011001_11110001 : OUT <= 0;  //25 / 241 = 0
    16'b00011001_11110010 : OUT <= 0;  //25 / 242 = 0
    16'b00011001_11110011 : OUT <= 0;  //25 / 243 = 0
    16'b00011001_11110100 : OUT <= 0;  //25 / 244 = 0
    16'b00011001_11110101 : OUT <= 0;  //25 / 245 = 0
    16'b00011001_11110110 : OUT <= 0;  //25 / 246 = 0
    16'b00011001_11110111 : OUT <= 0;  //25 / 247 = 0
    16'b00011001_11111000 : OUT <= 0;  //25 / 248 = 0
    16'b00011001_11111001 : OUT <= 0;  //25 / 249 = 0
    16'b00011001_11111010 : OUT <= 0;  //25 / 250 = 0
    16'b00011001_11111011 : OUT <= 0;  //25 / 251 = 0
    16'b00011001_11111100 : OUT <= 0;  //25 / 252 = 0
    16'b00011001_11111101 : OUT <= 0;  //25 / 253 = 0
    16'b00011001_11111110 : OUT <= 0;  //25 / 254 = 0
    16'b00011001_11111111 : OUT <= 0;  //25 / 255 = 0
    16'b00011010_00000000 : OUT <= 0;  //26 / 0 = 0
    16'b00011010_00000001 : OUT <= 26;  //26 / 1 = 26
    16'b00011010_00000010 : OUT <= 13;  //26 / 2 = 13
    16'b00011010_00000011 : OUT <= 8;  //26 / 3 = 8
    16'b00011010_00000100 : OUT <= 6;  //26 / 4 = 6
    16'b00011010_00000101 : OUT <= 5;  //26 / 5 = 5
    16'b00011010_00000110 : OUT <= 4;  //26 / 6 = 4
    16'b00011010_00000111 : OUT <= 3;  //26 / 7 = 3
    16'b00011010_00001000 : OUT <= 3;  //26 / 8 = 3
    16'b00011010_00001001 : OUT <= 2;  //26 / 9 = 2
    16'b00011010_00001010 : OUT <= 2;  //26 / 10 = 2
    16'b00011010_00001011 : OUT <= 2;  //26 / 11 = 2
    16'b00011010_00001100 : OUT <= 2;  //26 / 12 = 2
    16'b00011010_00001101 : OUT <= 2;  //26 / 13 = 2
    16'b00011010_00001110 : OUT <= 1;  //26 / 14 = 1
    16'b00011010_00001111 : OUT <= 1;  //26 / 15 = 1
    16'b00011010_00010000 : OUT <= 1;  //26 / 16 = 1
    16'b00011010_00010001 : OUT <= 1;  //26 / 17 = 1
    16'b00011010_00010010 : OUT <= 1;  //26 / 18 = 1
    16'b00011010_00010011 : OUT <= 1;  //26 / 19 = 1
    16'b00011010_00010100 : OUT <= 1;  //26 / 20 = 1
    16'b00011010_00010101 : OUT <= 1;  //26 / 21 = 1
    16'b00011010_00010110 : OUT <= 1;  //26 / 22 = 1
    16'b00011010_00010111 : OUT <= 1;  //26 / 23 = 1
    16'b00011010_00011000 : OUT <= 1;  //26 / 24 = 1
    16'b00011010_00011001 : OUT <= 1;  //26 / 25 = 1
    16'b00011010_00011010 : OUT <= 1;  //26 / 26 = 1
    16'b00011010_00011011 : OUT <= 0;  //26 / 27 = 0
    16'b00011010_00011100 : OUT <= 0;  //26 / 28 = 0
    16'b00011010_00011101 : OUT <= 0;  //26 / 29 = 0
    16'b00011010_00011110 : OUT <= 0;  //26 / 30 = 0
    16'b00011010_00011111 : OUT <= 0;  //26 / 31 = 0
    16'b00011010_00100000 : OUT <= 0;  //26 / 32 = 0
    16'b00011010_00100001 : OUT <= 0;  //26 / 33 = 0
    16'b00011010_00100010 : OUT <= 0;  //26 / 34 = 0
    16'b00011010_00100011 : OUT <= 0;  //26 / 35 = 0
    16'b00011010_00100100 : OUT <= 0;  //26 / 36 = 0
    16'b00011010_00100101 : OUT <= 0;  //26 / 37 = 0
    16'b00011010_00100110 : OUT <= 0;  //26 / 38 = 0
    16'b00011010_00100111 : OUT <= 0;  //26 / 39 = 0
    16'b00011010_00101000 : OUT <= 0;  //26 / 40 = 0
    16'b00011010_00101001 : OUT <= 0;  //26 / 41 = 0
    16'b00011010_00101010 : OUT <= 0;  //26 / 42 = 0
    16'b00011010_00101011 : OUT <= 0;  //26 / 43 = 0
    16'b00011010_00101100 : OUT <= 0;  //26 / 44 = 0
    16'b00011010_00101101 : OUT <= 0;  //26 / 45 = 0
    16'b00011010_00101110 : OUT <= 0;  //26 / 46 = 0
    16'b00011010_00101111 : OUT <= 0;  //26 / 47 = 0
    16'b00011010_00110000 : OUT <= 0;  //26 / 48 = 0
    16'b00011010_00110001 : OUT <= 0;  //26 / 49 = 0
    16'b00011010_00110010 : OUT <= 0;  //26 / 50 = 0
    16'b00011010_00110011 : OUT <= 0;  //26 / 51 = 0
    16'b00011010_00110100 : OUT <= 0;  //26 / 52 = 0
    16'b00011010_00110101 : OUT <= 0;  //26 / 53 = 0
    16'b00011010_00110110 : OUT <= 0;  //26 / 54 = 0
    16'b00011010_00110111 : OUT <= 0;  //26 / 55 = 0
    16'b00011010_00111000 : OUT <= 0;  //26 / 56 = 0
    16'b00011010_00111001 : OUT <= 0;  //26 / 57 = 0
    16'b00011010_00111010 : OUT <= 0;  //26 / 58 = 0
    16'b00011010_00111011 : OUT <= 0;  //26 / 59 = 0
    16'b00011010_00111100 : OUT <= 0;  //26 / 60 = 0
    16'b00011010_00111101 : OUT <= 0;  //26 / 61 = 0
    16'b00011010_00111110 : OUT <= 0;  //26 / 62 = 0
    16'b00011010_00111111 : OUT <= 0;  //26 / 63 = 0
    16'b00011010_01000000 : OUT <= 0;  //26 / 64 = 0
    16'b00011010_01000001 : OUT <= 0;  //26 / 65 = 0
    16'b00011010_01000010 : OUT <= 0;  //26 / 66 = 0
    16'b00011010_01000011 : OUT <= 0;  //26 / 67 = 0
    16'b00011010_01000100 : OUT <= 0;  //26 / 68 = 0
    16'b00011010_01000101 : OUT <= 0;  //26 / 69 = 0
    16'b00011010_01000110 : OUT <= 0;  //26 / 70 = 0
    16'b00011010_01000111 : OUT <= 0;  //26 / 71 = 0
    16'b00011010_01001000 : OUT <= 0;  //26 / 72 = 0
    16'b00011010_01001001 : OUT <= 0;  //26 / 73 = 0
    16'b00011010_01001010 : OUT <= 0;  //26 / 74 = 0
    16'b00011010_01001011 : OUT <= 0;  //26 / 75 = 0
    16'b00011010_01001100 : OUT <= 0;  //26 / 76 = 0
    16'b00011010_01001101 : OUT <= 0;  //26 / 77 = 0
    16'b00011010_01001110 : OUT <= 0;  //26 / 78 = 0
    16'b00011010_01001111 : OUT <= 0;  //26 / 79 = 0
    16'b00011010_01010000 : OUT <= 0;  //26 / 80 = 0
    16'b00011010_01010001 : OUT <= 0;  //26 / 81 = 0
    16'b00011010_01010010 : OUT <= 0;  //26 / 82 = 0
    16'b00011010_01010011 : OUT <= 0;  //26 / 83 = 0
    16'b00011010_01010100 : OUT <= 0;  //26 / 84 = 0
    16'b00011010_01010101 : OUT <= 0;  //26 / 85 = 0
    16'b00011010_01010110 : OUT <= 0;  //26 / 86 = 0
    16'b00011010_01010111 : OUT <= 0;  //26 / 87 = 0
    16'b00011010_01011000 : OUT <= 0;  //26 / 88 = 0
    16'b00011010_01011001 : OUT <= 0;  //26 / 89 = 0
    16'b00011010_01011010 : OUT <= 0;  //26 / 90 = 0
    16'b00011010_01011011 : OUT <= 0;  //26 / 91 = 0
    16'b00011010_01011100 : OUT <= 0;  //26 / 92 = 0
    16'b00011010_01011101 : OUT <= 0;  //26 / 93 = 0
    16'b00011010_01011110 : OUT <= 0;  //26 / 94 = 0
    16'b00011010_01011111 : OUT <= 0;  //26 / 95 = 0
    16'b00011010_01100000 : OUT <= 0;  //26 / 96 = 0
    16'b00011010_01100001 : OUT <= 0;  //26 / 97 = 0
    16'b00011010_01100010 : OUT <= 0;  //26 / 98 = 0
    16'b00011010_01100011 : OUT <= 0;  //26 / 99 = 0
    16'b00011010_01100100 : OUT <= 0;  //26 / 100 = 0
    16'b00011010_01100101 : OUT <= 0;  //26 / 101 = 0
    16'b00011010_01100110 : OUT <= 0;  //26 / 102 = 0
    16'b00011010_01100111 : OUT <= 0;  //26 / 103 = 0
    16'b00011010_01101000 : OUT <= 0;  //26 / 104 = 0
    16'b00011010_01101001 : OUT <= 0;  //26 / 105 = 0
    16'b00011010_01101010 : OUT <= 0;  //26 / 106 = 0
    16'b00011010_01101011 : OUT <= 0;  //26 / 107 = 0
    16'b00011010_01101100 : OUT <= 0;  //26 / 108 = 0
    16'b00011010_01101101 : OUT <= 0;  //26 / 109 = 0
    16'b00011010_01101110 : OUT <= 0;  //26 / 110 = 0
    16'b00011010_01101111 : OUT <= 0;  //26 / 111 = 0
    16'b00011010_01110000 : OUT <= 0;  //26 / 112 = 0
    16'b00011010_01110001 : OUT <= 0;  //26 / 113 = 0
    16'b00011010_01110010 : OUT <= 0;  //26 / 114 = 0
    16'b00011010_01110011 : OUT <= 0;  //26 / 115 = 0
    16'b00011010_01110100 : OUT <= 0;  //26 / 116 = 0
    16'b00011010_01110101 : OUT <= 0;  //26 / 117 = 0
    16'b00011010_01110110 : OUT <= 0;  //26 / 118 = 0
    16'b00011010_01110111 : OUT <= 0;  //26 / 119 = 0
    16'b00011010_01111000 : OUT <= 0;  //26 / 120 = 0
    16'b00011010_01111001 : OUT <= 0;  //26 / 121 = 0
    16'b00011010_01111010 : OUT <= 0;  //26 / 122 = 0
    16'b00011010_01111011 : OUT <= 0;  //26 / 123 = 0
    16'b00011010_01111100 : OUT <= 0;  //26 / 124 = 0
    16'b00011010_01111101 : OUT <= 0;  //26 / 125 = 0
    16'b00011010_01111110 : OUT <= 0;  //26 / 126 = 0
    16'b00011010_01111111 : OUT <= 0;  //26 / 127 = 0
    16'b00011010_10000000 : OUT <= 0;  //26 / 128 = 0
    16'b00011010_10000001 : OUT <= 0;  //26 / 129 = 0
    16'b00011010_10000010 : OUT <= 0;  //26 / 130 = 0
    16'b00011010_10000011 : OUT <= 0;  //26 / 131 = 0
    16'b00011010_10000100 : OUT <= 0;  //26 / 132 = 0
    16'b00011010_10000101 : OUT <= 0;  //26 / 133 = 0
    16'b00011010_10000110 : OUT <= 0;  //26 / 134 = 0
    16'b00011010_10000111 : OUT <= 0;  //26 / 135 = 0
    16'b00011010_10001000 : OUT <= 0;  //26 / 136 = 0
    16'b00011010_10001001 : OUT <= 0;  //26 / 137 = 0
    16'b00011010_10001010 : OUT <= 0;  //26 / 138 = 0
    16'b00011010_10001011 : OUT <= 0;  //26 / 139 = 0
    16'b00011010_10001100 : OUT <= 0;  //26 / 140 = 0
    16'b00011010_10001101 : OUT <= 0;  //26 / 141 = 0
    16'b00011010_10001110 : OUT <= 0;  //26 / 142 = 0
    16'b00011010_10001111 : OUT <= 0;  //26 / 143 = 0
    16'b00011010_10010000 : OUT <= 0;  //26 / 144 = 0
    16'b00011010_10010001 : OUT <= 0;  //26 / 145 = 0
    16'b00011010_10010010 : OUT <= 0;  //26 / 146 = 0
    16'b00011010_10010011 : OUT <= 0;  //26 / 147 = 0
    16'b00011010_10010100 : OUT <= 0;  //26 / 148 = 0
    16'b00011010_10010101 : OUT <= 0;  //26 / 149 = 0
    16'b00011010_10010110 : OUT <= 0;  //26 / 150 = 0
    16'b00011010_10010111 : OUT <= 0;  //26 / 151 = 0
    16'b00011010_10011000 : OUT <= 0;  //26 / 152 = 0
    16'b00011010_10011001 : OUT <= 0;  //26 / 153 = 0
    16'b00011010_10011010 : OUT <= 0;  //26 / 154 = 0
    16'b00011010_10011011 : OUT <= 0;  //26 / 155 = 0
    16'b00011010_10011100 : OUT <= 0;  //26 / 156 = 0
    16'b00011010_10011101 : OUT <= 0;  //26 / 157 = 0
    16'b00011010_10011110 : OUT <= 0;  //26 / 158 = 0
    16'b00011010_10011111 : OUT <= 0;  //26 / 159 = 0
    16'b00011010_10100000 : OUT <= 0;  //26 / 160 = 0
    16'b00011010_10100001 : OUT <= 0;  //26 / 161 = 0
    16'b00011010_10100010 : OUT <= 0;  //26 / 162 = 0
    16'b00011010_10100011 : OUT <= 0;  //26 / 163 = 0
    16'b00011010_10100100 : OUT <= 0;  //26 / 164 = 0
    16'b00011010_10100101 : OUT <= 0;  //26 / 165 = 0
    16'b00011010_10100110 : OUT <= 0;  //26 / 166 = 0
    16'b00011010_10100111 : OUT <= 0;  //26 / 167 = 0
    16'b00011010_10101000 : OUT <= 0;  //26 / 168 = 0
    16'b00011010_10101001 : OUT <= 0;  //26 / 169 = 0
    16'b00011010_10101010 : OUT <= 0;  //26 / 170 = 0
    16'b00011010_10101011 : OUT <= 0;  //26 / 171 = 0
    16'b00011010_10101100 : OUT <= 0;  //26 / 172 = 0
    16'b00011010_10101101 : OUT <= 0;  //26 / 173 = 0
    16'b00011010_10101110 : OUT <= 0;  //26 / 174 = 0
    16'b00011010_10101111 : OUT <= 0;  //26 / 175 = 0
    16'b00011010_10110000 : OUT <= 0;  //26 / 176 = 0
    16'b00011010_10110001 : OUT <= 0;  //26 / 177 = 0
    16'b00011010_10110010 : OUT <= 0;  //26 / 178 = 0
    16'b00011010_10110011 : OUT <= 0;  //26 / 179 = 0
    16'b00011010_10110100 : OUT <= 0;  //26 / 180 = 0
    16'b00011010_10110101 : OUT <= 0;  //26 / 181 = 0
    16'b00011010_10110110 : OUT <= 0;  //26 / 182 = 0
    16'b00011010_10110111 : OUT <= 0;  //26 / 183 = 0
    16'b00011010_10111000 : OUT <= 0;  //26 / 184 = 0
    16'b00011010_10111001 : OUT <= 0;  //26 / 185 = 0
    16'b00011010_10111010 : OUT <= 0;  //26 / 186 = 0
    16'b00011010_10111011 : OUT <= 0;  //26 / 187 = 0
    16'b00011010_10111100 : OUT <= 0;  //26 / 188 = 0
    16'b00011010_10111101 : OUT <= 0;  //26 / 189 = 0
    16'b00011010_10111110 : OUT <= 0;  //26 / 190 = 0
    16'b00011010_10111111 : OUT <= 0;  //26 / 191 = 0
    16'b00011010_11000000 : OUT <= 0;  //26 / 192 = 0
    16'b00011010_11000001 : OUT <= 0;  //26 / 193 = 0
    16'b00011010_11000010 : OUT <= 0;  //26 / 194 = 0
    16'b00011010_11000011 : OUT <= 0;  //26 / 195 = 0
    16'b00011010_11000100 : OUT <= 0;  //26 / 196 = 0
    16'b00011010_11000101 : OUT <= 0;  //26 / 197 = 0
    16'b00011010_11000110 : OUT <= 0;  //26 / 198 = 0
    16'b00011010_11000111 : OUT <= 0;  //26 / 199 = 0
    16'b00011010_11001000 : OUT <= 0;  //26 / 200 = 0
    16'b00011010_11001001 : OUT <= 0;  //26 / 201 = 0
    16'b00011010_11001010 : OUT <= 0;  //26 / 202 = 0
    16'b00011010_11001011 : OUT <= 0;  //26 / 203 = 0
    16'b00011010_11001100 : OUT <= 0;  //26 / 204 = 0
    16'b00011010_11001101 : OUT <= 0;  //26 / 205 = 0
    16'b00011010_11001110 : OUT <= 0;  //26 / 206 = 0
    16'b00011010_11001111 : OUT <= 0;  //26 / 207 = 0
    16'b00011010_11010000 : OUT <= 0;  //26 / 208 = 0
    16'b00011010_11010001 : OUT <= 0;  //26 / 209 = 0
    16'b00011010_11010010 : OUT <= 0;  //26 / 210 = 0
    16'b00011010_11010011 : OUT <= 0;  //26 / 211 = 0
    16'b00011010_11010100 : OUT <= 0;  //26 / 212 = 0
    16'b00011010_11010101 : OUT <= 0;  //26 / 213 = 0
    16'b00011010_11010110 : OUT <= 0;  //26 / 214 = 0
    16'b00011010_11010111 : OUT <= 0;  //26 / 215 = 0
    16'b00011010_11011000 : OUT <= 0;  //26 / 216 = 0
    16'b00011010_11011001 : OUT <= 0;  //26 / 217 = 0
    16'b00011010_11011010 : OUT <= 0;  //26 / 218 = 0
    16'b00011010_11011011 : OUT <= 0;  //26 / 219 = 0
    16'b00011010_11011100 : OUT <= 0;  //26 / 220 = 0
    16'b00011010_11011101 : OUT <= 0;  //26 / 221 = 0
    16'b00011010_11011110 : OUT <= 0;  //26 / 222 = 0
    16'b00011010_11011111 : OUT <= 0;  //26 / 223 = 0
    16'b00011010_11100000 : OUT <= 0;  //26 / 224 = 0
    16'b00011010_11100001 : OUT <= 0;  //26 / 225 = 0
    16'b00011010_11100010 : OUT <= 0;  //26 / 226 = 0
    16'b00011010_11100011 : OUT <= 0;  //26 / 227 = 0
    16'b00011010_11100100 : OUT <= 0;  //26 / 228 = 0
    16'b00011010_11100101 : OUT <= 0;  //26 / 229 = 0
    16'b00011010_11100110 : OUT <= 0;  //26 / 230 = 0
    16'b00011010_11100111 : OUT <= 0;  //26 / 231 = 0
    16'b00011010_11101000 : OUT <= 0;  //26 / 232 = 0
    16'b00011010_11101001 : OUT <= 0;  //26 / 233 = 0
    16'b00011010_11101010 : OUT <= 0;  //26 / 234 = 0
    16'b00011010_11101011 : OUT <= 0;  //26 / 235 = 0
    16'b00011010_11101100 : OUT <= 0;  //26 / 236 = 0
    16'b00011010_11101101 : OUT <= 0;  //26 / 237 = 0
    16'b00011010_11101110 : OUT <= 0;  //26 / 238 = 0
    16'b00011010_11101111 : OUT <= 0;  //26 / 239 = 0
    16'b00011010_11110000 : OUT <= 0;  //26 / 240 = 0
    16'b00011010_11110001 : OUT <= 0;  //26 / 241 = 0
    16'b00011010_11110010 : OUT <= 0;  //26 / 242 = 0
    16'b00011010_11110011 : OUT <= 0;  //26 / 243 = 0
    16'b00011010_11110100 : OUT <= 0;  //26 / 244 = 0
    16'b00011010_11110101 : OUT <= 0;  //26 / 245 = 0
    16'b00011010_11110110 : OUT <= 0;  //26 / 246 = 0
    16'b00011010_11110111 : OUT <= 0;  //26 / 247 = 0
    16'b00011010_11111000 : OUT <= 0;  //26 / 248 = 0
    16'b00011010_11111001 : OUT <= 0;  //26 / 249 = 0
    16'b00011010_11111010 : OUT <= 0;  //26 / 250 = 0
    16'b00011010_11111011 : OUT <= 0;  //26 / 251 = 0
    16'b00011010_11111100 : OUT <= 0;  //26 / 252 = 0
    16'b00011010_11111101 : OUT <= 0;  //26 / 253 = 0
    16'b00011010_11111110 : OUT <= 0;  //26 / 254 = 0
    16'b00011010_11111111 : OUT <= 0;  //26 / 255 = 0
    16'b00011011_00000000 : OUT <= 0;  //27 / 0 = 0
    16'b00011011_00000001 : OUT <= 27;  //27 / 1 = 27
    16'b00011011_00000010 : OUT <= 13;  //27 / 2 = 13
    16'b00011011_00000011 : OUT <= 9;  //27 / 3 = 9
    16'b00011011_00000100 : OUT <= 6;  //27 / 4 = 6
    16'b00011011_00000101 : OUT <= 5;  //27 / 5 = 5
    16'b00011011_00000110 : OUT <= 4;  //27 / 6 = 4
    16'b00011011_00000111 : OUT <= 3;  //27 / 7 = 3
    16'b00011011_00001000 : OUT <= 3;  //27 / 8 = 3
    16'b00011011_00001001 : OUT <= 3;  //27 / 9 = 3
    16'b00011011_00001010 : OUT <= 2;  //27 / 10 = 2
    16'b00011011_00001011 : OUT <= 2;  //27 / 11 = 2
    16'b00011011_00001100 : OUT <= 2;  //27 / 12 = 2
    16'b00011011_00001101 : OUT <= 2;  //27 / 13 = 2
    16'b00011011_00001110 : OUT <= 1;  //27 / 14 = 1
    16'b00011011_00001111 : OUT <= 1;  //27 / 15 = 1
    16'b00011011_00010000 : OUT <= 1;  //27 / 16 = 1
    16'b00011011_00010001 : OUT <= 1;  //27 / 17 = 1
    16'b00011011_00010010 : OUT <= 1;  //27 / 18 = 1
    16'b00011011_00010011 : OUT <= 1;  //27 / 19 = 1
    16'b00011011_00010100 : OUT <= 1;  //27 / 20 = 1
    16'b00011011_00010101 : OUT <= 1;  //27 / 21 = 1
    16'b00011011_00010110 : OUT <= 1;  //27 / 22 = 1
    16'b00011011_00010111 : OUT <= 1;  //27 / 23 = 1
    16'b00011011_00011000 : OUT <= 1;  //27 / 24 = 1
    16'b00011011_00011001 : OUT <= 1;  //27 / 25 = 1
    16'b00011011_00011010 : OUT <= 1;  //27 / 26 = 1
    16'b00011011_00011011 : OUT <= 1;  //27 / 27 = 1
    16'b00011011_00011100 : OUT <= 0;  //27 / 28 = 0
    16'b00011011_00011101 : OUT <= 0;  //27 / 29 = 0
    16'b00011011_00011110 : OUT <= 0;  //27 / 30 = 0
    16'b00011011_00011111 : OUT <= 0;  //27 / 31 = 0
    16'b00011011_00100000 : OUT <= 0;  //27 / 32 = 0
    16'b00011011_00100001 : OUT <= 0;  //27 / 33 = 0
    16'b00011011_00100010 : OUT <= 0;  //27 / 34 = 0
    16'b00011011_00100011 : OUT <= 0;  //27 / 35 = 0
    16'b00011011_00100100 : OUT <= 0;  //27 / 36 = 0
    16'b00011011_00100101 : OUT <= 0;  //27 / 37 = 0
    16'b00011011_00100110 : OUT <= 0;  //27 / 38 = 0
    16'b00011011_00100111 : OUT <= 0;  //27 / 39 = 0
    16'b00011011_00101000 : OUT <= 0;  //27 / 40 = 0
    16'b00011011_00101001 : OUT <= 0;  //27 / 41 = 0
    16'b00011011_00101010 : OUT <= 0;  //27 / 42 = 0
    16'b00011011_00101011 : OUT <= 0;  //27 / 43 = 0
    16'b00011011_00101100 : OUT <= 0;  //27 / 44 = 0
    16'b00011011_00101101 : OUT <= 0;  //27 / 45 = 0
    16'b00011011_00101110 : OUT <= 0;  //27 / 46 = 0
    16'b00011011_00101111 : OUT <= 0;  //27 / 47 = 0
    16'b00011011_00110000 : OUT <= 0;  //27 / 48 = 0
    16'b00011011_00110001 : OUT <= 0;  //27 / 49 = 0
    16'b00011011_00110010 : OUT <= 0;  //27 / 50 = 0
    16'b00011011_00110011 : OUT <= 0;  //27 / 51 = 0
    16'b00011011_00110100 : OUT <= 0;  //27 / 52 = 0
    16'b00011011_00110101 : OUT <= 0;  //27 / 53 = 0
    16'b00011011_00110110 : OUT <= 0;  //27 / 54 = 0
    16'b00011011_00110111 : OUT <= 0;  //27 / 55 = 0
    16'b00011011_00111000 : OUT <= 0;  //27 / 56 = 0
    16'b00011011_00111001 : OUT <= 0;  //27 / 57 = 0
    16'b00011011_00111010 : OUT <= 0;  //27 / 58 = 0
    16'b00011011_00111011 : OUT <= 0;  //27 / 59 = 0
    16'b00011011_00111100 : OUT <= 0;  //27 / 60 = 0
    16'b00011011_00111101 : OUT <= 0;  //27 / 61 = 0
    16'b00011011_00111110 : OUT <= 0;  //27 / 62 = 0
    16'b00011011_00111111 : OUT <= 0;  //27 / 63 = 0
    16'b00011011_01000000 : OUT <= 0;  //27 / 64 = 0
    16'b00011011_01000001 : OUT <= 0;  //27 / 65 = 0
    16'b00011011_01000010 : OUT <= 0;  //27 / 66 = 0
    16'b00011011_01000011 : OUT <= 0;  //27 / 67 = 0
    16'b00011011_01000100 : OUT <= 0;  //27 / 68 = 0
    16'b00011011_01000101 : OUT <= 0;  //27 / 69 = 0
    16'b00011011_01000110 : OUT <= 0;  //27 / 70 = 0
    16'b00011011_01000111 : OUT <= 0;  //27 / 71 = 0
    16'b00011011_01001000 : OUT <= 0;  //27 / 72 = 0
    16'b00011011_01001001 : OUT <= 0;  //27 / 73 = 0
    16'b00011011_01001010 : OUT <= 0;  //27 / 74 = 0
    16'b00011011_01001011 : OUT <= 0;  //27 / 75 = 0
    16'b00011011_01001100 : OUT <= 0;  //27 / 76 = 0
    16'b00011011_01001101 : OUT <= 0;  //27 / 77 = 0
    16'b00011011_01001110 : OUT <= 0;  //27 / 78 = 0
    16'b00011011_01001111 : OUT <= 0;  //27 / 79 = 0
    16'b00011011_01010000 : OUT <= 0;  //27 / 80 = 0
    16'b00011011_01010001 : OUT <= 0;  //27 / 81 = 0
    16'b00011011_01010010 : OUT <= 0;  //27 / 82 = 0
    16'b00011011_01010011 : OUT <= 0;  //27 / 83 = 0
    16'b00011011_01010100 : OUT <= 0;  //27 / 84 = 0
    16'b00011011_01010101 : OUT <= 0;  //27 / 85 = 0
    16'b00011011_01010110 : OUT <= 0;  //27 / 86 = 0
    16'b00011011_01010111 : OUT <= 0;  //27 / 87 = 0
    16'b00011011_01011000 : OUT <= 0;  //27 / 88 = 0
    16'b00011011_01011001 : OUT <= 0;  //27 / 89 = 0
    16'b00011011_01011010 : OUT <= 0;  //27 / 90 = 0
    16'b00011011_01011011 : OUT <= 0;  //27 / 91 = 0
    16'b00011011_01011100 : OUT <= 0;  //27 / 92 = 0
    16'b00011011_01011101 : OUT <= 0;  //27 / 93 = 0
    16'b00011011_01011110 : OUT <= 0;  //27 / 94 = 0
    16'b00011011_01011111 : OUT <= 0;  //27 / 95 = 0
    16'b00011011_01100000 : OUT <= 0;  //27 / 96 = 0
    16'b00011011_01100001 : OUT <= 0;  //27 / 97 = 0
    16'b00011011_01100010 : OUT <= 0;  //27 / 98 = 0
    16'b00011011_01100011 : OUT <= 0;  //27 / 99 = 0
    16'b00011011_01100100 : OUT <= 0;  //27 / 100 = 0
    16'b00011011_01100101 : OUT <= 0;  //27 / 101 = 0
    16'b00011011_01100110 : OUT <= 0;  //27 / 102 = 0
    16'b00011011_01100111 : OUT <= 0;  //27 / 103 = 0
    16'b00011011_01101000 : OUT <= 0;  //27 / 104 = 0
    16'b00011011_01101001 : OUT <= 0;  //27 / 105 = 0
    16'b00011011_01101010 : OUT <= 0;  //27 / 106 = 0
    16'b00011011_01101011 : OUT <= 0;  //27 / 107 = 0
    16'b00011011_01101100 : OUT <= 0;  //27 / 108 = 0
    16'b00011011_01101101 : OUT <= 0;  //27 / 109 = 0
    16'b00011011_01101110 : OUT <= 0;  //27 / 110 = 0
    16'b00011011_01101111 : OUT <= 0;  //27 / 111 = 0
    16'b00011011_01110000 : OUT <= 0;  //27 / 112 = 0
    16'b00011011_01110001 : OUT <= 0;  //27 / 113 = 0
    16'b00011011_01110010 : OUT <= 0;  //27 / 114 = 0
    16'b00011011_01110011 : OUT <= 0;  //27 / 115 = 0
    16'b00011011_01110100 : OUT <= 0;  //27 / 116 = 0
    16'b00011011_01110101 : OUT <= 0;  //27 / 117 = 0
    16'b00011011_01110110 : OUT <= 0;  //27 / 118 = 0
    16'b00011011_01110111 : OUT <= 0;  //27 / 119 = 0
    16'b00011011_01111000 : OUT <= 0;  //27 / 120 = 0
    16'b00011011_01111001 : OUT <= 0;  //27 / 121 = 0
    16'b00011011_01111010 : OUT <= 0;  //27 / 122 = 0
    16'b00011011_01111011 : OUT <= 0;  //27 / 123 = 0
    16'b00011011_01111100 : OUT <= 0;  //27 / 124 = 0
    16'b00011011_01111101 : OUT <= 0;  //27 / 125 = 0
    16'b00011011_01111110 : OUT <= 0;  //27 / 126 = 0
    16'b00011011_01111111 : OUT <= 0;  //27 / 127 = 0
    16'b00011011_10000000 : OUT <= 0;  //27 / 128 = 0
    16'b00011011_10000001 : OUT <= 0;  //27 / 129 = 0
    16'b00011011_10000010 : OUT <= 0;  //27 / 130 = 0
    16'b00011011_10000011 : OUT <= 0;  //27 / 131 = 0
    16'b00011011_10000100 : OUT <= 0;  //27 / 132 = 0
    16'b00011011_10000101 : OUT <= 0;  //27 / 133 = 0
    16'b00011011_10000110 : OUT <= 0;  //27 / 134 = 0
    16'b00011011_10000111 : OUT <= 0;  //27 / 135 = 0
    16'b00011011_10001000 : OUT <= 0;  //27 / 136 = 0
    16'b00011011_10001001 : OUT <= 0;  //27 / 137 = 0
    16'b00011011_10001010 : OUT <= 0;  //27 / 138 = 0
    16'b00011011_10001011 : OUT <= 0;  //27 / 139 = 0
    16'b00011011_10001100 : OUT <= 0;  //27 / 140 = 0
    16'b00011011_10001101 : OUT <= 0;  //27 / 141 = 0
    16'b00011011_10001110 : OUT <= 0;  //27 / 142 = 0
    16'b00011011_10001111 : OUT <= 0;  //27 / 143 = 0
    16'b00011011_10010000 : OUT <= 0;  //27 / 144 = 0
    16'b00011011_10010001 : OUT <= 0;  //27 / 145 = 0
    16'b00011011_10010010 : OUT <= 0;  //27 / 146 = 0
    16'b00011011_10010011 : OUT <= 0;  //27 / 147 = 0
    16'b00011011_10010100 : OUT <= 0;  //27 / 148 = 0
    16'b00011011_10010101 : OUT <= 0;  //27 / 149 = 0
    16'b00011011_10010110 : OUT <= 0;  //27 / 150 = 0
    16'b00011011_10010111 : OUT <= 0;  //27 / 151 = 0
    16'b00011011_10011000 : OUT <= 0;  //27 / 152 = 0
    16'b00011011_10011001 : OUT <= 0;  //27 / 153 = 0
    16'b00011011_10011010 : OUT <= 0;  //27 / 154 = 0
    16'b00011011_10011011 : OUT <= 0;  //27 / 155 = 0
    16'b00011011_10011100 : OUT <= 0;  //27 / 156 = 0
    16'b00011011_10011101 : OUT <= 0;  //27 / 157 = 0
    16'b00011011_10011110 : OUT <= 0;  //27 / 158 = 0
    16'b00011011_10011111 : OUT <= 0;  //27 / 159 = 0
    16'b00011011_10100000 : OUT <= 0;  //27 / 160 = 0
    16'b00011011_10100001 : OUT <= 0;  //27 / 161 = 0
    16'b00011011_10100010 : OUT <= 0;  //27 / 162 = 0
    16'b00011011_10100011 : OUT <= 0;  //27 / 163 = 0
    16'b00011011_10100100 : OUT <= 0;  //27 / 164 = 0
    16'b00011011_10100101 : OUT <= 0;  //27 / 165 = 0
    16'b00011011_10100110 : OUT <= 0;  //27 / 166 = 0
    16'b00011011_10100111 : OUT <= 0;  //27 / 167 = 0
    16'b00011011_10101000 : OUT <= 0;  //27 / 168 = 0
    16'b00011011_10101001 : OUT <= 0;  //27 / 169 = 0
    16'b00011011_10101010 : OUT <= 0;  //27 / 170 = 0
    16'b00011011_10101011 : OUT <= 0;  //27 / 171 = 0
    16'b00011011_10101100 : OUT <= 0;  //27 / 172 = 0
    16'b00011011_10101101 : OUT <= 0;  //27 / 173 = 0
    16'b00011011_10101110 : OUT <= 0;  //27 / 174 = 0
    16'b00011011_10101111 : OUT <= 0;  //27 / 175 = 0
    16'b00011011_10110000 : OUT <= 0;  //27 / 176 = 0
    16'b00011011_10110001 : OUT <= 0;  //27 / 177 = 0
    16'b00011011_10110010 : OUT <= 0;  //27 / 178 = 0
    16'b00011011_10110011 : OUT <= 0;  //27 / 179 = 0
    16'b00011011_10110100 : OUT <= 0;  //27 / 180 = 0
    16'b00011011_10110101 : OUT <= 0;  //27 / 181 = 0
    16'b00011011_10110110 : OUT <= 0;  //27 / 182 = 0
    16'b00011011_10110111 : OUT <= 0;  //27 / 183 = 0
    16'b00011011_10111000 : OUT <= 0;  //27 / 184 = 0
    16'b00011011_10111001 : OUT <= 0;  //27 / 185 = 0
    16'b00011011_10111010 : OUT <= 0;  //27 / 186 = 0
    16'b00011011_10111011 : OUT <= 0;  //27 / 187 = 0
    16'b00011011_10111100 : OUT <= 0;  //27 / 188 = 0
    16'b00011011_10111101 : OUT <= 0;  //27 / 189 = 0
    16'b00011011_10111110 : OUT <= 0;  //27 / 190 = 0
    16'b00011011_10111111 : OUT <= 0;  //27 / 191 = 0
    16'b00011011_11000000 : OUT <= 0;  //27 / 192 = 0
    16'b00011011_11000001 : OUT <= 0;  //27 / 193 = 0
    16'b00011011_11000010 : OUT <= 0;  //27 / 194 = 0
    16'b00011011_11000011 : OUT <= 0;  //27 / 195 = 0
    16'b00011011_11000100 : OUT <= 0;  //27 / 196 = 0
    16'b00011011_11000101 : OUT <= 0;  //27 / 197 = 0
    16'b00011011_11000110 : OUT <= 0;  //27 / 198 = 0
    16'b00011011_11000111 : OUT <= 0;  //27 / 199 = 0
    16'b00011011_11001000 : OUT <= 0;  //27 / 200 = 0
    16'b00011011_11001001 : OUT <= 0;  //27 / 201 = 0
    16'b00011011_11001010 : OUT <= 0;  //27 / 202 = 0
    16'b00011011_11001011 : OUT <= 0;  //27 / 203 = 0
    16'b00011011_11001100 : OUT <= 0;  //27 / 204 = 0
    16'b00011011_11001101 : OUT <= 0;  //27 / 205 = 0
    16'b00011011_11001110 : OUT <= 0;  //27 / 206 = 0
    16'b00011011_11001111 : OUT <= 0;  //27 / 207 = 0
    16'b00011011_11010000 : OUT <= 0;  //27 / 208 = 0
    16'b00011011_11010001 : OUT <= 0;  //27 / 209 = 0
    16'b00011011_11010010 : OUT <= 0;  //27 / 210 = 0
    16'b00011011_11010011 : OUT <= 0;  //27 / 211 = 0
    16'b00011011_11010100 : OUT <= 0;  //27 / 212 = 0
    16'b00011011_11010101 : OUT <= 0;  //27 / 213 = 0
    16'b00011011_11010110 : OUT <= 0;  //27 / 214 = 0
    16'b00011011_11010111 : OUT <= 0;  //27 / 215 = 0
    16'b00011011_11011000 : OUT <= 0;  //27 / 216 = 0
    16'b00011011_11011001 : OUT <= 0;  //27 / 217 = 0
    16'b00011011_11011010 : OUT <= 0;  //27 / 218 = 0
    16'b00011011_11011011 : OUT <= 0;  //27 / 219 = 0
    16'b00011011_11011100 : OUT <= 0;  //27 / 220 = 0
    16'b00011011_11011101 : OUT <= 0;  //27 / 221 = 0
    16'b00011011_11011110 : OUT <= 0;  //27 / 222 = 0
    16'b00011011_11011111 : OUT <= 0;  //27 / 223 = 0
    16'b00011011_11100000 : OUT <= 0;  //27 / 224 = 0
    16'b00011011_11100001 : OUT <= 0;  //27 / 225 = 0
    16'b00011011_11100010 : OUT <= 0;  //27 / 226 = 0
    16'b00011011_11100011 : OUT <= 0;  //27 / 227 = 0
    16'b00011011_11100100 : OUT <= 0;  //27 / 228 = 0
    16'b00011011_11100101 : OUT <= 0;  //27 / 229 = 0
    16'b00011011_11100110 : OUT <= 0;  //27 / 230 = 0
    16'b00011011_11100111 : OUT <= 0;  //27 / 231 = 0
    16'b00011011_11101000 : OUT <= 0;  //27 / 232 = 0
    16'b00011011_11101001 : OUT <= 0;  //27 / 233 = 0
    16'b00011011_11101010 : OUT <= 0;  //27 / 234 = 0
    16'b00011011_11101011 : OUT <= 0;  //27 / 235 = 0
    16'b00011011_11101100 : OUT <= 0;  //27 / 236 = 0
    16'b00011011_11101101 : OUT <= 0;  //27 / 237 = 0
    16'b00011011_11101110 : OUT <= 0;  //27 / 238 = 0
    16'b00011011_11101111 : OUT <= 0;  //27 / 239 = 0
    16'b00011011_11110000 : OUT <= 0;  //27 / 240 = 0
    16'b00011011_11110001 : OUT <= 0;  //27 / 241 = 0
    16'b00011011_11110010 : OUT <= 0;  //27 / 242 = 0
    16'b00011011_11110011 : OUT <= 0;  //27 / 243 = 0
    16'b00011011_11110100 : OUT <= 0;  //27 / 244 = 0
    16'b00011011_11110101 : OUT <= 0;  //27 / 245 = 0
    16'b00011011_11110110 : OUT <= 0;  //27 / 246 = 0
    16'b00011011_11110111 : OUT <= 0;  //27 / 247 = 0
    16'b00011011_11111000 : OUT <= 0;  //27 / 248 = 0
    16'b00011011_11111001 : OUT <= 0;  //27 / 249 = 0
    16'b00011011_11111010 : OUT <= 0;  //27 / 250 = 0
    16'b00011011_11111011 : OUT <= 0;  //27 / 251 = 0
    16'b00011011_11111100 : OUT <= 0;  //27 / 252 = 0
    16'b00011011_11111101 : OUT <= 0;  //27 / 253 = 0
    16'b00011011_11111110 : OUT <= 0;  //27 / 254 = 0
    16'b00011011_11111111 : OUT <= 0;  //27 / 255 = 0
    16'b00011100_00000000 : OUT <= 0;  //28 / 0 = 0
    16'b00011100_00000001 : OUT <= 28;  //28 / 1 = 28
    16'b00011100_00000010 : OUT <= 14;  //28 / 2 = 14
    16'b00011100_00000011 : OUT <= 9;  //28 / 3 = 9
    16'b00011100_00000100 : OUT <= 7;  //28 / 4 = 7
    16'b00011100_00000101 : OUT <= 5;  //28 / 5 = 5
    16'b00011100_00000110 : OUT <= 4;  //28 / 6 = 4
    16'b00011100_00000111 : OUT <= 4;  //28 / 7 = 4
    16'b00011100_00001000 : OUT <= 3;  //28 / 8 = 3
    16'b00011100_00001001 : OUT <= 3;  //28 / 9 = 3
    16'b00011100_00001010 : OUT <= 2;  //28 / 10 = 2
    16'b00011100_00001011 : OUT <= 2;  //28 / 11 = 2
    16'b00011100_00001100 : OUT <= 2;  //28 / 12 = 2
    16'b00011100_00001101 : OUT <= 2;  //28 / 13 = 2
    16'b00011100_00001110 : OUT <= 2;  //28 / 14 = 2
    16'b00011100_00001111 : OUT <= 1;  //28 / 15 = 1
    16'b00011100_00010000 : OUT <= 1;  //28 / 16 = 1
    16'b00011100_00010001 : OUT <= 1;  //28 / 17 = 1
    16'b00011100_00010010 : OUT <= 1;  //28 / 18 = 1
    16'b00011100_00010011 : OUT <= 1;  //28 / 19 = 1
    16'b00011100_00010100 : OUT <= 1;  //28 / 20 = 1
    16'b00011100_00010101 : OUT <= 1;  //28 / 21 = 1
    16'b00011100_00010110 : OUT <= 1;  //28 / 22 = 1
    16'b00011100_00010111 : OUT <= 1;  //28 / 23 = 1
    16'b00011100_00011000 : OUT <= 1;  //28 / 24 = 1
    16'b00011100_00011001 : OUT <= 1;  //28 / 25 = 1
    16'b00011100_00011010 : OUT <= 1;  //28 / 26 = 1
    16'b00011100_00011011 : OUT <= 1;  //28 / 27 = 1
    16'b00011100_00011100 : OUT <= 1;  //28 / 28 = 1
    16'b00011100_00011101 : OUT <= 0;  //28 / 29 = 0
    16'b00011100_00011110 : OUT <= 0;  //28 / 30 = 0
    16'b00011100_00011111 : OUT <= 0;  //28 / 31 = 0
    16'b00011100_00100000 : OUT <= 0;  //28 / 32 = 0
    16'b00011100_00100001 : OUT <= 0;  //28 / 33 = 0
    16'b00011100_00100010 : OUT <= 0;  //28 / 34 = 0
    16'b00011100_00100011 : OUT <= 0;  //28 / 35 = 0
    16'b00011100_00100100 : OUT <= 0;  //28 / 36 = 0
    16'b00011100_00100101 : OUT <= 0;  //28 / 37 = 0
    16'b00011100_00100110 : OUT <= 0;  //28 / 38 = 0
    16'b00011100_00100111 : OUT <= 0;  //28 / 39 = 0
    16'b00011100_00101000 : OUT <= 0;  //28 / 40 = 0
    16'b00011100_00101001 : OUT <= 0;  //28 / 41 = 0
    16'b00011100_00101010 : OUT <= 0;  //28 / 42 = 0
    16'b00011100_00101011 : OUT <= 0;  //28 / 43 = 0
    16'b00011100_00101100 : OUT <= 0;  //28 / 44 = 0
    16'b00011100_00101101 : OUT <= 0;  //28 / 45 = 0
    16'b00011100_00101110 : OUT <= 0;  //28 / 46 = 0
    16'b00011100_00101111 : OUT <= 0;  //28 / 47 = 0
    16'b00011100_00110000 : OUT <= 0;  //28 / 48 = 0
    16'b00011100_00110001 : OUT <= 0;  //28 / 49 = 0
    16'b00011100_00110010 : OUT <= 0;  //28 / 50 = 0
    16'b00011100_00110011 : OUT <= 0;  //28 / 51 = 0
    16'b00011100_00110100 : OUT <= 0;  //28 / 52 = 0
    16'b00011100_00110101 : OUT <= 0;  //28 / 53 = 0
    16'b00011100_00110110 : OUT <= 0;  //28 / 54 = 0
    16'b00011100_00110111 : OUT <= 0;  //28 / 55 = 0
    16'b00011100_00111000 : OUT <= 0;  //28 / 56 = 0
    16'b00011100_00111001 : OUT <= 0;  //28 / 57 = 0
    16'b00011100_00111010 : OUT <= 0;  //28 / 58 = 0
    16'b00011100_00111011 : OUT <= 0;  //28 / 59 = 0
    16'b00011100_00111100 : OUT <= 0;  //28 / 60 = 0
    16'b00011100_00111101 : OUT <= 0;  //28 / 61 = 0
    16'b00011100_00111110 : OUT <= 0;  //28 / 62 = 0
    16'b00011100_00111111 : OUT <= 0;  //28 / 63 = 0
    16'b00011100_01000000 : OUT <= 0;  //28 / 64 = 0
    16'b00011100_01000001 : OUT <= 0;  //28 / 65 = 0
    16'b00011100_01000010 : OUT <= 0;  //28 / 66 = 0
    16'b00011100_01000011 : OUT <= 0;  //28 / 67 = 0
    16'b00011100_01000100 : OUT <= 0;  //28 / 68 = 0
    16'b00011100_01000101 : OUT <= 0;  //28 / 69 = 0
    16'b00011100_01000110 : OUT <= 0;  //28 / 70 = 0
    16'b00011100_01000111 : OUT <= 0;  //28 / 71 = 0
    16'b00011100_01001000 : OUT <= 0;  //28 / 72 = 0
    16'b00011100_01001001 : OUT <= 0;  //28 / 73 = 0
    16'b00011100_01001010 : OUT <= 0;  //28 / 74 = 0
    16'b00011100_01001011 : OUT <= 0;  //28 / 75 = 0
    16'b00011100_01001100 : OUT <= 0;  //28 / 76 = 0
    16'b00011100_01001101 : OUT <= 0;  //28 / 77 = 0
    16'b00011100_01001110 : OUT <= 0;  //28 / 78 = 0
    16'b00011100_01001111 : OUT <= 0;  //28 / 79 = 0
    16'b00011100_01010000 : OUT <= 0;  //28 / 80 = 0
    16'b00011100_01010001 : OUT <= 0;  //28 / 81 = 0
    16'b00011100_01010010 : OUT <= 0;  //28 / 82 = 0
    16'b00011100_01010011 : OUT <= 0;  //28 / 83 = 0
    16'b00011100_01010100 : OUT <= 0;  //28 / 84 = 0
    16'b00011100_01010101 : OUT <= 0;  //28 / 85 = 0
    16'b00011100_01010110 : OUT <= 0;  //28 / 86 = 0
    16'b00011100_01010111 : OUT <= 0;  //28 / 87 = 0
    16'b00011100_01011000 : OUT <= 0;  //28 / 88 = 0
    16'b00011100_01011001 : OUT <= 0;  //28 / 89 = 0
    16'b00011100_01011010 : OUT <= 0;  //28 / 90 = 0
    16'b00011100_01011011 : OUT <= 0;  //28 / 91 = 0
    16'b00011100_01011100 : OUT <= 0;  //28 / 92 = 0
    16'b00011100_01011101 : OUT <= 0;  //28 / 93 = 0
    16'b00011100_01011110 : OUT <= 0;  //28 / 94 = 0
    16'b00011100_01011111 : OUT <= 0;  //28 / 95 = 0
    16'b00011100_01100000 : OUT <= 0;  //28 / 96 = 0
    16'b00011100_01100001 : OUT <= 0;  //28 / 97 = 0
    16'b00011100_01100010 : OUT <= 0;  //28 / 98 = 0
    16'b00011100_01100011 : OUT <= 0;  //28 / 99 = 0
    16'b00011100_01100100 : OUT <= 0;  //28 / 100 = 0
    16'b00011100_01100101 : OUT <= 0;  //28 / 101 = 0
    16'b00011100_01100110 : OUT <= 0;  //28 / 102 = 0
    16'b00011100_01100111 : OUT <= 0;  //28 / 103 = 0
    16'b00011100_01101000 : OUT <= 0;  //28 / 104 = 0
    16'b00011100_01101001 : OUT <= 0;  //28 / 105 = 0
    16'b00011100_01101010 : OUT <= 0;  //28 / 106 = 0
    16'b00011100_01101011 : OUT <= 0;  //28 / 107 = 0
    16'b00011100_01101100 : OUT <= 0;  //28 / 108 = 0
    16'b00011100_01101101 : OUT <= 0;  //28 / 109 = 0
    16'b00011100_01101110 : OUT <= 0;  //28 / 110 = 0
    16'b00011100_01101111 : OUT <= 0;  //28 / 111 = 0
    16'b00011100_01110000 : OUT <= 0;  //28 / 112 = 0
    16'b00011100_01110001 : OUT <= 0;  //28 / 113 = 0
    16'b00011100_01110010 : OUT <= 0;  //28 / 114 = 0
    16'b00011100_01110011 : OUT <= 0;  //28 / 115 = 0
    16'b00011100_01110100 : OUT <= 0;  //28 / 116 = 0
    16'b00011100_01110101 : OUT <= 0;  //28 / 117 = 0
    16'b00011100_01110110 : OUT <= 0;  //28 / 118 = 0
    16'b00011100_01110111 : OUT <= 0;  //28 / 119 = 0
    16'b00011100_01111000 : OUT <= 0;  //28 / 120 = 0
    16'b00011100_01111001 : OUT <= 0;  //28 / 121 = 0
    16'b00011100_01111010 : OUT <= 0;  //28 / 122 = 0
    16'b00011100_01111011 : OUT <= 0;  //28 / 123 = 0
    16'b00011100_01111100 : OUT <= 0;  //28 / 124 = 0
    16'b00011100_01111101 : OUT <= 0;  //28 / 125 = 0
    16'b00011100_01111110 : OUT <= 0;  //28 / 126 = 0
    16'b00011100_01111111 : OUT <= 0;  //28 / 127 = 0
    16'b00011100_10000000 : OUT <= 0;  //28 / 128 = 0
    16'b00011100_10000001 : OUT <= 0;  //28 / 129 = 0
    16'b00011100_10000010 : OUT <= 0;  //28 / 130 = 0
    16'b00011100_10000011 : OUT <= 0;  //28 / 131 = 0
    16'b00011100_10000100 : OUT <= 0;  //28 / 132 = 0
    16'b00011100_10000101 : OUT <= 0;  //28 / 133 = 0
    16'b00011100_10000110 : OUT <= 0;  //28 / 134 = 0
    16'b00011100_10000111 : OUT <= 0;  //28 / 135 = 0
    16'b00011100_10001000 : OUT <= 0;  //28 / 136 = 0
    16'b00011100_10001001 : OUT <= 0;  //28 / 137 = 0
    16'b00011100_10001010 : OUT <= 0;  //28 / 138 = 0
    16'b00011100_10001011 : OUT <= 0;  //28 / 139 = 0
    16'b00011100_10001100 : OUT <= 0;  //28 / 140 = 0
    16'b00011100_10001101 : OUT <= 0;  //28 / 141 = 0
    16'b00011100_10001110 : OUT <= 0;  //28 / 142 = 0
    16'b00011100_10001111 : OUT <= 0;  //28 / 143 = 0
    16'b00011100_10010000 : OUT <= 0;  //28 / 144 = 0
    16'b00011100_10010001 : OUT <= 0;  //28 / 145 = 0
    16'b00011100_10010010 : OUT <= 0;  //28 / 146 = 0
    16'b00011100_10010011 : OUT <= 0;  //28 / 147 = 0
    16'b00011100_10010100 : OUT <= 0;  //28 / 148 = 0
    16'b00011100_10010101 : OUT <= 0;  //28 / 149 = 0
    16'b00011100_10010110 : OUT <= 0;  //28 / 150 = 0
    16'b00011100_10010111 : OUT <= 0;  //28 / 151 = 0
    16'b00011100_10011000 : OUT <= 0;  //28 / 152 = 0
    16'b00011100_10011001 : OUT <= 0;  //28 / 153 = 0
    16'b00011100_10011010 : OUT <= 0;  //28 / 154 = 0
    16'b00011100_10011011 : OUT <= 0;  //28 / 155 = 0
    16'b00011100_10011100 : OUT <= 0;  //28 / 156 = 0
    16'b00011100_10011101 : OUT <= 0;  //28 / 157 = 0
    16'b00011100_10011110 : OUT <= 0;  //28 / 158 = 0
    16'b00011100_10011111 : OUT <= 0;  //28 / 159 = 0
    16'b00011100_10100000 : OUT <= 0;  //28 / 160 = 0
    16'b00011100_10100001 : OUT <= 0;  //28 / 161 = 0
    16'b00011100_10100010 : OUT <= 0;  //28 / 162 = 0
    16'b00011100_10100011 : OUT <= 0;  //28 / 163 = 0
    16'b00011100_10100100 : OUT <= 0;  //28 / 164 = 0
    16'b00011100_10100101 : OUT <= 0;  //28 / 165 = 0
    16'b00011100_10100110 : OUT <= 0;  //28 / 166 = 0
    16'b00011100_10100111 : OUT <= 0;  //28 / 167 = 0
    16'b00011100_10101000 : OUT <= 0;  //28 / 168 = 0
    16'b00011100_10101001 : OUT <= 0;  //28 / 169 = 0
    16'b00011100_10101010 : OUT <= 0;  //28 / 170 = 0
    16'b00011100_10101011 : OUT <= 0;  //28 / 171 = 0
    16'b00011100_10101100 : OUT <= 0;  //28 / 172 = 0
    16'b00011100_10101101 : OUT <= 0;  //28 / 173 = 0
    16'b00011100_10101110 : OUT <= 0;  //28 / 174 = 0
    16'b00011100_10101111 : OUT <= 0;  //28 / 175 = 0
    16'b00011100_10110000 : OUT <= 0;  //28 / 176 = 0
    16'b00011100_10110001 : OUT <= 0;  //28 / 177 = 0
    16'b00011100_10110010 : OUT <= 0;  //28 / 178 = 0
    16'b00011100_10110011 : OUT <= 0;  //28 / 179 = 0
    16'b00011100_10110100 : OUT <= 0;  //28 / 180 = 0
    16'b00011100_10110101 : OUT <= 0;  //28 / 181 = 0
    16'b00011100_10110110 : OUT <= 0;  //28 / 182 = 0
    16'b00011100_10110111 : OUT <= 0;  //28 / 183 = 0
    16'b00011100_10111000 : OUT <= 0;  //28 / 184 = 0
    16'b00011100_10111001 : OUT <= 0;  //28 / 185 = 0
    16'b00011100_10111010 : OUT <= 0;  //28 / 186 = 0
    16'b00011100_10111011 : OUT <= 0;  //28 / 187 = 0
    16'b00011100_10111100 : OUT <= 0;  //28 / 188 = 0
    16'b00011100_10111101 : OUT <= 0;  //28 / 189 = 0
    16'b00011100_10111110 : OUT <= 0;  //28 / 190 = 0
    16'b00011100_10111111 : OUT <= 0;  //28 / 191 = 0
    16'b00011100_11000000 : OUT <= 0;  //28 / 192 = 0
    16'b00011100_11000001 : OUT <= 0;  //28 / 193 = 0
    16'b00011100_11000010 : OUT <= 0;  //28 / 194 = 0
    16'b00011100_11000011 : OUT <= 0;  //28 / 195 = 0
    16'b00011100_11000100 : OUT <= 0;  //28 / 196 = 0
    16'b00011100_11000101 : OUT <= 0;  //28 / 197 = 0
    16'b00011100_11000110 : OUT <= 0;  //28 / 198 = 0
    16'b00011100_11000111 : OUT <= 0;  //28 / 199 = 0
    16'b00011100_11001000 : OUT <= 0;  //28 / 200 = 0
    16'b00011100_11001001 : OUT <= 0;  //28 / 201 = 0
    16'b00011100_11001010 : OUT <= 0;  //28 / 202 = 0
    16'b00011100_11001011 : OUT <= 0;  //28 / 203 = 0
    16'b00011100_11001100 : OUT <= 0;  //28 / 204 = 0
    16'b00011100_11001101 : OUT <= 0;  //28 / 205 = 0
    16'b00011100_11001110 : OUT <= 0;  //28 / 206 = 0
    16'b00011100_11001111 : OUT <= 0;  //28 / 207 = 0
    16'b00011100_11010000 : OUT <= 0;  //28 / 208 = 0
    16'b00011100_11010001 : OUT <= 0;  //28 / 209 = 0
    16'b00011100_11010010 : OUT <= 0;  //28 / 210 = 0
    16'b00011100_11010011 : OUT <= 0;  //28 / 211 = 0
    16'b00011100_11010100 : OUT <= 0;  //28 / 212 = 0
    16'b00011100_11010101 : OUT <= 0;  //28 / 213 = 0
    16'b00011100_11010110 : OUT <= 0;  //28 / 214 = 0
    16'b00011100_11010111 : OUT <= 0;  //28 / 215 = 0
    16'b00011100_11011000 : OUT <= 0;  //28 / 216 = 0
    16'b00011100_11011001 : OUT <= 0;  //28 / 217 = 0
    16'b00011100_11011010 : OUT <= 0;  //28 / 218 = 0
    16'b00011100_11011011 : OUT <= 0;  //28 / 219 = 0
    16'b00011100_11011100 : OUT <= 0;  //28 / 220 = 0
    16'b00011100_11011101 : OUT <= 0;  //28 / 221 = 0
    16'b00011100_11011110 : OUT <= 0;  //28 / 222 = 0
    16'b00011100_11011111 : OUT <= 0;  //28 / 223 = 0
    16'b00011100_11100000 : OUT <= 0;  //28 / 224 = 0
    16'b00011100_11100001 : OUT <= 0;  //28 / 225 = 0
    16'b00011100_11100010 : OUT <= 0;  //28 / 226 = 0
    16'b00011100_11100011 : OUT <= 0;  //28 / 227 = 0
    16'b00011100_11100100 : OUT <= 0;  //28 / 228 = 0
    16'b00011100_11100101 : OUT <= 0;  //28 / 229 = 0
    16'b00011100_11100110 : OUT <= 0;  //28 / 230 = 0
    16'b00011100_11100111 : OUT <= 0;  //28 / 231 = 0
    16'b00011100_11101000 : OUT <= 0;  //28 / 232 = 0
    16'b00011100_11101001 : OUT <= 0;  //28 / 233 = 0
    16'b00011100_11101010 : OUT <= 0;  //28 / 234 = 0
    16'b00011100_11101011 : OUT <= 0;  //28 / 235 = 0
    16'b00011100_11101100 : OUT <= 0;  //28 / 236 = 0
    16'b00011100_11101101 : OUT <= 0;  //28 / 237 = 0
    16'b00011100_11101110 : OUT <= 0;  //28 / 238 = 0
    16'b00011100_11101111 : OUT <= 0;  //28 / 239 = 0
    16'b00011100_11110000 : OUT <= 0;  //28 / 240 = 0
    16'b00011100_11110001 : OUT <= 0;  //28 / 241 = 0
    16'b00011100_11110010 : OUT <= 0;  //28 / 242 = 0
    16'b00011100_11110011 : OUT <= 0;  //28 / 243 = 0
    16'b00011100_11110100 : OUT <= 0;  //28 / 244 = 0
    16'b00011100_11110101 : OUT <= 0;  //28 / 245 = 0
    16'b00011100_11110110 : OUT <= 0;  //28 / 246 = 0
    16'b00011100_11110111 : OUT <= 0;  //28 / 247 = 0
    16'b00011100_11111000 : OUT <= 0;  //28 / 248 = 0
    16'b00011100_11111001 : OUT <= 0;  //28 / 249 = 0
    16'b00011100_11111010 : OUT <= 0;  //28 / 250 = 0
    16'b00011100_11111011 : OUT <= 0;  //28 / 251 = 0
    16'b00011100_11111100 : OUT <= 0;  //28 / 252 = 0
    16'b00011100_11111101 : OUT <= 0;  //28 / 253 = 0
    16'b00011100_11111110 : OUT <= 0;  //28 / 254 = 0
    16'b00011100_11111111 : OUT <= 0;  //28 / 255 = 0
    16'b00011101_00000000 : OUT <= 0;  //29 / 0 = 0
    16'b00011101_00000001 : OUT <= 29;  //29 / 1 = 29
    16'b00011101_00000010 : OUT <= 14;  //29 / 2 = 14
    16'b00011101_00000011 : OUT <= 9;  //29 / 3 = 9
    16'b00011101_00000100 : OUT <= 7;  //29 / 4 = 7
    16'b00011101_00000101 : OUT <= 5;  //29 / 5 = 5
    16'b00011101_00000110 : OUT <= 4;  //29 / 6 = 4
    16'b00011101_00000111 : OUT <= 4;  //29 / 7 = 4
    16'b00011101_00001000 : OUT <= 3;  //29 / 8 = 3
    16'b00011101_00001001 : OUT <= 3;  //29 / 9 = 3
    16'b00011101_00001010 : OUT <= 2;  //29 / 10 = 2
    16'b00011101_00001011 : OUT <= 2;  //29 / 11 = 2
    16'b00011101_00001100 : OUT <= 2;  //29 / 12 = 2
    16'b00011101_00001101 : OUT <= 2;  //29 / 13 = 2
    16'b00011101_00001110 : OUT <= 2;  //29 / 14 = 2
    16'b00011101_00001111 : OUT <= 1;  //29 / 15 = 1
    16'b00011101_00010000 : OUT <= 1;  //29 / 16 = 1
    16'b00011101_00010001 : OUT <= 1;  //29 / 17 = 1
    16'b00011101_00010010 : OUT <= 1;  //29 / 18 = 1
    16'b00011101_00010011 : OUT <= 1;  //29 / 19 = 1
    16'b00011101_00010100 : OUT <= 1;  //29 / 20 = 1
    16'b00011101_00010101 : OUT <= 1;  //29 / 21 = 1
    16'b00011101_00010110 : OUT <= 1;  //29 / 22 = 1
    16'b00011101_00010111 : OUT <= 1;  //29 / 23 = 1
    16'b00011101_00011000 : OUT <= 1;  //29 / 24 = 1
    16'b00011101_00011001 : OUT <= 1;  //29 / 25 = 1
    16'b00011101_00011010 : OUT <= 1;  //29 / 26 = 1
    16'b00011101_00011011 : OUT <= 1;  //29 / 27 = 1
    16'b00011101_00011100 : OUT <= 1;  //29 / 28 = 1
    16'b00011101_00011101 : OUT <= 1;  //29 / 29 = 1
    16'b00011101_00011110 : OUT <= 0;  //29 / 30 = 0
    16'b00011101_00011111 : OUT <= 0;  //29 / 31 = 0
    16'b00011101_00100000 : OUT <= 0;  //29 / 32 = 0
    16'b00011101_00100001 : OUT <= 0;  //29 / 33 = 0
    16'b00011101_00100010 : OUT <= 0;  //29 / 34 = 0
    16'b00011101_00100011 : OUT <= 0;  //29 / 35 = 0
    16'b00011101_00100100 : OUT <= 0;  //29 / 36 = 0
    16'b00011101_00100101 : OUT <= 0;  //29 / 37 = 0
    16'b00011101_00100110 : OUT <= 0;  //29 / 38 = 0
    16'b00011101_00100111 : OUT <= 0;  //29 / 39 = 0
    16'b00011101_00101000 : OUT <= 0;  //29 / 40 = 0
    16'b00011101_00101001 : OUT <= 0;  //29 / 41 = 0
    16'b00011101_00101010 : OUT <= 0;  //29 / 42 = 0
    16'b00011101_00101011 : OUT <= 0;  //29 / 43 = 0
    16'b00011101_00101100 : OUT <= 0;  //29 / 44 = 0
    16'b00011101_00101101 : OUT <= 0;  //29 / 45 = 0
    16'b00011101_00101110 : OUT <= 0;  //29 / 46 = 0
    16'b00011101_00101111 : OUT <= 0;  //29 / 47 = 0
    16'b00011101_00110000 : OUT <= 0;  //29 / 48 = 0
    16'b00011101_00110001 : OUT <= 0;  //29 / 49 = 0
    16'b00011101_00110010 : OUT <= 0;  //29 / 50 = 0
    16'b00011101_00110011 : OUT <= 0;  //29 / 51 = 0
    16'b00011101_00110100 : OUT <= 0;  //29 / 52 = 0
    16'b00011101_00110101 : OUT <= 0;  //29 / 53 = 0
    16'b00011101_00110110 : OUT <= 0;  //29 / 54 = 0
    16'b00011101_00110111 : OUT <= 0;  //29 / 55 = 0
    16'b00011101_00111000 : OUT <= 0;  //29 / 56 = 0
    16'b00011101_00111001 : OUT <= 0;  //29 / 57 = 0
    16'b00011101_00111010 : OUT <= 0;  //29 / 58 = 0
    16'b00011101_00111011 : OUT <= 0;  //29 / 59 = 0
    16'b00011101_00111100 : OUT <= 0;  //29 / 60 = 0
    16'b00011101_00111101 : OUT <= 0;  //29 / 61 = 0
    16'b00011101_00111110 : OUT <= 0;  //29 / 62 = 0
    16'b00011101_00111111 : OUT <= 0;  //29 / 63 = 0
    16'b00011101_01000000 : OUT <= 0;  //29 / 64 = 0
    16'b00011101_01000001 : OUT <= 0;  //29 / 65 = 0
    16'b00011101_01000010 : OUT <= 0;  //29 / 66 = 0
    16'b00011101_01000011 : OUT <= 0;  //29 / 67 = 0
    16'b00011101_01000100 : OUT <= 0;  //29 / 68 = 0
    16'b00011101_01000101 : OUT <= 0;  //29 / 69 = 0
    16'b00011101_01000110 : OUT <= 0;  //29 / 70 = 0
    16'b00011101_01000111 : OUT <= 0;  //29 / 71 = 0
    16'b00011101_01001000 : OUT <= 0;  //29 / 72 = 0
    16'b00011101_01001001 : OUT <= 0;  //29 / 73 = 0
    16'b00011101_01001010 : OUT <= 0;  //29 / 74 = 0
    16'b00011101_01001011 : OUT <= 0;  //29 / 75 = 0
    16'b00011101_01001100 : OUT <= 0;  //29 / 76 = 0
    16'b00011101_01001101 : OUT <= 0;  //29 / 77 = 0
    16'b00011101_01001110 : OUT <= 0;  //29 / 78 = 0
    16'b00011101_01001111 : OUT <= 0;  //29 / 79 = 0
    16'b00011101_01010000 : OUT <= 0;  //29 / 80 = 0
    16'b00011101_01010001 : OUT <= 0;  //29 / 81 = 0
    16'b00011101_01010010 : OUT <= 0;  //29 / 82 = 0
    16'b00011101_01010011 : OUT <= 0;  //29 / 83 = 0
    16'b00011101_01010100 : OUT <= 0;  //29 / 84 = 0
    16'b00011101_01010101 : OUT <= 0;  //29 / 85 = 0
    16'b00011101_01010110 : OUT <= 0;  //29 / 86 = 0
    16'b00011101_01010111 : OUT <= 0;  //29 / 87 = 0
    16'b00011101_01011000 : OUT <= 0;  //29 / 88 = 0
    16'b00011101_01011001 : OUT <= 0;  //29 / 89 = 0
    16'b00011101_01011010 : OUT <= 0;  //29 / 90 = 0
    16'b00011101_01011011 : OUT <= 0;  //29 / 91 = 0
    16'b00011101_01011100 : OUT <= 0;  //29 / 92 = 0
    16'b00011101_01011101 : OUT <= 0;  //29 / 93 = 0
    16'b00011101_01011110 : OUT <= 0;  //29 / 94 = 0
    16'b00011101_01011111 : OUT <= 0;  //29 / 95 = 0
    16'b00011101_01100000 : OUT <= 0;  //29 / 96 = 0
    16'b00011101_01100001 : OUT <= 0;  //29 / 97 = 0
    16'b00011101_01100010 : OUT <= 0;  //29 / 98 = 0
    16'b00011101_01100011 : OUT <= 0;  //29 / 99 = 0
    16'b00011101_01100100 : OUT <= 0;  //29 / 100 = 0
    16'b00011101_01100101 : OUT <= 0;  //29 / 101 = 0
    16'b00011101_01100110 : OUT <= 0;  //29 / 102 = 0
    16'b00011101_01100111 : OUT <= 0;  //29 / 103 = 0
    16'b00011101_01101000 : OUT <= 0;  //29 / 104 = 0
    16'b00011101_01101001 : OUT <= 0;  //29 / 105 = 0
    16'b00011101_01101010 : OUT <= 0;  //29 / 106 = 0
    16'b00011101_01101011 : OUT <= 0;  //29 / 107 = 0
    16'b00011101_01101100 : OUT <= 0;  //29 / 108 = 0
    16'b00011101_01101101 : OUT <= 0;  //29 / 109 = 0
    16'b00011101_01101110 : OUT <= 0;  //29 / 110 = 0
    16'b00011101_01101111 : OUT <= 0;  //29 / 111 = 0
    16'b00011101_01110000 : OUT <= 0;  //29 / 112 = 0
    16'b00011101_01110001 : OUT <= 0;  //29 / 113 = 0
    16'b00011101_01110010 : OUT <= 0;  //29 / 114 = 0
    16'b00011101_01110011 : OUT <= 0;  //29 / 115 = 0
    16'b00011101_01110100 : OUT <= 0;  //29 / 116 = 0
    16'b00011101_01110101 : OUT <= 0;  //29 / 117 = 0
    16'b00011101_01110110 : OUT <= 0;  //29 / 118 = 0
    16'b00011101_01110111 : OUT <= 0;  //29 / 119 = 0
    16'b00011101_01111000 : OUT <= 0;  //29 / 120 = 0
    16'b00011101_01111001 : OUT <= 0;  //29 / 121 = 0
    16'b00011101_01111010 : OUT <= 0;  //29 / 122 = 0
    16'b00011101_01111011 : OUT <= 0;  //29 / 123 = 0
    16'b00011101_01111100 : OUT <= 0;  //29 / 124 = 0
    16'b00011101_01111101 : OUT <= 0;  //29 / 125 = 0
    16'b00011101_01111110 : OUT <= 0;  //29 / 126 = 0
    16'b00011101_01111111 : OUT <= 0;  //29 / 127 = 0
    16'b00011101_10000000 : OUT <= 0;  //29 / 128 = 0
    16'b00011101_10000001 : OUT <= 0;  //29 / 129 = 0
    16'b00011101_10000010 : OUT <= 0;  //29 / 130 = 0
    16'b00011101_10000011 : OUT <= 0;  //29 / 131 = 0
    16'b00011101_10000100 : OUT <= 0;  //29 / 132 = 0
    16'b00011101_10000101 : OUT <= 0;  //29 / 133 = 0
    16'b00011101_10000110 : OUT <= 0;  //29 / 134 = 0
    16'b00011101_10000111 : OUT <= 0;  //29 / 135 = 0
    16'b00011101_10001000 : OUT <= 0;  //29 / 136 = 0
    16'b00011101_10001001 : OUT <= 0;  //29 / 137 = 0
    16'b00011101_10001010 : OUT <= 0;  //29 / 138 = 0
    16'b00011101_10001011 : OUT <= 0;  //29 / 139 = 0
    16'b00011101_10001100 : OUT <= 0;  //29 / 140 = 0
    16'b00011101_10001101 : OUT <= 0;  //29 / 141 = 0
    16'b00011101_10001110 : OUT <= 0;  //29 / 142 = 0
    16'b00011101_10001111 : OUT <= 0;  //29 / 143 = 0
    16'b00011101_10010000 : OUT <= 0;  //29 / 144 = 0
    16'b00011101_10010001 : OUT <= 0;  //29 / 145 = 0
    16'b00011101_10010010 : OUT <= 0;  //29 / 146 = 0
    16'b00011101_10010011 : OUT <= 0;  //29 / 147 = 0
    16'b00011101_10010100 : OUT <= 0;  //29 / 148 = 0
    16'b00011101_10010101 : OUT <= 0;  //29 / 149 = 0
    16'b00011101_10010110 : OUT <= 0;  //29 / 150 = 0
    16'b00011101_10010111 : OUT <= 0;  //29 / 151 = 0
    16'b00011101_10011000 : OUT <= 0;  //29 / 152 = 0
    16'b00011101_10011001 : OUT <= 0;  //29 / 153 = 0
    16'b00011101_10011010 : OUT <= 0;  //29 / 154 = 0
    16'b00011101_10011011 : OUT <= 0;  //29 / 155 = 0
    16'b00011101_10011100 : OUT <= 0;  //29 / 156 = 0
    16'b00011101_10011101 : OUT <= 0;  //29 / 157 = 0
    16'b00011101_10011110 : OUT <= 0;  //29 / 158 = 0
    16'b00011101_10011111 : OUT <= 0;  //29 / 159 = 0
    16'b00011101_10100000 : OUT <= 0;  //29 / 160 = 0
    16'b00011101_10100001 : OUT <= 0;  //29 / 161 = 0
    16'b00011101_10100010 : OUT <= 0;  //29 / 162 = 0
    16'b00011101_10100011 : OUT <= 0;  //29 / 163 = 0
    16'b00011101_10100100 : OUT <= 0;  //29 / 164 = 0
    16'b00011101_10100101 : OUT <= 0;  //29 / 165 = 0
    16'b00011101_10100110 : OUT <= 0;  //29 / 166 = 0
    16'b00011101_10100111 : OUT <= 0;  //29 / 167 = 0
    16'b00011101_10101000 : OUT <= 0;  //29 / 168 = 0
    16'b00011101_10101001 : OUT <= 0;  //29 / 169 = 0
    16'b00011101_10101010 : OUT <= 0;  //29 / 170 = 0
    16'b00011101_10101011 : OUT <= 0;  //29 / 171 = 0
    16'b00011101_10101100 : OUT <= 0;  //29 / 172 = 0
    16'b00011101_10101101 : OUT <= 0;  //29 / 173 = 0
    16'b00011101_10101110 : OUT <= 0;  //29 / 174 = 0
    16'b00011101_10101111 : OUT <= 0;  //29 / 175 = 0
    16'b00011101_10110000 : OUT <= 0;  //29 / 176 = 0
    16'b00011101_10110001 : OUT <= 0;  //29 / 177 = 0
    16'b00011101_10110010 : OUT <= 0;  //29 / 178 = 0
    16'b00011101_10110011 : OUT <= 0;  //29 / 179 = 0
    16'b00011101_10110100 : OUT <= 0;  //29 / 180 = 0
    16'b00011101_10110101 : OUT <= 0;  //29 / 181 = 0
    16'b00011101_10110110 : OUT <= 0;  //29 / 182 = 0
    16'b00011101_10110111 : OUT <= 0;  //29 / 183 = 0
    16'b00011101_10111000 : OUT <= 0;  //29 / 184 = 0
    16'b00011101_10111001 : OUT <= 0;  //29 / 185 = 0
    16'b00011101_10111010 : OUT <= 0;  //29 / 186 = 0
    16'b00011101_10111011 : OUT <= 0;  //29 / 187 = 0
    16'b00011101_10111100 : OUT <= 0;  //29 / 188 = 0
    16'b00011101_10111101 : OUT <= 0;  //29 / 189 = 0
    16'b00011101_10111110 : OUT <= 0;  //29 / 190 = 0
    16'b00011101_10111111 : OUT <= 0;  //29 / 191 = 0
    16'b00011101_11000000 : OUT <= 0;  //29 / 192 = 0
    16'b00011101_11000001 : OUT <= 0;  //29 / 193 = 0
    16'b00011101_11000010 : OUT <= 0;  //29 / 194 = 0
    16'b00011101_11000011 : OUT <= 0;  //29 / 195 = 0
    16'b00011101_11000100 : OUT <= 0;  //29 / 196 = 0
    16'b00011101_11000101 : OUT <= 0;  //29 / 197 = 0
    16'b00011101_11000110 : OUT <= 0;  //29 / 198 = 0
    16'b00011101_11000111 : OUT <= 0;  //29 / 199 = 0
    16'b00011101_11001000 : OUT <= 0;  //29 / 200 = 0
    16'b00011101_11001001 : OUT <= 0;  //29 / 201 = 0
    16'b00011101_11001010 : OUT <= 0;  //29 / 202 = 0
    16'b00011101_11001011 : OUT <= 0;  //29 / 203 = 0
    16'b00011101_11001100 : OUT <= 0;  //29 / 204 = 0
    16'b00011101_11001101 : OUT <= 0;  //29 / 205 = 0
    16'b00011101_11001110 : OUT <= 0;  //29 / 206 = 0
    16'b00011101_11001111 : OUT <= 0;  //29 / 207 = 0
    16'b00011101_11010000 : OUT <= 0;  //29 / 208 = 0
    16'b00011101_11010001 : OUT <= 0;  //29 / 209 = 0
    16'b00011101_11010010 : OUT <= 0;  //29 / 210 = 0
    16'b00011101_11010011 : OUT <= 0;  //29 / 211 = 0
    16'b00011101_11010100 : OUT <= 0;  //29 / 212 = 0
    16'b00011101_11010101 : OUT <= 0;  //29 / 213 = 0
    16'b00011101_11010110 : OUT <= 0;  //29 / 214 = 0
    16'b00011101_11010111 : OUT <= 0;  //29 / 215 = 0
    16'b00011101_11011000 : OUT <= 0;  //29 / 216 = 0
    16'b00011101_11011001 : OUT <= 0;  //29 / 217 = 0
    16'b00011101_11011010 : OUT <= 0;  //29 / 218 = 0
    16'b00011101_11011011 : OUT <= 0;  //29 / 219 = 0
    16'b00011101_11011100 : OUT <= 0;  //29 / 220 = 0
    16'b00011101_11011101 : OUT <= 0;  //29 / 221 = 0
    16'b00011101_11011110 : OUT <= 0;  //29 / 222 = 0
    16'b00011101_11011111 : OUT <= 0;  //29 / 223 = 0
    16'b00011101_11100000 : OUT <= 0;  //29 / 224 = 0
    16'b00011101_11100001 : OUT <= 0;  //29 / 225 = 0
    16'b00011101_11100010 : OUT <= 0;  //29 / 226 = 0
    16'b00011101_11100011 : OUT <= 0;  //29 / 227 = 0
    16'b00011101_11100100 : OUT <= 0;  //29 / 228 = 0
    16'b00011101_11100101 : OUT <= 0;  //29 / 229 = 0
    16'b00011101_11100110 : OUT <= 0;  //29 / 230 = 0
    16'b00011101_11100111 : OUT <= 0;  //29 / 231 = 0
    16'b00011101_11101000 : OUT <= 0;  //29 / 232 = 0
    16'b00011101_11101001 : OUT <= 0;  //29 / 233 = 0
    16'b00011101_11101010 : OUT <= 0;  //29 / 234 = 0
    16'b00011101_11101011 : OUT <= 0;  //29 / 235 = 0
    16'b00011101_11101100 : OUT <= 0;  //29 / 236 = 0
    16'b00011101_11101101 : OUT <= 0;  //29 / 237 = 0
    16'b00011101_11101110 : OUT <= 0;  //29 / 238 = 0
    16'b00011101_11101111 : OUT <= 0;  //29 / 239 = 0
    16'b00011101_11110000 : OUT <= 0;  //29 / 240 = 0
    16'b00011101_11110001 : OUT <= 0;  //29 / 241 = 0
    16'b00011101_11110010 : OUT <= 0;  //29 / 242 = 0
    16'b00011101_11110011 : OUT <= 0;  //29 / 243 = 0
    16'b00011101_11110100 : OUT <= 0;  //29 / 244 = 0
    16'b00011101_11110101 : OUT <= 0;  //29 / 245 = 0
    16'b00011101_11110110 : OUT <= 0;  //29 / 246 = 0
    16'b00011101_11110111 : OUT <= 0;  //29 / 247 = 0
    16'b00011101_11111000 : OUT <= 0;  //29 / 248 = 0
    16'b00011101_11111001 : OUT <= 0;  //29 / 249 = 0
    16'b00011101_11111010 : OUT <= 0;  //29 / 250 = 0
    16'b00011101_11111011 : OUT <= 0;  //29 / 251 = 0
    16'b00011101_11111100 : OUT <= 0;  //29 / 252 = 0
    16'b00011101_11111101 : OUT <= 0;  //29 / 253 = 0
    16'b00011101_11111110 : OUT <= 0;  //29 / 254 = 0
    16'b00011101_11111111 : OUT <= 0;  //29 / 255 = 0
    16'b00011110_00000000 : OUT <= 0;  //30 / 0 = 0
    16'b00011110_00000001 : OUT <= 30;  //30 / 1 = 30
    16'b00011110_00000010 : OUT <= 15;  //30 / 2 = 15
    16'b00011110_00000011 : OUT <= 10;  //30 / 3 = 10
    16'b00011110_00000100 : OUT <= 7;  //30 / 4 = 7
    16'b00011110_00000101 : OUT <= 6;  //30 / 5 = 6
    16'b00011110_00000110 : OUT <= 5;  //30 / 6 = 5
    16'b00011110_00000111 : OUT <= 4;  //30 / 7 = 4
    16'b00011110_00001000 : OUT <= 3;  //30 / 8 = 3
    16'b00011110_00001001 : OUT <= 3;  //30 / 9 = 3
    16'b00011110_00001010 : OUT <= 3;  //30 / 10 = 3
    16'b00011110_00001011 : OUT <= 2;  //30 / 11 = 2
    16'b00011110_00001100 : OUT <= 2;  //30 / 12 = 2
    16'b00011110_00001101 : OUT <= 2;  //30 / 13 = 2
    16'b00011110_00001110 : OUT <= 2;  //30 / 14 = 2
    16'b00011110_00001111 : OUT <= 2;  //30 / 15 = 2
    16'b00011110_00010000 : OUT <= 1;  //30 / 16 = 1
    16'b00011110_00010001 : OUT <= 1;  //30 / 17 = 1
    16'b00011110_00010010 : OUT <= 1;  //30 / 18 = 1
    16'b00011110_00010011 : OUT <= 1;  //30 / 19 = 1
    16'b00011110_00010100 : OUT <= 1;  //30 / 20 = 1
    16'b00011110_00010101 : OUT <= 1;  //30 / 21 = 1
    16'b00011110_00010110 : OUT <= 1;  //30 / 22 = 1
    16'b00011110_00010111 : OUT <= 1;  //30 / 23 = 1
    16'b00011110_00011000 : OUT <= 1;  //30 / 24 = 1
    16'b00011110_00011001 : OUT <= 1;  //30 / 25 = 1
    16'b00011110_00011010 : OUT <= 1;  //30 / 26 = 1
    16'b00011110_00011011 : OUT <= 1;  //30 / 27 = 1
    16'b00011110_00011100 : OUT <= 1;  //30 / 28 = 1
    16'b00011110_00011101 : OUT <= 1;  //30 / 29 = 1
    16'b00011110_00011110 : OUT <= 1;  //30 / 30 = 1
    16'b00011110_00011111 : OUT <= 0;  //30 / 31 = 0
    16'b00011110_00100000 : OUT <= 0;  //30 / 32 = 0
    16'b00011110_00100001 : OUT <= 0;  //30 / 33 = 0
    16'b00011110_00100010 : OUT <= 0;  //30 / 34 = 0
    16'b00011110_00100011 : OUT <= 0;  //30 / 35 = 0
    16'b00011110_00100100 : OUT <= 0;  //30 / 36 = 0
    16'b00011110_00100101 : OUT <= 0;  //30 / 37 = 0
    16'b00011110_00100110 : OUT <= 0;  //30 / 38 = 0
    16'b00011110_00100111 : OUT <= 0;  //30 / 39 = 0
    16'b00011110_00101000 : OUT <= 0;  //30 / 40 = 0
    16'b00011110_00101001 : OUT <= 0;  //30 / 41 = 0
    16'b00011110_00101010 : OUT <= 0;  //30 / 42 = 0
    16'b00011110_00101011 : OUT <= 0;  //30 / 43 = 0
    16'b00011110_00101100 : OUT <= 0;  //30 / 44 = 0
    16'b00011110_00101101 : OUT <= 0;  //30 / 45 = 0
    16'b00011110_00101110 : OUT <= 0;  //30 / 46 = 0
    16'b00011110_00101111 : OUT <= 0;  //30 / 47 = 0
    16'b00011110_00110000 : OUT <= 0;  //30 / 48 = 0
    16'b00011110_00110001 : OUT <= 0;  //30 / 49 = 0
    16'b00011110_00110010 : OUT <= 0;  //30 / 50 = 0
    16'b00011110_00110011 : OUT <= 0;  //30 / 51 = 0
    16'b00011110_00110100 : OUT <= 0;  //30 / 52 = 0
    16'b00011110_00110101 : OUT <= 0;  //30 / 53 = 0
    16'b00011110_00110110 : OUT <= 0;  //30 / 54 = 0
    16'b00011110_00110111 : OUT <= 0;  //30 / 55 = 0
    16'b00011110_00111000 : OUT <= 0;  //30 / 56 = 0
    16'b00011110_00111001 : OUT <= 0;  //30 / 57 = 0
    16'b00011110_00111010 : OUT <= 0;  //30 / 58 = 0
    16'b00011110_00111011 : OUT <= 0;  //30 / 59 = 0
    16'b00011110_00111100 : OUT <= 0;  //30 / 60 = 0
    16'b00011110_00111101 : OUT <= 0;  //30 / 61 = 0
    16'b00011110_00111110 : OUT <= 0;  //30 / 62 = 0
    16'b00011110_00111111 : OUT <= 0;  //30 / 63 = 0
    16'b00011110_01000000 : OUT <= 0;  //30 / 64 = 0
    16'b00011110_01000001 : OUT <= 0;  //30 / 65 = 0
    16'b00011110_01000010 : OUT <= 0;  //30 / 66 = 0
    16'b00011110_01000011 : OUT <= 0;  //30 / 67 = 0
    16'b00011110_01000100 : OUT <= 0;  //30 / 68 = 0
    16'b00011110_01000101 : OUT <= 0;  //30 / 69 = 0
    16'b00011110_01000110 : OUT <= 0;  //30 / 70 = 0
    16'b00011110_01000111 : OUT <= 0;  //30 / 71 = 0
    16'b00011110_01001000 : OUT <= 0;  //30 / 72 = 0
    16'b00011110_01001001 : OUT <= 0;  //30 / 73 = 0
    16'b00011110_01001010 : OUT <= 0;  //30 / 74 = 0
    16'b00011110_01001011 : OUT <= 0;  //30 / 75 = 0
    16'b00011110_01001100 : OUT <= 0;  //30 / 76 = 0
    16'b00011110_01001101 : OUT <= 0;  //30 / 77 = 0
    16'b00011110_01001110 : OUT <= 0;  //30 / 78 = 0
    16'b00011110_01001111 : OUT <= 0;  //30 / 79 = 0
    16'b00011110_01010000 : OUT <= 0;  //30 / 80 = 0
    16'b00011110_01010001 : OUT <= 0;  //30 / 81 = 0
    16'b00011110_01010010 : OUT <= 0;  //30 / 82 = 0
    16'b00011110_01010011 : OUT <= 0;  //30 / 83 = 0
    16'b00011110_01010100 : OUT <= 0;  //30 / 84 = 0
    16'b00011110_01010101 : OUT <= 0;  //30 / 85 = 0
    16'b00011110_01010110 : OUT <= 0;  //30 / 86 = 0
    16'b00011110_01010111 : OUT <= 0;  //30 / 87 = 0
    16'b00011110_01011000 : OUT <= 0;  //30 / 88 = 0
    16'b00011110_01011001 : OUT <= 0;  //30 / 89 = 0
    16'b00011110_01011010 : OUT <= 0;  //30 / 90 = 0
    16'b00011110_01011011 : OUT <= 0;  //30 / 91 = 0
    16'b00011110_01011100 : OUT <= 0;  //30 / 92 = 0
    16'b00011110_01011101 : OUT <= 0;  //30 / 93 = 0
    16'b00011110_01011110 : OUT <= 0;  //30 / 94 = 0
    16'b00011110_01011111 : OUT <= 0;  //30 / 95 = 0
    16'b00011110_01100000 : OUT <= 0;  //30 / 96 = 0
    16'b00011110_01100001 : OUT <= 0;  //30 / 97 = 0
    16'b00011110_01100010 : OUT <= 0;  //30 / 98 = 0
    16'b00011110_01100011 : OUT <= 0;  //30 / 99 = 0
    16'b00011110_01100100 : OUT <= 0;  //30 / 100 = 0
    16'b00011110_01100101 : OUT <= 0;  //30 / 101 = 0
    16'b00011110_01100110 : OUT <= 0;  //30 / 102 = 0
    16'b00011110_01100111 : OUT <= 0;  //30 / 103 = 0
    16'b00011110_01101000 : OUT <= 0;  //30 / 104 = 0
    16'b00011110_01101001 : OUT <= 0;  //30 / 105 = 0
    16'b00011110_01101010 : OUT <= 0;  //30 / 106 = 0
    16'b00011110_01101011 : OUT <= 0;  //30 / 107 = 0
    16'b00011110_01101100 : OUT <= 0;  //30 / 108 = 0
    16'b00011110_01101101 : OUT <= 0;  //30 / 109 = 0
    16'b00011110_01101110 : OUT <= 0;  //30 / 110 = 0
    16'b00011110_01101111 : OUT <= 0;  //30 / 111 = 0
    16'b00011110_01110000 : OUT <= 0;  //30 / 112 = 0
    16'b00011110_01110001 : OUT <= 0;  //30 / 113 = 0
    16'b00011110_01110010 : OUT <= 0;  //30 / 114 = 0
    16'b00011110_01110011 : OUT <= 0;  //30 / 115 = 0
    16'b00011110_01110100 : OUT <= 0;  //30 / 116 = 0
    16'b00011110_01110101 : OUT <= 0;  //30 / 117 = 0
    16'b00011110_01110110 : OUT <= 0;  //30 / 118 = 0
    16'b00011110_01110111 : OUT <= 0;  //30 / 119 = 0
    16'b00011110_01111000 : OUT <= 0;  //30 / 120 = 0
    16'b00011110_01111001 : OUT <= 0;  //30 / 121 = 0
    16'b00011110_01111010 : OUT <= 0;  //30 / 122 = 0
    16'b00011110_01111011 : OUT <= 0;  //30 / 123 = 0
    16'b00011110_01111100 : OUT <= 0;  //30 / 124 = 0
    16'b00011110_01111101 : OUT <= 0;  //30 / 125 = 0
    16'b00011110_01111110 : OUT <= 0;  //30 / 126 = 0
    16'b00011110_01111111 : OUT <= 0;  //30 / 127 = 0
    16'b00011110_10000000 : OUT <= 0;  //30 / 128 = 0
    16'b00011110_10000001 : OUT <= 0;  //30 / 129 = 0
    16'b00011110_10000010 : OUT <= 0;  //30 / 130 = 0
    16'b00011110_10000011 : OUT <= 0;  //30 / 131 = 0
    16'b00011110_10000100 : OUT <= 0;  //30 / 132 = 0
    16'b00011110_10000101 : OUT <= 0;  //30 / 133 = 0
    16'b00011110_10000110 : OUT <= 0;  //30 / 134 = 0
    16'b00011110_10000111 : OUT <= 0;  //30 / 135 = 0
    16'b00011110_10001000 : OUT <= 0;  //30 / 136 = 0
    16'b00011110_10001001 : OUT <= 0;  //30 / 137 = 0
    16'b00011110_10001010 : OUT <= 0;  //30 / 138 = 0
    16'b00011110_10001011 : OUT <= 0;  //30 / 139 = 0
    16'b00011110_10001100 : OUT <= 0;  //30 / 140 = 0
    16'b00011110_10001101 : OUT <= 0;  //30 / 141 = 0
    16'b00011110_10001110 : OUT <= 0;  //30 / 142 = 0
    16'b00011110_10001111 : OUT <= 0;  //30 / 143 = 0
    16'b00011110_10010000 : OUT <= 0;  //30 / 144 = 0
    16'b00011110_10010001 : OUT <= 0;  //30 / 145 = 0
    16'b00011110_10010010 : OUT <= 0;  //30 / 146 = 0
    16'b00011110_10010011 : OUT <= 0;  //30 / 147 = 0
    16'b00011110_10010100 : OUT <= 0;  //30 / 148 = 0
    16'b00011110_10010101 : OUT <= 0;  //30 / 149 = 0
    16'b00011110_10010110 : OUT <= 0;  //30 / 150 = 0
    16'b00011110_10010111 : OUT <= 0;  //30 / 151 = 0
    16'b00011110_10011000 : OUT <= 0;  //30 / 152 = 0
    16'b00011110_10011001 : OUT <= 0;  //30 / 153 = 0
    16'b00011110_10011010 : OUT <= 0;  //30 / 154 = 0
    16'b00011110_10011011 : OUT <= 0;  //30 / 155 = 0
    16'b00011110_10011100 : OUT <= 0;  //30 / 156 = 0
    16'b00011110_10011101 : OUT <= 0;  //30 / 157 = 0
    16'b00011110_10011110 : OUT <= 0;  //30 / 158 = 0
    16'b00011110_10011111 : OUT <= 0;  //30 / 159 = 0
    16'b00011110_10100000 : OUT <= 0;  //30 / 160 = 0
    16'b00011110_10100001 : OUT <= 0;  //30 / 161 = 0
    16'b00011110_10100010 : OUT <= 0;  //30 / 162 = 0
    16'b00011110_10100011 : OUT <= 0;  //30 / 163 = 0
    16'b00011110_10100100 : OUT <= 0;  //30 / 164 = 0
    16'b00011110_10100101 : OUT <= 0;  //30 / 165 = 0
    16'b00011110_10100110 : OUT <= 0;  //30 / 166 = 0
    16'b00011110_10100111 : OUT <= 0;  //30 / 167 = 0
    16'b00011110_10101000 : OUT <= 0;  //30 / 168 = 0
    16'b00011110_10101001 : OUT <= 0;  //30 / 169 = 0
    16'b00011110_10101010 : OUT <= 0;  //30 / 170 = 0
    16'b00011110_10101011 : OUT <= 0;  //30 / 171 = 0
    16'b00011110_10101100 : OUT <= 0;  //30 / 172 = 0
    16'b00011110_10101101 : OUT <= 0;  //30 / 173 = 0
    16'b00011110_10101110 : OUT <= 0;  //30 / 174 = 0
    16'b00011110_10101111 : OUT <= 0;  //30 / 175 = 0
    16'b00011110_10110000 : OUT <= 0;  //30 / 176 = 0
    16'b00011110_10110001 : OUT <= 0;  //30 / 177 = 0
    16'b00011110_10110010 : OUT <= 0;  //30 / 178 = 0
    16'b00011110_10110011 : OUT <= 0;  //30 / 179 = 0
    16'b00011110_10110100 : OUT <= 0;  //30 / 180 = 0
    16'b00011110_10110101 : OUT <= 0;  //30 / 181 = 0
    16'b00011110_10110110 : OUT <= 0;  //30 / 182 = 0
    16'b00011110_10110111 : OUT <= 0;  //30 / 183 = 0
    16'b00011110_10111000 : OUT <= 0;  //30 / 184 = 0
    16'b00011110_10111001 : OUT <= 0;  //30 / 185 = 0
    16'b00011110_10111010 : OUT <= 0;  //30 / 186 = 0
    16'b00011110_10111011 : OUT <= 0;  //30 / 187 = 0
    16'b00011110_10111100 : OUT <= 0;  //30 / 188 = 0
    16'b00011110_10111101 : OUT <= 0;  //30 / 189 = 0
    16'b00011110_10111110 : OUT <= 0;  //30 / 190 = 0
    16'b00011110_10111111 : OUT <= 0;  //30 / 191 = 0
    16'b00011110_11000000 : OUT <= 0;  //30 / 192 = 0
    16'b00011110_11000001 : OUT <= 0;  //30 / 193 = 0
    16'b00011110_11000010 : OUT <= 0;  //30 / 194 = 0
    16'b00011110_11000011 : OUT <= 0;  //30 / 195 = 0
    16'b00011110_11000100 : OUT <= 0;  //30 / 196 = 0
    16'b00011110_11000101 : OUT <= 0;  //30 / 197 = 0
    16'b00011110_11000110 : OUT <= 0;  //30 / 198 = 0
    16'b00011110_11000111 : OUT <= 0;  //30 / 199 = 0
    16'b00011110_11001000 : OUT <= 0;  //30 / 200 = 0
    16'b00011110_11001001 : OUT <= 0;  //30 / 201 = 0
    16'b00011110_11001010 : OUT <= 0;  //30 / 202 = 0
    16'b00011110_11001011 : OUT <= 0;  //30 / 203 = 0
    16'b00011110_11001100 : OUT <= 0;  //30 / 204 = 0
    16'b00011110_11001101 : OUT <= 0;  //30 / 205 = 0
    16'b00011110_11001110 : OUT <= 0;  //30 / 206 = 0
    16'b00011110_11001111 : OUT <= 0;  //30 / 207 = 0
    16'b00011110_11010000 : OUT <= 0;  //30 / 208 = 0
    16'b00011110_11010001 : OUT <= 0;  //30 / 209 = 0
    16'b00011110_11010010 : OUT <= 0;  //30 / 210 = 0
    16'b00011110_11010011 : OUT <= 0;  //30 / 211 = 0
    16'b00011110_11010100 : OUT <= 0;  //30 / 212 = 0
    16'b00011110_11010101 : OUT <= 0;  //30 / 213 = 0
    16'b00011110_11010110 : OUT <= 0;  //30 / 214 = 0
    16'b00011110_11010111 : OUT <= 0;  //30 / 215 = 0
    16'b00011110_11011000 : OUT <= 0;  //30 / 216 = 0
    16'b00011110_11011001 : OUT <= 0;  //30 / 217 = 0
    16'b00011110_11011010 : OUT <= 0;  //30 / 218 = 0
    16'b00011110_11011011 : OUT <= 0;  //30 / 219 = 0
    16'b00011110_11011100 : OUT <= 0;  //30 / 220 = 0
    16'b00011110_11011101 : OUT <= 0;  //30 / 221 = 0
    16'b00011110_11011110 : OUT <= 0;  //30 / 222 = 0
    16'b00011110_11011111 : OUT <= 0;  //30 / 223 = 0
    16'b00011110_11100000 : OUT <= 0;  //30 / 224 = 0
    16'b00011110_11100001 : OUT <= 0;  //30 / 225 = 0
    16'b00011110_11100010 : OUT <= 0;  //30 / 226 = 0
    16'b00011110_11100011 : OUT <= 0;  //30 / 227 = 0
    16'b00011110_11100100 : OUT <= 0;  //30 / 228 = 0
    16'b00011110_11100101 : OUT <= 0;  //30 / 229 = 0
    16'b00011110_11100110 : OUT <= 0;  //30 / 230 = 0
    16'b00011110_11100111 : OUT <= 0;  //30 / 231 = 0
    16'b00011110_11101000 : OUT <= 0;  //30 / 232 = 0
    16'b00011110_11101001 : OUT <= 0;  //30 / 233 = 0
    16'b00011110_11101010 : OUT <= 0;  //30 / 234 = 0
    16'b00011110_11101011 : OUT <= 0;  //30 / 235 = 0
    16'b00011110_11101100 : OUT <= 0;  //30 / 236 = 0
    16'b00011110_11101101 : OUT <= 0;  //30 / 237 = 0
    16'b00011110_11101110 : OUT <= 0;  //30 / 238 = 0
    16'b00011110_11101111 : OUT <= 0;  //30 / 239 = 0
    16'b00011110_11110000 : OUT <= 0;  //30 / 240 = 0
    16'b00011110_11110001 : OUT <= 0;  //30 / 241 = 0
    16'b00011110_11110010 : OUT <= 0;  //30 / 242 = 0
    16'b00011110_11110011 : OUT <= 0;  //30 / 243 = 0
    16'b00011110_11110100 : OUT <= 0;  //30 / 244 = 0
    16'b00011110_11110101 : OUT <= 0;  //30 / 245 = 0
    16'b00011110_11110110 : OUT <= 0;  //30 / 246 = 0
    16'b00011110_11110111 : OUT <= 0;  //30 / 247 = 0
    16'b00011110_11111000 : OUT <= 0;  //30 / 248 = 0
    16'b00011110_11111001 : OUT <= 0;  //30 / 249 = 0
    16'b00011110_11111010 : OUT <= 0;  //30 / 250 = 0
    16'b00011110_11111011 : OUT <= 0;  //30 / 251 = 0
    16'b00011110_11111100 : OUT <= 0;  //30 / 252 = 0
    16'b00011110_11111101 : OUT <= 0;  //30 / 253 = 0
    16'b00011110_11111110 : OUT <= 0;  //30 / 254 = 0
    16'b00011110_11111111 : OUT <= 0;  //30 / 255 = 0
    16'b00011111_00000000 : OUT <= 0;  //31 / 0 = 0
    16'b00011111_00000001 : OUT <= 31;  //31 / 1 = 31
    16'b00011111_00000010 : OUT <= 15;  //31 / 2 = 15
    16'b00011111_00000011 : OUT <= 10;  //31 / 3 = 10
    16'b00011111_00000100 : OUT <= 7;  //31 / 4 = 7
    16'b00011111_00000101 : OUT <= 6;  //31 / 5 = 6
    16'b00011111_00000110 : OUT <= 5;  //31 / 6 = 5
    16'b00011111_00000111 : OUT <= 4;  //31 / 7 = 4
    16'b00011111_00001000 : OUT <= 3;  //31 / 8 = 3
    16'b00011111_00001001 : OUT <= 3;  //31 / 9 = 3
    16'b00011111_00001010 : OUT <= 3;  //31 / 10 = 3
    16'b00011111_00001011 : OUT <= 2;  //31 / 11 = 2
    16'b00011111_00001100 : OUT <= 2;  //31 / 12 = 2
    16'b00011111_00001101 : OUT <= 2;  //31 / 13 = 2
    16'b00011111_00001110 : OUT <= 2;  //31 / 14 = 2
    16'b00011111_00001111 : OUT <= 2;  //31 / 15 = 2
    16'b00011111_00010000 : OUT <= 1;  //31 / 16 = 1
    16'b00011111_00010001 : OUT <= 1;  //31 / 17 = 1
    16'b00011111_00010010 : OUT <= 1;  //31 / 18 = 1
    16'b00011111_00010011 : OUT <= 1;  //31 / 19 = 1
    16'b00011111_00010100 : OUT <= 1;  //31 / 20 = 1
    16'b00011111_00010101 : OUT <= 1;  //31 / 21 = 1
    16'b00011111_00010110 : OUT <= 1;  //31 / 22 = 1
    16'b00011111_00010111 : OUT <= 1;  //31 / 23 = 1
    16'b00011111_00011000 : OUT <= 1;  //31 / 24 = 1
    16'b00011111_00011001 : OUT <= 1;  //31 / 25 = 1
    16'b00011111_00011010 : OUT <= 1;  //31 / 26 = 1
    16'b00011111_00011011 : OUT <= 1;  //31 / 27 = 1
    16'b00011111_00011100 : OUT <= 1;  //31 / 28 = 1
    16'b00011111_00011101 : OUT <= 1;  //31 / 29 = 1
    16'b00011111_00011110 : OUT <= 1;  //31 / 30 = 1
    16'b00011111_00011111 : OUT <= 1;  //31 / 31 = 1
    16'b00011111_00100000 : OUT <= 0;  //31 / 32 = 0
    16'b00011111_00100001 : OUT <= 0;  //31 / 33 = 0
    16'b00011111_00100010 : OUT <= 0;  //31 / 34 = 0
    16'b00011111_00100011 : OUT <= 0;  //31 / 35 = 0
    16'b00011111_00100100 : OUT <= 0;  //31 / 36 = 0
    16'b00011111_00100101 : OUT <= 0;  //31 / 37 = 0
    16'b00011111_00100110 : OUT <= 0;  //31 / 38 = 0
    16'b00011111_00100111 : OUT <= 0;  //31 / 39 = 0
    16'b00011111_00101000 : OUT <= 0;  //31 / 40 = 0
    16'b00011111_00101001 : OUT <= 0;  //31 / 41 = 0
    16'b00011111_00101010 : OUT <= 0;  //31 / 42 = 0
    16'b00011111_00101011 : OUT <= 0;  //31 / 43 = 0
    16'b00011111_00101100 : OUT <= 0;  //31 / 44 = 0
    16'b00011111_00101101 : OUT <= 0;  //31 / 45 = 0
    16'b00011111_00101110 : OUT <= 0;  //31 / 46 = 0
    16'b00011111_00101111 : OUT <= 0;  //31 / 47 = 0
    16'b00011111_00110000 : OUT <= 0;  //31 / 48 = 0
    16'b00011111_00110001 : OUT <= 0;  //31 / 49 = 0
    16'b00011111_00110010 : OUT <= 0;  //31 / 50 = 0
    16'b00011111_00110011 : OUT <= 0;  //31 / 51 = 0
    16'b00011111_00110100 : OUT <= 0;  //31 / 52 = 0
    16'b00011111_00110101 : OUT <= 0;  //31 / 53 = 0
    16'b00011111_00110110 : OUT <= 0;  //31 / 54 = 0
    16'b00011111_00110111 : OUT <= 0;  //31 / 55 = 0
    16'b00011111_00111000 : OUT <= 0;  //31 / 56 = 0
    16'b00011111_00111001 : OUT <= 0;  //31 / 57 = 0
    16'b00011111_00111010 : OUT <= 0;  //31 / 58 = 0
    16'b00011111_00111011 : OUT <= 0;  //31 / 59 = 0
    16'b00011111_00111100 : OUT <= 0;  //31 / 60 = 0
    16'b00011111_00111101 : OUT <= 0;  //31 / 61 = 0
    16'b00011111_00111110 : OUT <= 0;  //31 / 62 = 0
    16'b00011111_00111111 : OUT <= 0;  //31 / 63 = 0
    16'b00011111_01000000 : OUT <= 0;  //31 / 64 = 0
    16'b00011111_01000001 : OUT <= 0;  //31 / 65 = 0
    16'b00011111_01000010 : OUT <= 0;  //31 / 66 = 0
    16'b00011111_01000011 : OUT <= 0;  //31 / 67 = 0
    16'b00011111_01000100 : OUT <= 0;  //31 / 68 = 0
    16'b00011111_01000101 : OUT <= 0;  //31 / 69 = 0
    16'b00011111_01000110 : OUT <= 0;  //31 / 70 = 0
    16'b00011111_01000111 : OUT <= 0;  //31 / 71 = 0
    16'b00011111_01001000 : OUT <= 0;  //31 / 72 = 0
    16'b00011111_01001001 : OUT <= 0;  //31 / 73 = 0
    16'b00011111_01001010 : OUT <= 0;  //31 / 74 = 0
    16'b00011111_01001011 : OUT <= 0;  //31 / 75 = 0
    16'b00011111_01001100 : OUT <= 0;  //31 / 76 = 0
    16'b00011111_01001101 : OUT <= 0;  //31 / 77 = 0
    16'b00011111_01001110 : OUT <= 0;  //31 / 78 = 0
    16'b00011111_01001111 : OUT <= 0;  //31 / 79 = 0
    16'b00011111_01010000 : OUT <= 0;  //31 / 80 = 0
    16'b00011111_01010001 : OUT <= 0;  //31 / 81 = 0
    16'b00011111_01010010 : OUT <= 0;  //31 / 82 = 0
    16'b00011111_01010011 : OUT <= 0;  //31 / 83 = 0
    16'b00011111_01010100 : OUT <= 0;  //31 / 84 = 0
    16'b00011111_01010101 : OUT <= 0;  //31 / 85 = 0
    16'b00011111_01010110 : OUT <= 0;  //31 / 86 = 0
    16'b00011111_01010111 : OUT <= 0;  //31 / 87 = 0
    16'b00011111_01011000 : OUT <= 0;  //31 / 88 = 0
    16'b00011111_01011001 : OUT <= 0;  //31 / 89 = 0
    16'b00011111_01011010 : OUT <= 0;  //31 / 90 = 0
    16'b00011111_01011011 : OUT <= 0;  //31 / 91 = 0
    16'b00011111_01011100 : OUT <= 0;  //31 / 92 = 0
    16'b00011111_01011101 : OUT <= 0;  //31 / 93 = 0
    16'b00011111_01011110 : OUT <= 0;  //31 / 94 = 0
    16'b00011111_01011111 : OUT <= 0;  //31 / 95 = 0
    16'b00011111_01100000 : OUT <= 0;  //31 / 96 = 0
    16'b00011111_01100001 : OUT <= 0;  //31 / 97 = 0
    16'b00011111_01100010 : OUT <= 0;  //31 / 98 = 0
    16'b00011111_01100011 : OUT <= 0;  //31 / 99 = 0
    16'b00011111_01100100 : OUT <= 0;  //31 / 100 = 0
    16'b00011111_01100101 : OUT <= 0;  //31 / 101 = 0
    16'b00011111_01100110 : OUT <= 0;  //31 / 102 = 0
    16'b00011111_01100111 : OUT <= 0;  //31 / 103 = 0
    16'b00011111_01101000 : OUT <= 0;  //31 / 104 = 0
    16'b00011111_01101001 : OUT <= 0;  //31 / 105 = 0
    16'b00011111_01101010 : OUT <= 0;  //31 / 106 = 0
    16'b00011111_01101011 : OUT <= 0;  //31 / 107 = 0
    16'b00011111_01101100 : OUT <= 0;  //31 / 108 = 0
    16'b00011111_01101101 : OUT <= 0;  //31 / 109 = 0
    16'b00011111_01101110 : OUT <= 0;  //31 / 110 = 0
    16'b00011111_01101111 : OUT <= 0;  //31 / 111 = 0
    16'b00011111_01110000 : OUT <= 0;  //31 / 112 = 0
    16'b00011111_01110001 : OUT <= 0;  //31 / 113 = 0
    16'b00011111_01110010 : OUT <= 0;  //31 / 114 = 0
    16'b00011111_01110011 : OUT <= 0;  //31 / 115 = 0
    16'b00011111_01110100 : OUT <= 0;  //31 / 116 = 0
    16'b00011111_01110101 : OUT <= 0;  //31 / 117 = 0
    16'b00011111_01110110 : OUT <= 0;  //31 / 118 = 0
    16'b00011111_01110111 : OUT <= 0;  //31 / 119 = 0
    16'b00011111_01111000 : OUT <= 0;  //31 / 120 = 0
    16'b00011111_01111001 : OUT <= 0;  //31 / 121 = 0
    16'b00011111_01111010 : OUT <= 0;  //31 / 122 = 0
    16'b00011111_01111011 : OUT <= 0;  //31 / 123 = 0
    16'b00011111_01111100 : OUT <= 0;  //31 / 124 = 0
    16'b00011111_01111101 : OUT <= 0;  //31 / 125 = 0
    16'b00011111_01111110 : OUT <= 0;  //31 / 126 = 0
    16'b00011111_01111111 : OUT <= 0;  //31 / 127 = 0
    16'b00011111_10000000 : OUT <= 0;  //31 / 128 = 0
    16'b00011111_10000001 : OUT <= 0;  //31 / 129 = 0
    16'b00011111_10000010 : OUT <= 0;  //31 / 130 = 0
    16'b00011111_10000011 : OUT <= 0;  //31 / 131 = 0
    16'b00011111_10000100 : OUT <= 0;  //31 / 132 = 0
    16'b00011111_10000101 : OUT <= 0;  //31 / 133 = 0
    16'b00011111_10000110 : OUT <= 0;  //31 / 134 = 0
    16'b00011111_10000111 : OUT <= 0;  //31 / 135 = 0
    16'b00011111_10001000 : OUT <= 0;  //31 / 136 = 0
    16'b00011111_10001001 : OUT <= 0;  //31 / 137 = 0
    16'b00011111_10001010 : OUT <= 0;  //31 / 138 = 0
    16'b00011111_10001011 : OUT <= 0;  //31 / 139 = 0
    16'b00011111_10001100 : OUT <= 0;  //31 / 140 = 0
    16'b00011111_10001101 : OUT <= 0;  //31 / 141 = 0
    16'b00011111_10001110 : OUT <= 0;  //31 / 142 = 0
    16'b00011111_10001111 : OUT <= 0;  //31 / 143 = 0
    16'b00011111_10010000 : OUT <= 0;  //31 / 144 = 0
    16'b00011111_10010001 : OUT <= 0;  //31 / 145 = 0
    16'b00011111_10010010 : OUT <= 0;  //31 / 146 = 0
    16'b00011111_10010011 : OUT <= 0;  //31 / 147 = 0
    16'b00011111_10010100 : OUT <= 0;  //31 / 148 = 0
    16'b00011111_10010101 : OUT <= 0;  //31 / 149 = 0
    16'b00011111_10010110 : OUT <= 0;  //31 / 150 = 0
    16'b00011111_10010111 : OUT <= 0;  //31 / 151 = 0
    16'b00011111_10011000 : OUT <= 0;  //31 / 152 = 0
    16'b00011111_10011001 : OUT <= 0;  //31 / 153 = 0
    16'b00011111_10011010 : OUT <= 0;  //31 / 154 = 0
    16'b00011111_10011011 : OUT <= 0;  //31 / 155 = 0
    16'b00011111_10011100 : OUT <= 0;  //31 / 156 = 0
    16'b00011111_10011101 : OUT <= 0;  //31 / 157 = 0
    16'b00011111_10011110 : OUT <= 0;  //31 / 158 = 0
    16'b00011111_10011111 : OUT <= 0;  //31 / 159 = 0
    16'b00011111_10100000 : OUT <= 0;  //31 / 160 = 0
    16'b00011111_10100001 : OUT <= 0;  //31 / 161 = 0
    16'b00011111_10100010 : OUT <= 0;  //31 / 162 = 0
    16'b00011111_10100011 : OUT <= 0;  //31 / 163 = 0
    16'b00011111_10100100 : OUT <= 0;  //31 / 164 = 0
    16'b00011111_10100101 : OUT <= 0;  //31 / 165 = 0
    16'b00011111_10100110 : OUT <= 0;  //31 / 166 = 0
    16'b00011111_10100111 : OUT <= 0;  //31 / 167 = 0
    16'b00011111_10101000 : OUT <= 0;  //31 / 168 = 0
    16'b00011111_10101001 : OUT <= 0;  //31 / 169 = 0
    16'b00011111_10101010 : OUT <= 0;  //31 / 170 = 0
    16'b00011111_10101011 : OUT <= 0;  //31 / 171 = 0
    16'b00011111_10101100 : OUT <= 0;  //31 / 172 = 0
    16'b00011111_10101101 : OUT <= 0;  //31 / 173 = 0
    16'b00011111_10101110 : OUT <= 0;  //31 / 174 = 0
    16'b00011111_10101111 : OUT <= 0;  //31 / 175 = 0
    16'b00011111_10110000 : OUT <= 0;  //31 / 176 = 0
    16'b00011111_10110001 : OUT <= 0;  //31 / 177 = 0
    16'b00011111_10110010 : OUT <= 0;  //31 / 178 = 0
    16'b00011111_10110011 : OUT <= 0;  //31 / 179 = 0
    16'b00011111_10110100 : OUT <= 0;  //31 / 180 = 0
    16'b00011111_10110101 : OUT <= 0;  //31 / 181 = 0
    16'b00011111_10110110 : OUT <= 0;  //31 / 182 = 0
    16'b00011111_10110111 : OUT <= 0;  //31 / 183 = 0
    16'b00011111_10111000 : OUT <= 0;  //31 / 184 = 0
    16'b00011111_10111001 : OUT <= 0;  //31 / 185 = 0
    16'b00011111_10111010 : OUT <= 0;  //31 / 186 = 0
    16'b00011111_10111011 : OUT <= 0;  //31 / 187 = 0
    16'b00011111_10111100 : OUT <= 0;  //31 / 188 = 0
    16'b00011111_10111101 : OUT <= 0;  //31 / 189 = 0
    16'b00011111_10111110 : OUT <= 0;  //31 / 190 = 0
    16'b00011111_10111111 : OUT <= 0;  //31 / 191 = 0
    16'b00011111_11000000 : OUT <= 0;  //31 / 192 = 0
    16'b00011111_11000001 : OUT <= 0;  //31 / 193 = 0
    16'b00011111_11000010 : OUT <= 0;  //31 / 194 = 0
    16'b00011111_11000011 : OUT <= 0;  //31 / 195 = 0
    16'b00011111_11000100 : OUT <= 0;  //31 / 196 = 0
    16'b00011111_11000101 : OUT <= 0;  //31 / 197 = 0
    16'b00011111_11000110 : OUT <= 0;  //31 / 198 = 0
    16'b00011111_11000111 : OUT <= 0;  //31 / 199 = 0
    16'b00011111_11001000 : OUT <= 0;  //31 / 200 = 0
    16'b00011111_11001001 : OUT <= 0;  //31 / 201 = 0
    16'b00011111_11001010 : OUT <= 0;  //31 / 202 = 0
    16'b00011111_11001011 : OUT <= 0;  //31 / 203 = 0
    16'b00011111_11001100 : OUT <= 0;  //31 / 204 = 0
    16'b00011111_11001101 : OUT <= 0;  //31 / 205 = 0
    16'b00011111_11001110 : OUT <= 0;  //31 / 206 = 0
    16'b00011111_11001111 : OUT <= 0;  //31 / 207 = 0
    16'b00011111_11010000 : OUT <= 0;  //31 / 208 = 0
    16'b00011111_11010001 : OUT <= 0;  //31 / 209 = 0
    16'b00011111_11010010 : OUT <= 0;  //31 / 210 = 0
    16'b00011111_11010011 : OUT <= 0;  //31 / 211 = 0
    16'b00011111_11010100 : OUT <= 0;  //31 / 212 = 0
    16'b00011111_11010101 : OUT <= 0;  //31 / 213 = 0
    16'b00011111_11010110 : OUT <= 0;  //31 / 214 = 0
    16'b00011111_11010111 : OUT <= 0;  //31 / 215 = 0
    16'b00011111_11011000 : OUT <= 0;  //31 / 216 = 0
    16'b00011111_11011001 : OUT <= 0;  //31 / 217 = 0
    16'b00011111_11011010 : OUT <= 0;  //31 / 218 = 0
    16'b00011111_11011011 : OUT <= 0;  //31 / 219 = 0
    16'b00011111_11011100 : OUT <= 0;  //31 / 220 = 0
    16'b00011111_11011101 : OUT <= 0;  //31 / 221 = 0
    16'b00011111_11011110 : OUT <= 0;  //31 / 222 = 0
    16'b00011111_11011111 : OUT <= 0;  //31 / 223 = 0
    16'b00011111_11100000 : OUT <= 0;  //31 / 224 = 0
    16'b00011111_11100001 : OUT <= 0;  //31 / 225 = 0
    16'b00011111_11100010 : OUT <= 0;  //31 / 226 = 0
    16'b00011111_11100011 : OUT <= 0;  //31 / 227 = 0
    16'b00011111_11100100 : OUT <= 0;  //31 / 228 = 0
    16'b00011111_11100101 : OUT <= 0;  //31 / 229 = 0
    16'b00011111_11100110 : OUT <= 0;  //31 / 230 = 0
    16'b00011111_11100111 : OUT <= 0;  //31 / 231 = 0
    16'b00011111_11101000 : OUT <= 0;  //31 / 232 = 0
    16'b00011111_11101001 : OUT <= 0;  //31 / 233 = 0
    16'b00011111_11101010 : OUT <= 0;  //31 / 234 = 0
    16'b00011111_11101011 : OUT <= 0;  //31 / 235 = 0
    16'b00011111_11101100 : OUT <= 0;  //31 / 236 = 0
    16'b00011111_11101101 : OUT <= 0;  //31 / 237 = 0
    16'b00011111_11101110 : OUT <= 0;  //31 / 238 = 0
    16'b00011111_11101111 : OUT <= 0;  //31 / 239 = 0
    16'b00011111_11110000 : OUT <= 0;  //31 / 240 = 0
    16'b00011111_11110001 : OUT <= 0;  //31 / 241 = 0
    16'b00011111_11110010 : OUT <= 0;  //31 / 242 = 0
    16'b00011111_11110011 : OUT <= 0;  //31 / 243 = 0
    16'b00011111_11110100 : OUT <= 0;  //31 / 244 = 0
    16'b00011111_11110101 : OUT <= 0;  //31 / 245 = 0
    16'b00011111_11110110 : OUT <= 0;  //31 / 246 = 0
    16'b00011111_11110111 : OUT <= 0;  //31 / 247 = 0
    16'b00011111_11111000 : OUT <= 0;  //31 / 248 = 0
    16'b00011111_11111001 : OUT <= 0;  //31 / 249 = 0
    16'b00011111_11111010 : OUT <= 0;  //31 / 250 = 0
    16'b00011111_11111011 : OUT <= 0;  //31 / 251 = 0
    16'b00011111_11111100 : OUT <= 0;  //31 / 252 = 0
    16'b00011111_11111101 : OUT <= 0;  //31 / 253 = 0
    16'b00011111_11111110 : OUT <= 0;  //31 / 254 = 0
    16'b00011111_11111111 : OUT <= 0;  //31 / 255 = 0
    16'b00100000_00000000 : OUT <= 0;  //32 / 0 = 0
    16'b00100000_00000001 : OUT <= 32;  //32 / 1 = 32
    16'b00100000_00000010 : OUT <= 16;  //32 / 2 = 16
    16'b00100000_00000011 : OUT <= 10;  //32 / 3 = 10
    16'b00100000_00000100 : OUT <= 8;  //32 / 4 = 8
    16'b00100000_00000101 : OUT <= 6;  //32 / 5 = 6
    16'b00100000_00000110 : OUT <= 5;  //32 / 6 = 5
    16'b00100000_00000111 : OUT <= 4;  //32 / 7 = 4
    16'b00100000_00001000 : OUT <= 4;  //32 / 8 = 4
    16'b00100000_00001001 : OUT <= 3;  //32 / 9 = 3
    16'b00100000_00001010 : OUT <= 3;  //32 / 10 = 3
    16'b00100000_00001011 : OUT <= 2;  //32 / 11 = 2
    16'b00100000_00001100 : OUT <= 2;  //32 / 12 = 2
    16'b00100000_00001101 : OUT <= 2;  //32 / 13 = 2
    16'b00100000_00001110 : OUT <= 2;  //32 / 14 = 2
    16'b00100000_00001111 : OUT <= 2;  //32 / 15 = 2
    16'b00100000_00010000 : OUT <= 2;  //32 / 16 = 2
    16'b00100000_00010001 : OUT <= 1;  //32 / 17 = 1
    16'b00100000_00010010 : OUT <= 1;  //32 / 18 = 1
    16'b00100000_00010011 : OUT <= 1;  //32 / 19 = 1
    16'b00100000_00010100 : OUT <= 1;  //32 / 20 = 1
    16'b00100000_00010101 : OUT <= 1;  //32 / 21 = 1
    16'b00100000_00010110 : OUT <= 1;  //32 / 22 = 1
    16'b00100000_00010111 : OUT <= 1;  //32 / 23 = 1
    16'b00100000_00011000 : OUT <= 1;  //32 / 24 = 1
    16'b00100000_00011001 : OUT <= 1;  //32 / 25 = 1
    16'b00100000_00011010 : OUT <= 1;  //32 / 26 = 1
    16'b00100000_00011011 : OUT <= 1;  //32 / 27 = 1
    16'b00100000_00011100 : OUT <= 1;  //32 / 28 = 1
    16'b00100000_00011101 : OUT <= 1;  //32 / 29 = 1
    16'b00100000_00011110 : OUT <= 1;  //32 / 30 = 1
    16'b00100000_00011111 : OUT <= 1;  //32 / 31 = 1
    16'b00100000_00100000 : OUT <= 1;  //32 / 32 = 1
    16'b00100000_00100001 : OUT <= 0;  //32 / 33 = 0
    16'b00100000_00100010 : OUT <= 0;  //32 / 34 = 0
    16'b00100000_00100011 : OUT <= 0;  //32 / 35 = 0
    16'b00100000_00100100 : OUT <= 0;  //32 / 36 = 0
    16'b00100000_00100101 : OUT <= 0;  //32 / 37 = 0
    16'b00100000_00100110 : OUT <= 0;  //32 / 38 = 0
    16'b00100000_00100111 : OUT <= 0;  //32 / 39 = 0
    16'b00100000_00101000 : OUT <= 0;  //32 / 40 = 0
    16'b00100000_00101001 : OUT <= 0;  //32 / 41 = 0
    16'b00100000_00101010 : OUT <= 0;  //32 / 42 = 0
    16'b00100000_00101011 : OUT <= 0;  //32 / 43 = 0
    16'b00100000_00101100 : OUT <= 0;  //32 / 44 = 0
    16'b00100000_00101101 : OUT <= 0;  //32 / 45 = 0
    16'b00100000_00101110 : OUT <= 0;  //32 / 46 = 0
    16'b00100000_00101111 : OUT <= 0;  //32 / 47 = 0
    16'b00100000_00110000 : OUT <= 0;  //32 / 48 = 0
    16'b00100000_00110001 : OUT <= 0;  //32 / 49 = 0
    16'b00100000_00110010 : OUT <= 0;  //32 / 50 = 0
    16'b00100000_00110011 : OUT <= 0;  //32 / 51 = 0
    16'b00100000_00110100 : OUT <= 0;  //32 / 52 = 0
    16'b00100000_00110101 : OUT <= 0;  //32 / 53 = 0
    16'b00100000_00110110 : OUT <= 0;  //32 / 54 = 0
    16'b00100000_00110111 : OUT <= 0;  //32 / 55 = 0
    16'b00100000_00111000 : OUT <= 0;  //32 / 56 = 0
    16'b00100000_00111001 : OUT <= 0;  //32 / 57 = 0
    16'b00100000_00111010 : OUT <= 0;  //32 / 58 = 0
    16'b00100000_00111011 : OUT <= 0;  //32 / 59 = 0
    16'b00100000_00111100 : OUT <= 0;  //32 / 60 = 0
    16'b00100000_00111101 : OUT <= 0;  //32 / 61 = 0
    16'b00100000_00111110 : OUT <= 0;  //32 / 62 = 0
    16'b00100000_00111111 : OUT <= 0;  //32 / 63 = 0
    16'b00100000_01000000 : OUT <= 0;  //32 / 64 = 0
    16'b00100000_01000001 : OUT <= 0;  //32 / 65 = 0
    16'b00100000_01000010 : OUT <= 0;  //32 / 66 = 0
    16'b00100000_01000011 : OUT <= 0;  //32 / 67 = 0
    16'b00100000_01000100 : OUT <= 0;  //32 / 68 = 0
    16'b00100000_01000101 : OUT <= 0;  //32 / 69 = 0
    16'b00100000_01000110 : OUT <= 0;  //32 / 70 = 0
    16'b00100000_01000111 : OUT <= 0;  //32 / 71 = 0
    16'b00100000_01001000 : OUT <= 0;  //32 / 72 = 0
    16'b00100000_01001001 : OUT <= 0;  //32 / 73 = 0
    16'b00100000_01001010 : OUT <= 0;  //32 / 74 = 0
    16'b00100000_01001011 : OUT <= 0;  //32 / 75 = 0
    16'b00100000_01001100 : OUT <= 0;  //32 / 76 = 0
    16'b00100000_01001101 : OUT <= 0;  //32 / 77 = 0
    16'b00100000_01001110 : OUT <= 0;  //32 / 78 = 0
    16'b00100000_01001111 : OUT <= 0;  //32 / 79 = 0
    16'b00100000_01010000 : OUT <= 0;  //32 / 80 = 0
    16'b00100000_01010001 : OUT <= 0;  //32 / 81 = 0
    16'b00100000_01010010 : OUT <= 0;  //32 / 82 = 0
    16'b00100000_01010011 : OUT <= 0;  //32 / 83 = 0
    16'b00100000_01010100 : OUT <= 0;  //32 / 84 = 0
    16'b00100000_01010101 : OUT <= 0;  //32 / 85 = 0
    16'b00100000_01010110 : OUT <= 0;  //32 / 86 = 0
    16'b00100000_01010111 : OUT <= 0;  //32 / 87 = 0
    16'b00100000_01011000 : OUT <= 0;  //32 / 88 = 0
    16'b00100000_01011001 : OUT <= 0;  //32 / 89 = 0
    16'b00100000_01011010 : OUT <= 0;  //32 / 90 = 0
    16'b00100000_01011011 : OUT <= 0;  //32 / 91 = 0
    16'b00100000_01011100 : OUT <= 0;  //32 / 92 = 0
    16'b00100000_01011101 : OUT <= 0;  //32 / 93 = 0
    16'b00100000_01011110 : OUT <= 0;  //32 / 94 = 0
    16'b00100000_01011111 : OUT <= 0;  //32 / 95 = 0
    16'b00100000_01100000 : OUT <= 0;  //32 / 96 = 0
    16'b00100000_01100001 : OUT <= 0;  //32 / 97 = 0
    16'b00100000_01100010 : OUT <= 0;  //32 / 98 = 0
    16'b00100000_01100011 : OUT <= 0;  //32 / 99 = 0
    16'b00100000_01100100 : OUT <= 0;  //32 / 100 = 0
    16'b00100000_01100101 : OUT <= 0;  //32 / 101 = 0
    16'b00100000_01100110 : OUT <= 0;  //32 / 102 = 0
    16'b00100000_01100111 : OUT <= 0;  //32 / 103 = 0
    16'b00100000_01101000 : OUT <= 0;  //32 / 104 = 0
    16'b00100000_01101001 : OUT <= 0;  //32 / 105 = 0
    16'b00100000_01101010 : OUT <= 0;  //32 / 106 = 0
    16'b00100000_01101011 : OUT <= 0;  //32 / 107 = 0
    16'b00100000_01101100 : OUT <= 0;  //32 / 108 = 0
    16'b00100000_01101101 : OUT <= 0;  //32 / 109 = 0
    16'b00100000_01101110 : OUT <= 0;  //32 / 110 = 0
    16'b00100000_01101111 : OUT <= 0;  //32 / 111 = 0
    16'b00100000_01110000 : OUT <= 0;  //32 / 112 = 0
    16'b00100000_01110001 : OUT <= 0;  //32 / 113 = 0
    16'b00100000_01110010 : OUT <= 0;  //32 / 114 = 0
    16'b00100000_01110011 : OUT <= 0;  //32 / 115 = 0
    16'b00100000_01110100 : OUT <= 0;  //32 / 116 = 0
    16'b00100000_01110101 : OUT <= 0;  //32 / 117 = 0
    16'b00100000_01110110 : OUT <= 0;  //32 / 118 = 0
    16'b00100000_01110111 : OUT <= 0;  //32 / 119 = 0
    16'b00100000_01111000 : OUT <= 0;  //32 / 120 = 0
    16'b00100000_01111001 : OUT <= 0;  //32 / 121 = 0
    16'b00100000_01111010 : OUT <= 0;  //32 / 122 = 0
    16'b00100000_01111011 : OUT <= 0;  //32 / 123 = 0
    16'b00100000_01111100 : OUT <= 0;  //32 / 124 = 0
    16'b00100000_01111101 : OUT <= 0;  //32 / 125 = 0
    16'b00100000_01111110 : OUT <= 0;  //32 / 126 = 0
    16'b00100000_01111111 : OUT <= 0;  //32 / 127 = 0
    16'b00100000_10000000 : OUT <= 0;  //32 / 128 = 0
    16'b00100000_10000001 : OUT <= 0;  //32 / 129 = 0
    16'b00100000_10000010 : OUT <= 0;  //32 / 130 = 0
    16'b00100000_10000011 : OUT <= 0;  //32 / 131 = 0
    16'b00100000_10000100 : OUT <= 0;  //32 / 132 = 0
    16'b00100000_10000101 : OUT <= 0;  //32 / 133 = 0
    16'b00100000_10000110 : OUT <= 0;  //32 / 134 = 0
    16'b00100000_10000111 : OUT <= 0;  //32 / 135 = 0
    16'b00100000_10001000 : OUT <= 0;  //32 / 136 = 0
    16'b00100000_10001001 : OUT <= 0;  //32 / 137 = 0
    16'b00100000_10001010 : OUT <= 0;  //32 / 138 = 0
    16'b00100000_10001011 : OUT <= 0;  //32 / 139 = 0
    16'b00100000_10001100 : OUT <= 0;  //32 / 140 = 0
    16'b00100000_10001101 : OUT <= 0;  //32 / 141 = 0
    16'b00100000_10001110 : OUT <= 0;  //32 / 142 = 0
    16'b00100000_10001111 : OUT <= 0;  //32 / 143 = 0
    16'b00100000_10010000 : OUT <= 0;  //32 / 144 = 0
    16'b00100000_10010001 : OUT <= 0;  //32 / 145 = 0
    16'b00100000_10010010 : OUT <= 0;  //32 / 146 = 0
    16'b00100000_10010011 : OUT <= 0;  //32 / 147 = 0
    16'b00100000_10010100 : OUT <= 0;  //32 / 148 = 0
    16'b00100000_10010101 : OUT <= 0;  //32 / 149 = 0
    16'b00100000_10010110 : OUT <= 0;  //32 / 150 = 0
    16'b00100000_10010111 : OUT <= 0;  //32 / 151 = 0
    16'b00100000_10011000 : OUT <= 0;  //32 / 152 = 0
    16'b00100000_10011001 : OUT <= 0;  //32 / 153 = 0
    16'b00100000_10011010 : OUT <= 0;  //32 / 154 = 0
    16'b00100000_10011011 : OUT <= 0;  //32 / 155 = 0
    16'b00100000_10011100 : OUT <= 0;  //32 / 156 = 0
    16'b00100000_10011101 : OUT <= 0;  //32 / 157 = 0
    16'b00100000_10011110 : OUT <= 0;  //32 / 158 = 0
    16'b00100000_10011111 : OUT <= 0;  //32 / 159 = 0
    16'b00100000_10100000 : OUT <= 0;  //32 / 160 = 0
    16'b00100000_10100001 : OUT <= 0;  //32 / 161 = 0
    16'b00100000_10100010 : OUT <= 0;  //32 / 162 = 0
    16'b00100000_10100011 : OUT <= 0;  //32 / 163 = 0
    16'b00100000_10100100 : OUT <= 0;  //32 / 164 = 0
    16'b00100000_10100101 : OUT <= 0;  //32 / 165 = 0
    16'b00100000_10100110 : OUT <= 0;  //32 / 166 = 0
    16'b00100000_10100111 : OUT <= 0;  //32 / 167 = 0
    16'b00100000_10101000 : OUT <= 0;  //32 / 168 = 0
    16'b00100000_10101001 : OUT <= 0;  //32 / 169 = 0
    16'b00100000_10101010 : OUT <= 0;  //32 / 170 = 0
    16'b00100000_10101011 : OUT <= 0;  //32 / 171 = 0
    16'b00100000_10101100 : OUT <= 0;  //32 / 172 = 0
    16'b00100000_10101101 : OUT <= 0;  //32 / 173 = 0
    16'b00100000_10101110 : OUT <= 0;  //32 / 174 = 0
    16'b00100000_10101111 : OUT <= 0;  //32 / 175 = 0
    16'b00100000_10110000 : OUT <= 0;  //32 / 176 = 0
    16'b00100000_10110001 : OUT <= 0;  //32 / 177 = 0
    16'b00100000_10110010 : OUT <= 0;  //32 / 178 = 0
    16'b00100000_10110011 : OUT <= 0;  //32 / 179 = 0
    16'b00100000_10110100 : OUT <= 0;  //32 / 180 = 0
    16'b00100000_10110101 : OUT <= 0;  //32 / 181 = 0
    16'b00100000_10110110 : OUT <= 0;  //32 / 182 = 0
    16'b00100000_10110111 : OUT <= 0;  //32 / 183 = 0
    16'b00100000_10111000 : OUT <= 0;  //32 / 184 = 0
    16'b00100000_10111001 : OUT <= 0;  //32 / 185 = 0
    16'b00100000_10111010 : OUT <= 0;  //32 / 186 = 0
    16'b00100000_10111011 : OUT <= 0;  //32 / 187 = 0
    16'b00100000_10111100 : OUT <= 0;  //32 / 188 = 0
    16'b00100000_10111101 : OUT <= 0;  //32 / 189 = 0
    16'b00100000_10111110 : OUT <= 0;  //32 / 190 = 0
    16'b00100000_10111111 : OUT <= 0;  //32 / 191 = 0
    16'b00100000_11000000 : OUT <= 0;  //32 / 192 = 0
    16'b00100000_11000001 : OUT <= 0;  //32 / 193 = 0
    16'b00100000_11000010 : OUT <= 0;  //32 / 194 = 0
    16'b00100000_11000011 : OUT <= 0;  //32 / 195 = 0
    16'b00100000_11000100 : OUT <= 0;  //32 / 196 = 0
    16'b00100000_11000101 : OUT <= 0;  //32 / 197 = 0
    16'b00100000_11000110 : OUT <= 0;  //32 / 198 = 0
    16'b00100000_11000111 : OUT <= 0;  //32 / 199 = 0
    16'b00100000_11001000 : OUT <= 0;  //32 / 200 = 0
    16'b00100000_11001001 : OUT <= 0;  //32 / 201 = 0
    16'b00100000_11001010 : OUT <= 0;  //32 / 202 = 0
    16'b00100000_11001011 : OUT <= 0;  //32 / 203 = 0
    16'b00100000_11001100 : OUT <= 0;  //32 / 204 = 0
    16'b00100000_11001101 : OUT <= 0;  //32 / 205 = 0
    16'b00100000_11001110 : OUT <= 0;  //32 / 206 = 0
    16'b00100000_11001111 : OUT <= 0;  //32 / 207 = 0
    16'b00100000_11010000 : OUT <= 0;  //32 / 208 = 0
    16'b00100000_11010001 : OUT <= 0;  //32 / 209 = 0
    16'b00100000_11010010 : OUT <= 0;  //32 / 210 = 0
    16'b00100000_11010011 : OUT <= 0;  //32 / 211 = 0
    16'b00100000_11010100 : OUT <= 0;  //32 / 212 = 0
    16'b00100000_11010101 : OUT <= 0;  //32 / 213 = 0
    16'b00100000_11010110 : OUT <= 0;  //32 / 214 = 0
    16'b00100000_11010111 : OUT <= 0;  //32 / 215 = 0
    16'b00100000_11011000 : OUT <= 0;  //32 / 216 = 0
    16'b00100000_11011001 : OUT <= 0;  //32 / 217 = 0
    16'b00100000_11011010 : OUT <= 0;  //32 / 218 = 0
    16'b00100000_11011011 : OUT <= 0;  //32 / 219 = 0
    16'b00100000_11011100 : OUT <= 0;  //32 / 220 = 0
    16'b00100000_11011101 : OUT <= 0;  //32 / 221 = 0
    16'b00100000_11011110 : OUT <= 0;  //32 / 222 = 0
    16'b00100000_11011111 : OUT <= 0;  //32 / 223 = 0
    16'b00100000_11100000 : OUT <= 0;  //32 / 224 = 0
    16'b00100000_11100001 : OUT <= 0;  //32 / 225 = 0
    16'b00100000_11100010 : OUT <= 0;  //32 / 226 = 0
    16'b00100000_11100011 : OUT <= 0;  //32 / 227 = 0
    16'b00100000_11100100 : OUT <= 0;  //32 / 228 = 0
    16'b00100000_11100101 : OUT <= 0;  //32 / 229 = 0
    16'b00100000_11100110 : OUT <= 0;  //32 / 230 = 0
    16'b00100000_11100111 : OUT <= 0;  //32 / 231 = 0
    16'b00100000_11101000 : OUT <= 0;  //32 / 232 = 0
    16'b00100000_11101001 : OUT <= 0;  //32 / 233 = 0
    16'b00100000_11101010 : OUT <= 0;  //32 / 234 = 0
    16'b00100000_11101011 : OUT <= 0;  //32 / 235 = 0
    16'b00100000_11101100 : OUT <= 0;  //32 / 236 = 0
    16'b00100000_11101101 : OUT <= 0;  //32 / 237 = 0
    16'b00100000_11101110 : OUT <= 0;  //32 / 238 = 0
    16'b00100000_11101111 : OUT <= 0;  //32 / 239 = 0
    16'b00100000_11110000 : OUT <= 0;  //32 / 240 = 0
    16'b00100000_11110001 : OUT <= 0;  //32 / 241 = 0
    16'b00100000_11110010 : OUT <= 0;  //32 / 242 = 0
    16'b00100000_11110011 : OUT <= 0;  //32 / 243 = 0
    16'b00100000_11110100 : OUT <= 0;  //32 / 244 = 0
    16'b00100000_11110101 : OUT <= 0;  //32 / 245 = 0
    16'b00100000_11110110 : OUT <= 0;  //32 / 246 = 0
    16'b00100000_11110111 : OUT <= 0;  //32 / 247 = 0
    16'b00100000_11111000 : OUT <= 0;  //32 / 248 = 0
    16'b00100000_11111001 : OUT <= 0;  //32 / 249 = 0
    16'b00100000_11111010 : OUT <= 0;  //32 / 250 = 0
    16'b00100000_11111011 : OUT <= 0;  //32 / 251 = 0
    16'b00100000_11111100 : OUT <= 0;  //32 / 252 = 0
    16'b00100000_11111101 : OUT <= 0;  //32 / 253 = 0
    16'b00100000_11111110 : OUT <= 0;  //32 / 254 = 0
    16'b00100000_11111111 : OUT <= 0;  //32 / 255 = 0
    16'b00100001_00000000 : OUT <= 0;  //33 / 0 = 0
    16'b00100001_00000001 : OUT <= 33;  //33 / 1 = 33
    16'b00100001_00000010 : OUT <= 16;  //33 / 2 = 16
    16'b00100001_00000011 : OUT <= 11;  //33 / 3 = 11
    16'b00100001_00000100 : OUT <= 8;  //33 / 4 = 8
    16'b00100001_00000101 : OUT <= 6;  //33 / 5 = 6
    16'b00100001_00000110 : OUT <= 5;  //33 / 6 = 5
    16'b00100001_00000111 : OUT <= 4;  //33 / 7 = 4
    16'b00100001_00001000 : OUT <= 4;  //33 / 8 = 4
    16'b00100001_00001001 : OUT <= 3;  //33 / 9 = 3
    16'b00100001_00001010 : OUT <= 3;  //33 / 10 = 3
    16'b00100001_00001011 : OUT <= 3;  //33 / 11 = 3
    16'b00100001_00001100 : OUT <= 2;  //33 / 12 = 2
    16'b00100001_00001101 : OUT <= 2;  //33 / 13 = 2
    16'b00100001_00001110 : OUT <= 2;  //33 / 14 = 2
    16'b00100001_00001111 : OUT <= 2;  //33 / 15 = 2
    16'b00100001_00010000 : OUT <= 2;  //33 / 16 = 2
    16'b00100001_00010001 : OUT <= 1;  //33 / 17 = 1
    16'b00100001_00010010 : OUT <= 1;  //33 / 18 = 1
    16'b00100001_00010011 : OUT <= 1;  //33 / 19 = 1
    16'b00100001_00010100 : OUT <= 1;  //33 / 20 = 1
    16'b00100001_00010101 : OUT <= 1;  //33 / 21 = 1
    16'b00100001_00010110 : OUT <= 1;  //33 / 22 = 1
    16'b00100001_00010111 : OUT <= 1;  //33 / 23 = 1
    16'b00100001_00011000 : OUT <= 1;  //33 / 24 = 1
    16'b00100001_00011001 : OUT <= 1;  //33 / 25 = 1
    16'b00100001_00011010 : OUT <= 1;  //33 / 26 = 1
    16'b00100001_00011011 : OUT <= 1;  //33 / 27 = 1
    16'b00100001_00011100 : OUT <= 1;  //33 / 28 = 1
    16'b00100001_00011101 : OUT <= 1;  //33 / 29 = 1
    16'b00100001_00011110 : OUT <= 1;  //33 / 30 = 1
    16'b00100001_00011111 : OUT <= 1;  //33 / 31 = 1
    16'b00100001_00100000 : OUT <= 1;  //33 / 32 = 1
    16'b00100001_00100001 : OUT <= 1;  //33 / 33 = 1
    16'b00100001_00100010 : OUT <= 0;  //33 / 34 = 0
    16'b00100001_00100011 : OUT <= 0;  //33 / 35 = 0
    16'b00100001_00100100 : OUT <= 0;  //33 / 36 = 0
    16'b00100001_00100101 : OUT <= 0;  //33 / 37 = 0
    16'b00100001_00100110 : OUT <= 0;  //33 / 38 = 0
    16'b00100001_00100111 : OUT <= 0;  //33 / 39 = 0
    16'b00100001_00101000 : OUT <= 0;  //33 / 40 = 0
    16'b00100001_00101001 : OUT <= 0;  //33 / 41 = 0
    16'b00100001_00101010 : OUT <= 0;  //33 / 42 = 0
    16'b00100001_00101011 : OUT <= 0;  //33 / 43 = 0
    16'b00100001_00101100 : OUT <= 0;  //33 / 44 = 0
    16'b00100001_00101101 : OUT <= 0;  //33 / 45 = 0
    16'b00100001_00101110 : OUT <= 0;  //33 / 46 = 0
    16'b00100001_00101111 : OUT <= 0;  //33 / 47 = 0
    16'b00100001_00110000 : OUT <= 0;  //33 / 48 = 0
    16'b00100001_00110001 : OUT <= 0;  //33 / 49 = 0
    16'b00100001_00110010 : OUT <= 0;  //33 / 50 = 0
    16'b00100001_00110011 : OUT <= 0;  //33 / 51 = 0
    16'b00100001_00110100 : OUT <= 0;  //33 / 52 = 0
    16'b00100001_00110101 : OUT <= 0;  //33 / 53 = 0
    16'b00100001_00110110 : OUT <= 0;  //33 / 54 = 0
    16'b00100001_00110111 : OUT <= 0;  //33 / 55 = 0
    16'b00100001_00111000 : OUT <= 0;  //33 / 56 = 0
    16'b00100001_00111001 : OUT <= 0;  //33 / 57 = 0
    16'b00100001_00111010 : OUT <= 0;  //33 / 58 = 0
    16'b00100001_00111011 : OUT <= 0;  //33 / 59 = 0
    16'b00100001_00111100 : OUT <= 0;  //33 / 60 = 0
    16'b00100001_00111101 : OUT <= 0;  //33 / 61 = 0
    16'b00100001_00111110 : OUT <= 0;  //33 / 62 = 0
    16'b00100001_00111111 : OUT <= 0;  //33 / 63 = 0
    16'b00100001_01000000 : OUT <= 0;  //33 / 64 = 0
    16'b00100001_01000001 : OUT <= 0;  //33 / 65 = 0
    16'b00100001_01000010 : OUT <= 0;  //33 / 66 = 0
    16'b00100001_01000011 : OUT <= 0;  //33 / 67 = 0
    16'b00100001_01000100 : OUT <= 0;  //33 / 68 = 0
    16'b00100001_01000101 : OUT <= 0;  //33 / 69 = 0
    16'b00100001_01000110 : OUT <= 0;  //33 / 70 = 0
    16'b00100001_01000111 : OUT <= 0;  //33 / 71 = 0
    16'b00100001_01001000 : OUT <= 0;  //33 / 72 = 0
    16'b00100001_01001001 : OUT <= 0;  //33 / 73 = 0
    16'b00100001_01001010 : OUT <= 0;  //33 / 74 = 0
    16'b00100001_01001011 : OUT <= 0;  //33 / 75 = 0
    16'b00100001_01001100 : OUT <= 0;  //33 / 76 = 0
    16'b00100001_01001101 : OUT <= 0;  //33 / 77 = 0
    16'b00100001_01001110 : OUT <= 0;  //33 / 78 = 0
    16'b00100001_01001111 : OUT <= 0;  //33 / 79 = 0
    16'b00100001_01010000 : OUT <= 0;  //33 / 80 = 0
    16'b00100001_01010001 : OUT <= 0;  //33 / 81 = 0
    16'b00100001_01010010 : OUT <= 0;  //33 / 82 = 0
    16'b00100001_01010011 : OUT <= 0;  //33 / 83 = 0
    16'b00100001_01010100 : OUT <= 0;  //33 / 84 = 0
    16'b00100001_01010101 : OUT <= 0;  //33 / 85 = 0
    16'b00100001_01010110 : OUT <= 0;  //33 / 86 = 0
    16'b00100001_01010111 : OUT <= 0;  //33 / 87 = 0
    16'b00100001_01011000 : OUT <= 0;  //33 / 88 = 0
    16'b00100001_01011001 : OUT <= 0;  //33 / 89 = 0
    16'b00100001_01011010 : OUT <= 0;  //33 / 90 = 0
    16'b00100001_01011011 : OUT <= 0;  //33 / 91 = 0
    16'b00100001_01011100 : OUT <= 0;  //33 / 92 = 0
    16'b00100001_01011101 : OUT <= 0;  //33 / 93 = 0
    16'b00100001_01011110 : OUT <= 0;  //33 / 94 = 0
    16'b00100001_01011111 : OUT <= 0;  //33 / 95 = 0
    16'b00100001_01100000 : OUT <= 0;  //33 / 96 = 0
    16'b00100001_01100001 : OUT <= 0;  //33 / 97 = 0
    16'b00100001_01100010 : OUT <= 0;  //33 / 98 = 0
    16'b00100001_01100011 : OUT <= 0;  //33 / 99 = 0
    16'b00100001_01100100 : OUT <= 0;  //33 / 100 = 0
    16'b00100001_01100101 : OUT <= 0;  //33 / 101 = 0
    16'b00100001_01100110 : OUT <= 0;  //33 / 102 = 0
    16'b00100001_01100111 : OUT <= 0;  //33 / 103 = 0
    16'b00100001_01101000 : OUT <= 0;  //33 / 104 = 0
    16'b00100001_01101001 : OUT <= 0;  //33 / 105 = 0
    16'b00100001_01101010 : OUT <= 0;  //33 / 106 = 0
    16'b00100001_01101011 : OUT <= 0;  //33 / 107 = 0
    16'b00100001_01101100 : OUT <= 0;  //33 / 108 = 0
    16'b00100001_01101101 : OUT <= 0;  //33 / 109 = 0
    16'b00100001_01101110 : OUT <= 0;  //33 / 110 = 0
    16'b00100001_01101111 : OUT <= 0;  //33 / 111 = 0
    16'b00100001_01110000 : OUT <= 0;  //33 / 112 = 0
    16'b00100001_01110001 : OUT <= 0;  //33 / 113 = 0
    16'b00100001_01110010 : OUT <= 0;  //33 / 114 = 0
    16'b00100001_01110011 : OUT <= 0;  //33 / 115 = 0
    16'b00100001_01110100 : OUT <= 0;  //33 / 116 = 0
    16'b00100001_01110101 : OUT <= 0;  //33 / 117 = 0
    16'b00100001_01110110 : OUT <= 0;  //33 / 118 = 0
    16'b00100001_01110111 : OUT <= 0;  //33 / 119 = 0
    16'b00100001_01111000 : OUT <= 0;  //33 / 120 = 0
    16'b00100001_01111001 : OUT <= 0;  //33 / 121 = 0
    16'b00100001_01111010 : OUT <= 0;  //33 / 122 = 0
    16'b00100001_01111011 : OUT <= 0;  //33 / 123 = 0
    16'b00100001_01111100 : OUT <= 0;  //33 / 124 = 0
    16'b00100001_01111101 : OUT <= 0;  //33 / 125 = 0
    16'b00100001_01111110 : OUT <= 0;  //33 / 126 = 0
    16'b00100001_01111111 : OUT <= 0;  //33 / 127 = 0
    16'b00100001_10000000 : OUT <= 0;  //33 / 128 = 0
    16'b00100001_10000001 : OUT <= 0;  //33 / 129 = 0
    16'b00100001_10000010 : OUT <= 0;  //33 / 130 = 0
    16'b00100001_10000011 : OUT <= 0;  //33 / 131 = 0
    16'b00100001_10000100 : OUT <= 0;  //33 / 132 = 0
    16'b00100001_10000101 : OUT <= 0;  //33 / 133 = 0
    16'b00100001_10000110 : OUT <= 0;  //33 / 134 = 0
    16'b00100001_10000111 : OUT <= 0;  //33 / 135 = 0
    16'b00100001_10001000 : OUT <= 0;  //33 / 136 = 0
    16'b00100001_10001001 : OUT <= 0;  //33 / 137 = 0
    16'b00100001_10001010 : OUT <= 0;  //33 / 138 = 0
    16'b00100001_10001011 : OUT <= 0;  //33 / 139 = 0
    16'b00100001_10001100 : OUT <= 0;  //33 / 140 = 0
    16'b00100001_10001101 : OUT <= 0;  //33 / 141 = 0
    16'b00100001_10001110 : OUT <= 0;  //33 / 142 = 0
    16'b00100001_10001111 : OUT <= 0;  //33 / 143 = 0
    16'b00100001_10010000 : OUT <= 0;  //33 / 144 = 0
    16'b00100001_10010001 : OUT <= 0;  //33 / 145 = 0
    16'b00100001_10010010 : OUT <= 0;  //33 / 146 = 0
    16'b00100001_10010011 : OUT <= 0;  //33 / 147 = 0
    16'b00100001_10010100 : OUT <= 0;  //33 / 148 = 0
    16'b00100001_10010101 : OUT <= 0;  //33 / 149 = 0
    16'b00100001_10010110 : OUT <= 0;  //33 / 150 = 0
    16'b00100001_10010111 : OUT <= 0;  //33 / 151 = 0
    16'b00100001_10011000 : OUT <= 0;  //33 / 152 = 0
    16'b00100001_10011001 : OUT <= 0;  //33 / 153 = 0
    16'b00100001_10011010 : OUT <= 0;  //33 / 154 = 0
    16'b00100001_10011011 : OUT <= 0;  //33 / 155 = 0
    16'b00100001_10011100 : OUT <= 0;  //33 / 156 = 0
    16'b00100001_10011101 : OUT <= 0;  //33 / 157 = 0
    16'b00100001_10011110 : OUT <= 0;  //33 / 158 = 0
    16'b00100001_10011111 : OUT <= 0;  //33 / 159 = 0
    16'b00100001_10100000 : OUT <= 0;  //33 / 160 = 0
    16'b00100001_10100001 : OUT <= 0;  //33 / 161 = 0
    16'b00100001_10100010 : OUT <= 0;  //33 / 162 = 0
    16'b00100001_10100011 : OUT <= 0;  //33 / 163 = 0
    16'b00100001_10100100 : OUT <= 0;  //33 / 164 = 0
    16'b00100001_10100101 : OUT <= 0;  //33 / 165 = 0
    16'b00100001_10100110 : OUT <= 0;  //33 / 166 = 0
    16'b00100001_10100111 : OUT <= 0;  //33 / 167 = 0
    16'b00100001_10101000 : OUT <= 0;  //33 / 168 = 0
    16'b00100001_10101001 : OUT <= 0;  //33 / 169 = 0
    16'b00100001_10101010 : OUT <= 0;  //33 / 170 = 0
    16'b00100001_10101011 : OUT <= 0;  //33 / 171 = 0
    16'b00100001_10101100 : OUT <= 0;  //33 / 172 = 0
    16'b00100001_10101101 : OUT <= 0;  //33 / 173 = 0
    16'b00100001_10101110 : OUT <= 0;  //33 / 174 = 0
    16'b00100001_10101111 : OUT <= 0;  //33 / 175 = 0
    16'b00100001_10110000 : OUT <= 0;  //33 / 176 = 0
    16'b00100001_10110001 : OUT <= 0;  //33 / 177 = 0
    16'b00100001_10110010 : OUT <= 0;  //33 / 178 = 0
    16'b00100001_10110011 : OUT <= 0;  //33 / 179 = 0
    16'b00100001_10110100 : OUT <= 0;  //33 / 180 = 0
    16'b00100001_10110101 : OUT <= 0;  //33 / 181 = 0
    16'b00100001_10110110 : OUT <= 0;  //33 / 182 = 0
    16'b00100001_10110111 : OUT <= 0;  //33 / 183 = 0
    16'b00100001_10111000 : OUT <= 0;  //33 / 184 = 0
    16'b00100001_10111001 : OUT <= 0;  //33 / 185 = 0
    16'b00100001_10111010 : OUT <= 0;  //33 / 186 = 0
    16'b00100001_10111011 : OUT <= 0;  //33 / 187 = 0
    16'b00100001_10111100 : OUT <= 0;  //33 / 188 = 0
    16'b00100001_10111101 : OUT <= 0;  //33 / 189 = 0
    16'b00100001_10111110 : OUT <= 0;  //33 / 190 = 0
    16'b00100001_10111111 : OUT <= 0;  //33 / 191 = 0
    16'b00100001_11000000 : OUT <= 0;  //33 / 192 = 0
    16'b00100001_11000001 : OUT <= 0;  //33 / 193 = 0
    16'b00100001_11000010 : OUT <= 0;  //33 / 194 = 0
    16'b00100001_11000011 : OUT <= 0;  //33 / 195 = 0
    16'b00100001_11000100 : OUT <= 0;  //33 / 196 = 0
    16'b00100001_11000101 : OUT <= 0;  //33 / 197 = 0
    16'b00100001_11000110 : OUT <= 0;  //33 / 198 = 0
    16'b00100001_11000111 : OUT <= 0;  //33 / 199 = 0
    16'b00100001_11001000 : OUT <= 0;  //33 / 200 = 0
    16'b00100001_11001001 : OUT <= 0;  //33 / 201 = 0
    16'b00100001_11001010 : OUT <= 0;  //33 / 202 = 0
    16'b00100001_11001011 : OUT <= 0;  //33 / 203 = 0
    16'b00100001_11001100 : OUT <= 0;  //33 / 204 = 0
    16'b00100001_11001101 : OUT <= 0;  //33 / 205 = 0
    16'b00100001_11001110 : OUT <= 0;  //33 / 206 = 0
    16'b00100001_11001111 : OUT <= 0;  //33 / 207 = 0
    16'b00100001_11010000 : OUT <= 0;  //33 / 208 = 0
    16'b00100001_11010001 : OUT <= 0;  //33 / 209 = 0
    16'b00100001_11010010 : OUT <= 0;  //33 / 210 = 0
    16'b00100001_11010011 : OUT <= 0;  //33 / 211 = 0
    16'b00100001_11010100 : OUT <= 0;  //33 / 212 = 0
    16'b00100001_11010101 : OUT <= 0;  //33 / 213 = 0
    16'b00100001_11010110 : OUT <= 0;  //33 / 214 = 0
    16'b00100001_11010111 : OUT <= 0;  //33 / 215 = 0
    16'b00100001_11011000 : OUT <= 0;  //33 / 216 = 0
    16'b00100001_11011001 : OUT <= 0;  //33 / 217 = 0
    16'b00100001_11011010 : OUT <= 0;  //33 / 218 = 0
    16'b00100001_11011011 : OUT <= 0;  //33 / 219 = 0
    16'b00100001_11011100 : OUT <= 0;  //33 / 220 = 0
    16'b00100001_11011101 : OUT <= 0;  //33 / 221 = 0
    16'b00100001_11011110 : OUT <= 0;  //33 / 222 = 0
    16'b00100001_11011111 : OUT <= 0;  //33 / 223 = 0
    16'b00100001_11100000 : OUT <= 0;  //33 / 224 = 0
    16'b00100001_11100001 : OUT <= 0;  //33 / 225 = 0
    16'b00100001_11100010 : OUT <= 0;  //33 / 226 = 0
    16'b00100001_11100011 : OUT <= 0;  //33 / 227 = 0
    16'b00100001_11100100 : OUT <= 0;  //33 / 228 = 0
    16'b00100001_11100101 : OUT <= 0;  //33 / 229 = 0
    16'b00100001_11100110 : OUT <= 0;  //33 / 230 = 0
    16'b00100001_11100111 : OUT <= 0;  //33 / 231 = 0
    16'b00100001_11101000 : OUT <= 0;  //33 / 232 = 0
    16'b00100001_11101001 : OUT <= 0;  //33 / 233 = 0
    16'b00100001_11101010 : OUT <= 0;  //33 / 234 = 0
    16'b00100001_11101011 : OUT <= 0;  //33 / 235 = 0
    16'b00100001_11101100 : OUT <= 0;  //33 / 236 = 0
    16'b00100001_11101101 : OUT <= 0;  //33 / 237 = 0
    16'b00100001_11101110 : OUT <= 0;  //33 / 238 = 0
    16'b00100001_11101111 : OUT <= 0;  //33 / 239 = 0
    16'b00100001_11110000 : OUT <= 0;  //33 / 240 = 0
    16'b00100001_11110001 : OUT <= 0;  //33 / 241 = 0
    16'b00100001_11110010 : OUT <= 0;  //33 / 242 = 0
    16'b00100001_11110011 : OUT <= 0;  //33 / 243 = 0
    16'b00100001_11110100 : OUT <= 0;  //33 / 244 = 0
    16'b00100001_11110101 : OUT <= 0;  //33 / 245 = 0
    16'b00100001_11110110 : OUT <= 0;  //33 / 246 = 0
    16'b00100001_11110111 : OUT <= 0;  //33 / 247 = 0
    16'b00100001_11111000 : OUT <= 0;  //33 / 248 = 0
    16'b00100001_11111001 : OUT <= 0;  //33 / 249 = 0
    16'b00100001_11111010 : OUT <= 0;  //33 / 250 = 0
    16'b00100001_11111011 : OUT <= 0;  //33 / 251 = 0
    16'b00100001_11111100 : OUT <= 0;  //33 / 252 = 0
    16'b00100001_11111101 : OUT <= 0;  //33 / 253 = 0
    16'b00100001_11111110 : OUT <= 0;  //33 / 254 = 0
    16'b00100001_11111111 : OUT <= 0;  //33 / 255 = 0
    16'b00100010_00000000 : OUT <= 0;  //34 / 0 = 0
    16'b00100010_00000001 : OUT <= 34;  //34 / 1 = 34
    16'b00100010_00000010 : OUT <= 17;  //34 / 2 = 17
    16'b00100010_00000011 : OUT <= 11;  //34 / 3 = 11
    16'b00100010_00000100 : OUT <= 8;  //34 / 4 = 8
    16'b00100010_00000101 : OUT <= 6;  //34 / 5 = 6
    16'b00100010_00000110 : OUT <= 5;  //34 / 6 = 5
    16'b00100010_00000111 : OUT <= 4;  //34 / 7 = 4
    16'b00100010_00001000 : OUT <= 4;  //34 / 8 = 4
    16'b00100010_00001001 : OUT <= 3;  //34 / 9 = 3
    16'b00100010_00001010 : OUT <= 3;  //34 / 10 = 3
    16'b00100010_00001011 : OUT <= 3;  //34 / 11 = 3
    16'b00100010_00001100 : OUT <= 2;  //34 / 12 = 2
    16'b00100010_00001101 : OUT <= 2;  //34 / 13 = 2
    16'b00100010_00001110 : OUT <= 2;  //34 / 14 = 2
    16'b00100010_00001111 : OUT <= 2;  //34 / 15 = 2
    16'b00100010_00010000 : OUT <= 2;  //34 / 16 = 2
    16'b00100010_00010001 : OUT <= 2;  //34 / 17 = 2
    16'b00100010_00010010 : OUT <= 1;  //34 / 18 = 1
    16'b00100010_00010011 : OUT <= 1;  //34 / 19 = 1
    16'b00100010_00010100 : OUT <= 1;  //34 / 20 = 1
    16'b00100010_00010101 : OUT <= 1;  //34 / 21 = 1
    16'b00100010_00010110 : OUT <= 1;  //34 / 22 = 1
    16'b00100010_00010111 : OUT <= 1;  //34 / 23 = 1
    16'b00100010_00011000 : OUT <= 1;  //34 / 24 = 1
    16'b00100010_00011001 : OUT <= 1;  //34 / 25 = 1
    16'b00100010_00011010 : OUT <= 1;  //34 / 26 = 1
    16'b00100010_00011011 : OUT <= 1;  //34 / 27 = 1
    16'b00100010_00011100 : OUT <= 1;  //34 / 28 = 1
    16'b00100010_00011101 : OUT <= 1;  //34 / 29 = 1
    16'b00100010_00011110 : OUT <= 1;  //34 / 30 = 1
    16'b00100010_00011111 : OUT <= 1;  //34 / 31 = 1
    16'b00100010_00100000 : OUT <= 1;  //34 / 32 = 1
    16'b00100010_00100001 : OUT <= 1;  //34 / 33 = 1
    16'b00100010_00100010 : OUT <= 1;  //34 / 34 = 1
    16'b00100010_00100011 : OUT <= 0;  //34 / 35 = 0
    16'b00100010_00100100 : OUT <= 0;  //34 / 36 = 0
    16'b00100010_00100101 : OUT <= 0;  //34 / 37 = 0
    16'b00100010_00100110 : OUT <= 0;  //34 / 38 = 0
    16'b00100010_00100111 : OUT <= 0;  //34 / 39 = 0
    16'b00100010_00101000 : OUT <= 0;  //34 / 40 = 0
    16'b00100010_00101001 : OUT <= 0;  //34 / 41 = 0
    16'b00100010_00101010 : OUT <= 0;  //34 / 42 = 0
    16'b00100010_00101011 : OUT <= 0;  //34 / 43 = 0
    16'b00100010_00101100 : OUT <= 0;  //34 / 44 = 0
    16'b00100010_00101101 : OUT <= 0;  //34 / 45 = 0
    16'b00100010_00101110 : OUT <= 0;  //34 / 46 = 0
    16'b00100010_00101111 : OUT <= 0;  //34 / 47 = 0
    16'b00100010_00110000 : OUT <= 0;  //34 / 48 = 0
    16'b00100010_00110001 : OUT <= 0;  //34 / 49 = 0
    16'b00100010_00110010 : OUT <= 0;  //34 / 50 = 0
    16'b00100010_00110011 : OUT <= 0;  //34 / 51 = 0
    16'b00100010_00110100 : OUT <= 0;  //34 / 52 = 0
    16'b00100010_00110101 : OUT <= 0;  //34 / 53 = 0
    16'b00100010_00110110 : OUT <= 0;  //34 / 54 = 0
    16'b00100010_00110111 : OUT <= 0;  //34 / 55 = 0
    16'b00100010_00111000 : OUT <= 0;  //34 / 56 = 0
    16'b00100010_00111001 : OUT <= 0;  //34 / 57 = 0
    16'b00100010_00111010 : OUT <= 0;  //34 / 58 = 0
    16'b00100010_00111011 : OUT <= 0;  //34 / 59 = 0
    16'b00100010_00111100 : OUT <= 0;  //34 / 60 = 0
    16'b00100010_00111101 : OUT <= 0;  //34 / 61 = 0
    16'b00100010_00111110 : OUT <= 0;  //34 / 62 = 0
    16'b00100010_00111111 : OUT <= 0;  //34 / 63 = 0
    16'b00100010_01000000 : OUT <= 0;  //34 / 64 = 0
    16'b00100010_01000001 : OUT <= 0;  //34 / 65 = 0
    16'b00100010_01000010 : OUT <= 0;  //34 / 66 = 0
    16'b00100010_01000011 : OUT <= 0;  //34 / 67 = 0
    16'b00100010_01000100 : OUT <= 0;  //34 / 68 = 0
    16'b00100010_01000101 : OUT <= 0;  //34 / 69 = 0
    16'b00100010_01000110 : OUT <= 0;  //34 / 70 = 0
    16'b00100010_01000111 : OUT <= 0;  //34 / 71 = 0
    16'b00100010_01001000 : OUT <= 0;  //34 / 72 = 0
    16'b00100010_01001001 : OUT <= 0;  //34 / 73 = 0
    16'b00100010_01001010 : OUT <= 0;  //34 / 74 = 0
    16'b00100010_01001011 : OUT <= 0;  //34 / 75 = 0
    16'b00100010_01001100 : OUT <= 0;  //34 / 76 = 0
    16'b00100010_01001101 : OUT <= 0;  //34 / 77 = 0
    16'b00100010_01001110 : OUT <= 0;  //34 / 78 = 0
    16'b00100010_01001111 : OUT <= 0;  //34 / 79 = 0
    16'b00100010_01010000 : OUT <= 0;  //34 / 80 = 0
    16'b00100010_01010001 : OUT <= 0;  //34 / 81 = 0
    16'b00100010_01010010 : OUT <= 0;  //34 / 82 = 0
    16'b00100010_01010011 : OUT <= 0;  //34 / 83 = 0
    16'b00100010_01010100 : OUT <= 0;  //34 / 84 = 0
    16'b00100010_01010101 : OUT <= 0;  //34 / 85 = 0
    16'b00100010_01010110 : OUT <= 0;  //34 / 86 = 0
    16'b00100010_01010111 : OUT <= 0;  //34 / 87 = 0
    16'b00100010_01011000 : OUT <= 0;  //34 / 88 = 0
    16'b00100010_01011001 : OUT <= 0;  //34 / 89 = 0
    16'b00100010_01011010 : OUT <= 0;  //34 / 90 = 0
    16'b00100010_01011011 : OUT <= 0;  //34 / 91 = 0
    16'b00100010_01011100 : OUT <= 0;  //34 / 92 = 0
    16'b00100010_01011101 : OUT <= 0;  //34 / 93 = 0
    16'b00100010_01011110 : OUT <= 0;  //34 / 94 = 0
    16'b00100010_01011111 : OUT <= 0;  //34 / 95 = 0
    16'b00100010_01100000 : OUT <= 0;  //34 / 96 = 0
    16'b00100010_01100001 : OUT <= 0;  //34 / 97 = 0
    16'b00100010_01100010 : OUT <= 0;  //34 / 98 = 0
    16'b00100010_01100011 : OUT <= 0;  //34 / 99 = 0
    16'b00100010_01100100 : OUT <= 0;  //34 / 100 = 0
    16'b00100010_01100101 : OUT <= 0;  //34 / 101 = 0
    16'b00100010_01100110 : OUT <= 0;  //34 / 102 = 0
    16'b00100010_01100111 : OUT <= 0;  //34 / 103 = 0
    16'b00100010_01101000 : OUT <= 0;  //34 / 104 = 0
    16'b00100010_01101001 : OUT <= 0;  //34 / 105 = 0
    16'b00100010_01101010 : OUT <= 0;  //34 / 106 = 0
    16'b00100010_01101011 : OUT <= 0;  //34 / 107 = 0
    16'b00100010_01101100 : OUT <= 0;  //34 / 108 = 0
    16'b00100010_01101101 : OUT <= 0;  //34 / 109 = 0
    16'b00100010_01101110 : OUT <= 0;  //34 / 110 = 0
    16'b00100010_01101111 : OUT <= 0;  //34 / 111 = 0
    16'b00100010_01110000 : OUT <= 0;  //34 / 112 = 0
    16'b00100010_01110001 : OUT <= 0;  //34 / 113 = 0
    16'b00100010_01110010 : OUT <= 0;  //34 / 114 = 0
    16'b00100010_01110011 : OUT <= 0;  //34 / 115 = 0
    16'b00100010_01110100 : OUT <= 0;  //34 / 116 = 0
    16'b00100010_01110101 : OUT <= 0;  //34 / 117 = 0
    16'b00100010_01110110 : OUT <= 0;  //34 / 118 = 0
    16'b00100010_01110111 : OUT <= 0;  //34 / 119 = 0
    16'b00100010_01111000 : OUT <= 0;  //34 / 120 = 0
    16'b00100010_01111001 : OUT <= 0;  //34 / 121 = 0
    16'b00100010_01111010 : OUT <= 0;  //34 / 122 = 0
    16'b00100010_01111011 : OUT <= 0;  //34 / 123 = 0
    16'b00100010_01111100 : OUT <= 0;  //34 / 124 = 0
    16'b00100010_01111101 : OUT <= 0;  //34 / 125 = 0
    16'b00100010_01111110 : OUT <= 0;  //34 / 126 = 0
    16'b00100010_01111111 : OUT <= 0;  //34 / 127 = 0
    16'b00100010_10000000 : OUT <= 0;  //34 / 128 = 0
    16'b00100010_10000001 : OUT <= 0;  //34 / 129 = 0
    16'b00100010_10000010 : OUT <= 0;  //34 / 130 = 0
    16'b00100010_10000011 : OUT <= 0;  //34 / 131 = 0
    16'b00100010_10000100 : OUT <= 0;  //34 / 132 = 0
    16'b00100010_10000101 : OUT <= 0;  //34 / 133 = 0
    16'b00100010_10000110 : OUT <= 0;  //34 / 134 = 0
    16'b00100010_10000111 : OUT <= 0;  //34 / 135 = 0
    16'b00100010_10001000 : OUT <= 0;  //34 / 136 = 0
    16'b00100010_10001001 : OUT <= 0;  //34 / 137 = 0
    16'b00100010_10001010 : OUT <= 0;  //34 / 138 = 0
    16'b00100010_10001011 : OUT <= 0;  //34 / 139 = 0
    16'b00100010_10001100 : OUT <= 0;  //34 / 140 = 0
    16'b00100010_10001101 : OUT <= 0;  //34 / 141 = 0
    16'b00100010_10001110 : OUT <= 0;  //34 / 142 = 0
    16'b00100010_10001111 : OUT <= 0;  //34 / 143 = 0
    16'b00100010_10010000 : OUT <= 0;  //34 / 144 = 0
    16'b00100010_10010001 : OUT <= 0;  //34 / 145 = 0
    16'b00100010_10010010 : OUT <= 0;  //34 / 146 = 0
    16'b00100010_10010011 : OUT <= 0;  //34 / 147 = 0
    16'b00100010_10010100 : OUT <= 0;  //34 / 148 = 0
    16'b00100010_10010101 : OUT <= 0;  //34 / 149 = 0
    16'b00100010_10010110 : OUT <= 0;  //34 / 150 = 0
    16'b00100010_10010111 : OUT <= 0;  //34 / 151 = 0
    16'b00100010_10011000 : OUT <= 0;  //34 / 152 = 0
    16'b00100010_10011001 : OUT <= 0;  //34 / 153 = 0
    16'b00100010_10011010 : OUT <= 0;  //34 / 154 = 0
    16'b00100010_10011011 : OUT <= 0;  //34 / 155 = 0
    16'b00100010_10011100 : OUT <= 0;  //34 / 156 = 0
    16'b00100010_10011101 : OUT <= 0;  //34 / 157 = 0
    16'b00100010_10011110 : OUT <= 0;  //34 / 158 = 0
    16'b00100010_10011111 : OUT <= 0;  //34 / 159 = 0
    16'b00100010_10100000 : OUT <= 0;  //34 / 160 = 0
    16'b00100010_10100001 : OUT <= 0;  //34 / 161 = 0
    16'b00100010_10100010 : OUT <= 0;  //34 / 162 = 0
    16'b00100010_10100011 : OUT <= 0;  //34 / 163 = 0
    16'b00100010_10100100 : OUT <= 0;  //34 / 164 = 0
    16'b00100010_10100101 : OUT <= 0;  //34 / 165 = 0
    16'b00100010_10100110 : OUT <= 0;  //34 / 166 = 0
    16'b00100010_10100111 : OUT <= 0;  //34 / 167 = 0
    16'b00100010_10101000 : OUT <= 0;  //34 / 168 = 0
    16'b00100010_10101001 : OUT <= 0;  //34 / 169 = 0
    16'b00100010_10101010 : OUT <= 0;  //34 / 170 = 0
    16'b00100010_10101011 : OUT <= 0;  //34 / 171 = 0
    16'b00100010_10101100 : OUT <= 0;  //34 / 172 = 0
    16'b00100010_10101101 : OUT <= 0;  //34 / 173 = 0
    16'b00100010_10101110 : OUT <= 0;  //34 / 174 = 0
    16'b00100010_10101111 : OUT <= 0;  //34 / 175 = 0
    16'b00100010_10110000 : OUT <= 0;  //34 / 176 = 0
    16'b00100010_10110001 : OUT <= 0;  //34 / 177 = 0
    16'b00100010_10110010 : OUT <= 0;  //34 / 178 = 0
    16'b00100010_10110011 : OUT <= 0;  //34 / 179 = 0
    16'b00100010_10110100 : OUT <= 0;  //34 / 180 = 0
    16'b00100010_10110101 : OUT <= 0;  //34 / 181 = 0
    16'b00100010_10110110 : OUT <= 0;  //34 / 182 = 0
    16'b00100010_10110111 : OUT <= 0;  //34 / 183 = 0
    16'b00100010_10111000 : OUT <= 0;  //34 / 184 = 0
    16'b00100010_10111001 : OUT <= 0;  //34 / 185 = 0
    16'b00100010_10111010 : OUT <= 0;  //34 / 186 = 0
    16'b00100010_10111011 : OUT <= 0;  //34 / 187 = 0
    16'b00100010_10111100 : OUT <= 0;  //34 / 188 = 0
    16'b00100010_10111101 : OUT <= 0;  //34 / 189 = 0
    16'b00100010_10111110 : OUT <= 0;  //34 / 190 = 0
    16'b00100010_10111111 : OUT <= 0;  //34 / 191 = 0
    16'b00100010_11000000 : OUT <= 0;  //34 / 192 = 0
    16'b00100010_11000001 : OUT <= 0;  //34 / 193 = 0
    16'b00100010_11000010 : OUT <= 0;  //34 / 194 = 0
    16'b00100010_11000011 : OUT <= 0;  //34 / 195 = 0
    16'b00100010_11000100 : OUT <= 0;  //34 / 196 = 0
    16'b00100010_11000101 : OUT <= 0;  //34 / 197 = 0
    16'b00100010_11000110 : OUT <= 0;  //34 / 198 = 0
    16'b00100010_11000111 : OUT <= 0;  //34 / 199 = 0
    16'b00100010_11001000 : OUT <= 0;  //34 / 200 = 0
    16'b00100010_11001001 : OUT <= 0;  //34 / 201 = 0
    16'b00100010_11001010 : OUT <= 0;  //34 / 202 = 0
    16'b00100010_11001011 : OUT <= 0;  //34 / 203 = 0
    16'b00100010_11001100 : OUT <= 0;  //34 / 204 = 0
    16'b00100010_11001101 : OUT <= 0;  //34 / 205 = 0
    16'b00100010_11001110 : OUT <= 0;  //34 / 206 = 0
    16'b00100010_11001111 : OUT <= 0;  //34 / 207 = 0
    16'b00100010_11010000 : OUT <= 0;  //34 / 208 = 0
    16'b00100010_11010001 : OUT <= 0;  //34 / 209 = 0
    16'b00100010_11010010 : OUT <= 0;  //34 / 210 = 0
    16'b00100010_11010011 : OUT <= 0;  //34 / 211 = 0
    16'b00100010_11010100 : OUT <= 0;  //34 / 212 = 0
    16'b00100010_11010101 : OUT <= 0;  //34 / 213 = 0
    16'b00100010_11010110 : OUT <= 0;  //34 / 214 = 0
    16'b00100010_11010111 : OUT <= 0;  //34 / 215 = 0
    16'b00100010_11011000 : OUT <= 0;  //34 / 216 = 0
    16'b00100010_11011001 : OUT <= 0;  //34 / 217 = 0
    16'b00100010_11011010 : OUT <= 0;  //34 / 218 = 0
    16'b00100010_11011011 : OUT <= 0;  //34 / 219 = 0
    16'b00100010_11011100 : OUT <= 0;  //34 / 220 = 0
    16'b00100010_11011101 : OUT <= 0;  //34 / 221 = 0
    16'b00100010_11011110 : OUT <= 0;  //34 / 222 = 0
    16'b00100010_11011111 : OUT <= 0;  //34 / 223 = 0
    16'b00100010_11100000 : OUT <= 0;  //34 / 224 = 0
    16'b00100010_11100001 : OUT <= 0;  //34 / 225 = 0
    16'b00100010_11100010 : OUT <= 0;  //34 / 226 = 0
    16'b00100010_11100011 : OUT <= 0;  //34 / 227 = 0
    16'b00100010_11100100 : OUT <= 0;  //34 / 228 = 0
    16'b00100010_11100101 : OUT <= 0;  //34 / 229 = 0
    16'b00100010_11100110 : OUT <= 0;  //34 / 230 = 0
    16'b00100010_11100111 : OUT <= 0;  //34 / 231 = 0
    16'b00100010_11101000 : OUT <= 0;  //34 / 232 = 0
    16'b00100010_11101001 : OUT <= 0;  //34 / 233 = 0
    16'b00100010_11101010 : OUT <= 0;  //34 / 234 = 0
    16'b00100010_11101011 : OUT <= 0;  //34 / 235 = 0
    16'b00100010_11101100 : OUT <= 0;  //34 / 236 = 0
    16'b00100010_11101101 : OUT <= 0;  //34 / 237 = 0
    16'b00100010_11101110 : OUT <= 0;  //34 / 238 = 0
    16'b00100010_11101111 : OUT <= 0;  //34 / 239 = 0
    16'b00100010_11110000 : OUT <= 0;  //34 / 240 = 0
    16'b00100010_11110001 : OUT <= 0;  //34 / 241 = 0
    16'b00100010_11110010 : OUT <= 0;  //34 / 242 = 0
    16'b00100010_11110011 : OUT <= 0;  //34 / 243 = 0
    16'b00100010_11110100 : OUT <= 0;  //34 / 244 = 0
    16'b00100010_11110101 : OUT <= 0;  //34 / 245 = 0
    16'b00100010_11110110 : OUT <= 0;  //34 / 246 = 0
    16'b00100010_11110111 : OUT <= 0;  //34 / 247 = 0
    16'b00100010_11111000 : OUT <= 0;  //34 / 248 = 0
    16'b00100010_11111001 : OUT <= 0;  //34 / 249 = 0
    16'b00100010_11111010 : OUT <= 0;  //34 / 250 = 0
    16'b00100010_11111011 : OUT <= 0;  //34 / 251 = 0
    16'b00100010_11111100 : OUT <= 0;  //34 / 252 = 0
    16'b00100010_11111101 : OUT <= 0;  //34 / 253 = 0
    16'b00100010_11111110 : OUT <= 0;  //34 / 254 = 0
    16'b00100010_11111111 : OUT <= 0;  //34 / 255 = 0
    16'b00100011_00000000 : OUT <= 0;  //35 / 0 = 0
    16'b00100011_00000001 : OUT <= 35;  //35 / 1 = 35
    16'b00100011_00000010 : OUT <= 17;  //35 / 2 = 17
    16'b00100011_00000011 : OUT <= 11;  //35 / 3 = 11
    16'b00100011_00000100 : OUT <= 8;  //35 / 4 = 8
    16'b00100011_00000101 : OUT <= 7;  //35 / 5 = 7
    16'b00100011_00000110 : OUT <= 5;  //35 / 6 = 5
    16'b00100011_00000111 : OUT <= 5;  //35 / 7 = 5
    16'b00100011_00001000 : OUT <= 4;  //35 / 8 = 4
    16'b00100011_00001001 : OUT <= 3;  //35 / 9 = 3
    16'b00100011_00001010 : OUT <= 3;  //35 / 10 = 3
    16'b00100011_00001011 : OUT <= 3;  //35 / 11 = 3
    16'b00100011_00001100 : OUT <= 2;  //35 / 12 = 2
    16'b00100011_00001101 : OUT <= 2;  //35 / 13 = 2
    16'b00100011_00001110 : OUT <= 2;  //35 / 14 = 2
    16'b00100011_00001111 : OUT <= 2;  //35 / 15 = 2
    16'b00100011_00010000 : OUT <= 2;  //35 / 16 = 2
    16'b00100011_00010001 : OUT <= 2;  //35 / 17 = 2
    16'b00100011_00010010 : OUT <= 1;  //35 / 18 = 1
    16'b00100011_00010011 : OUT <= 1;  //35 / 19 = 1
    16'b00100011_00010100 : OUT <= 1;  //35 / 20 = 1
    16'b00100011_00010101 : OUT <= 1;  //35 / 21 = 1
    16'b00100011_00010110 : OUT <= 1;  //35 / 22 = 1
    16'b00100011_00010111 : OUT <= 1;  //35 / 23 = 1
    16'b00100011_00011000 : OUT <= 1;  //35 / 24 = 1
    16'b00100011_00011001 : OUT <= 1;  //35 / 25 = 1
    16'b00100011_00011010 : OUT <= 1;  //35 / 26 = 1
    16'b00100011_00011011 : OUT <= 1;  //35 / 27 = 1
    16'b00100011_00011100 : OUT <= 1;  //35 / 28 = 1
    16'b00100011_00011101 : OUT <= 1;  //35 / 29 = 1
    16'b00100011_00011110 : OUT <= 1;  //35 / 30 = 1
    16'b00100011_00011111 : OUT <= 1;  //35 / 31 = 1
    16'b00100011_00100000 : OUT <= 1;  //35 / 32 = 1
    16'b00100011_00100001 : OUT <= 1;  //35 / 33 = 1
    16'b00100011_00100010 : OUT <= 1;  //35 / 34 = 1
    16'b00100011_00100011 : OUT <= 1;  //35 / 35 = 1
    16'b00100011_00100100 : OUT <= 0;  //35 / 36 = 0
    16'b00100011_00100101 : OUT <= 0;  //35 / 37 = 0
    16'b00100011_00100110 : OUT <= 0;  //35 / 38 = 0
    16'b00100011_00100111 : OUT <= 0;  //35 / 39 = 0
    16'b00100011_00101000 : OUT <= 0;  //35 / 40 = 0
    16'b00100011_00101001 : OUT <= 0;  //35 / 41 = 0
    16'b00100011_00101010 : OUT <= 0;  //35 / 42 = 0
    16'b00100011_00101011 : OUT <= 0;  //35 / 43 = 0
    16'b00100011_00101100 : OUT <= 0;  //35 / 44 = 0
    16'b00100011_00101101 : OUT <= 0;  //35 / 45 = 0
    16'b00100011_00101110 : OUT <= 0;  //35 / 46 = 0
    16'b00100011_00101111 : OUT <= 0;  //35 / 47 = 0
    16'b00100011_00110000 : OUT <= 0;  //35 / 48 = 0
    16'b00100011_00110001 : OUT <= 0;  //35 / 49 = 0
    16'b00100011_00110010 : OUT <= 0;  //35 / 50 = 0
    16'b00100011_00110011 : OUT <= 0;  //35 / 51 = 0
    16'b00100011_00110100 : OUT <= 0;  //35 / 52 = 0
    16'b00100011_00110101 : OUT <= 0;  //35 / 53 = 0
    16'b00100011_00110110 : OUT <= 0;  //35 / 54 = 0
    16'b00100011_00110111 : OUT <= 0;  //35 / 55 = 0
    16'b00100011_00111000 : OUT <= 0;  //35 / 56 = 0
    16'b00100011_00111001 : OUT <= 0;  //35 / 57 = 0
    16'b00100011_00111010 : OUT <= 0;  //35 / 58 = 0
    16'b00100011_00111011 : OUT <= 0;  //35 / 59 = 0
    16'b00100011_00111100 : OUT <= 0;  //35 / 60 = 0
    16'b00100011_00111101 : OUT <= 0;  //35 / 61 = 0
    16'b00100011_00111110 : OUT <= 0;  //35 / 62 = 0
    16'b00100011_00111111 : OUT <= 0;  //35 / 63 = 0
    16'b00100011_01000000 : OUT <= 0;  //35 / 64 = 0
    16'b00100011_01000001 : OUT <= 0;  //35 / 65 = 0
    16'b00100011_01000010 : OUT <= 0;  //35 / 66 = 0
    16'b00100011_01000011 : OUT <= 0;  //35 / 67 = 0
    16'b00100011_01000100 : OUT <= 0;  //35 / 68 = 0
    16'b00100011_01000101 : OUT <= 0;  //35 / 69 = 0
    16'b00100011_01000110 : OUT <= 0;  //35 / 70 = 0
    16'b00100011_01000111 : OUT <= 0;  //35 / 71 = 0
    16'b00100011_01001000 : OUT <= 0;  //35 / 72 = 0
    16'b00100011_01001001 : OUT <= 0;  //35 / 73 = 0
    16'b00100011_01001010 : OUT <= 0;  //35 / 74 = 0
    16'b00100011_01001011 : OUT <= 0;  //35 / 75 = 0
    16'b00100011_01001100 : OUT <= 0;  //35 / 76 = 0
    16'b00100011_01001101 : OUT <= 0;  //35 / 77 = 0
    16'b00100011_01001110 : OUT <= 0;  //35 / 78 = 0
    16'b00100011_01001111 : OUT <= 0;  //35 / 79 = 0
    16'b00100011_01010000 : OUT <= 0;  //35 / 80 = 0
    16'b00100011_01010001 : OUT <= 0;  //35 / 81 = 0
    16'b00100011_01010010 : OUT <= 0;  //35 / 82 = 0
    16'b00100011_01010011 : OUT <= 0;  //35 / 83 = 0
    16'b00100011_01010100 : OUT <= 0;  //35 / 84 = 0
    16'b00100011_01010101 : OUT <= 0;  //35 / 85 = 0
    16'b00100011_01010110 : OUT <= 0;  //35 / 86 = 0
    16'b00100011_01010111 : OUT <= 0;  //35 / 87 = 0
    16'b00100011_01011000 : OUT <= 0;  //35 / 88 = 0
    16'b00100011_01011001 : OUT <= 0;  //35 / 89 = 0
    16'b00100011_01011010 : OUT <= 0;  //35 / 90 = 0
    16'b00100011_01011011 : OUT <= 0;  //35 / 91 = 0
    16'b00100011_01011100 : OUT <= 0;  //35 / 92 = 0
    16'b00100011_01011101 : OUT <= 0;  //35 / 93 = 0
    16'b00100011_01011110 : OUT <= 0;  //35 / 94 = 0
    16'b00100011_01011111 : OUT <= 0;  //35 / 95 = 0
    16'b00100011_01100000 : OUT <= 0;  //35 / 96 = 0
    16'b00100011_01100001 : OUT <= 0;  //35 / 97 = 0
    16'b00100011_01100010 : OUT <= 0;  //35 / 98 = 0
    16'b00100011_01100011 : OUT <= 0;  //35 / 99 = 0
    16'b00100011_01100100 : OUT <= 0;  //35 / 100 = 0
    16'b00100011_01100101 : OUT <= 0;  //35 / 101 = 0
    16'b00100011_01100110 : OUT <= 0;  //35 / 102 = 0
    16'b00100011_01100111 : OUT <= 0;  //35 / 103 = 0
    16'b00100011_01101000 : OUT <= 0;  //35 / 104 = 0
    16'b00100011_01101001 : OUT <= 0;  //35 / 105 = 0
    16'b00100011_01101010 : OUT <= 0;  //35 / 106 = 0
    16'b00100011_01101011 : OUT <= 0;  //35 / 107 = 0
    16'b00100011_01101100 : OUT <= 0;  //35 / 108 = 0
    16'b00100011_01101101 : OUT <= 0;  //35 / 109 = 0
    16'b00100011_01101110 : OUT <= 0;  //35 / 110 = 0
    16'b00100011_01101111 : OUT <= 0;  //35 / 111 = 0
    16'b00100011_01110000 : OUT <= 0;  //35 / 112 = 0
    16'b00100011_01110001 : OUT <= 0;  //35 / 113 = 0
    16'b00100011_01110010 : OUT <= 0;  //35 / 114 = 0
    16'b00100011_01110011 : OUT <= 0;  //35 / 115 = 0
    16'b00100011_01110100 : OUT <= 0;  //35 / 116 = 0
    16'b00100011_01110101 : OUT <= 0;  //35 / 117 = 0
    16'b00100011_01110110 : OUT <= 0;  //35 / 118 = 0
    16'b00100011_01110111 : OUT <= 0;  //35 / 119 = 0
    16'b00100011_01111000 : OUT <= 0;  //35 / 120 = 0
    16'b00100011_01111001 : OUT <= 0;  //35 / 121 = 0
    16'b00100011_01111010 : OUT <= 0;  //35 / 122 = 0
    16'b00100011_01111011 : OUT <= 0;  //35 / 123 = 0
    16'b00100011_01111100 : OUT <= 0;  //35 / 124 = 0
    16'b00100011_01111101 : OUT <= 0;  //35 / 125 = 0
    16'b00100011_01111110 : OUT <= 0;  //35 / 126 = 0
    16'b00100011_01111111 : OUT <= 0;  //35 / 127 = 0
    16'b00100011_10000000 : OUT <= 0;  //35 / 128 = 0
    16'b00100011_10000001 : OUT <= 0;  //35 / 129 = 0
    16'b00100011_10000010 : OUT <= 0;  //35 / 130 = 0
    16'b00100011_10000011 : OUT <= 0;  //35 / 131 = 0
    16'b00100011_10000100 : OUT <= 0;  //35 / 132 = 0
    16'b00100011_10000101 : OUT <= 0;  //35 / 133 = 0
    16'b00100011_10000110 : OUT <= 0;  //35 / 134 = 0
    16'b00100011_10000111 : OUT <= 0;  //35 / 135 = 0
    16'b00100011_10001000 : OUT <= 0;  //35 / 136 = 0
    16'b00100011_10001001 : OUT <= 0;  //35 / 137 = 0
    16'b00100011_10001010 : OUT <= 0;  //35 / 138 = 0
    16'b00100011_10001011 : OUT <= 0;  //35 / 139 = 0
    16'b00100011_10001100 : OUT <= 0;  //35 / 140 = 0
    16'b00100011_10001101 : OUT <= 0;  //35 / 141 = 0
    16'b00100011_10001110 : OUT <= 0;  //35 / 142 = 0
    16'b00100011_10001111 : OUT <= 0;  //35 / 143 = 0
    16'b00100011_10010000 : OUT <= 0;  //35 / 144 = 0
    16'b00100011_10010001 : OUT <= 0;  //35 / 145 = 0
    16'b00100011_10010010 : OUT <= 0;  //35 / 146 = 0
    16'b00100011_10010011 : OUT <= 0;  //35 / 147 = 0
    16'b00100011_10010100 : OUT <= 0;  //35 / 148 = 0
    16'b00100011_10010101 : OUT <= 0;  //35 / 149 = 0
    16'b00100011_10010110 : OUT <= 0;  //35 / 150 = 0
    16'b00100011_10010111 : OUT <= 0;  //35 / 151 = 0
    16'b00100011_10011000 : OUT <= 0;  //35 / 152 = 0
    16'b00100011_10011001 : OUT <= 0;  //35 / 153 = 0
    16'b00100011_10011010 : OUT <= 0;  //35 / 154 = 0
    16'b00100011_10011011 : OUT <= 0;  //35 / 155 = 0
    16'b00100011_10011100 : OUT <= 0;  //35 / 156 = 0
    16'b00100011_10011101 : OUT <= 0;  //35 / 157 = 0
    16'b00100011_10011110 : OUT <= 0;  //35 / 158 = 0
    16'b00100011_10011111 : OUT <= 0;  //35 / 159 = 0
    16'b00100011_10100000 : OUT <= 0;  //35 / 160 = 0
    16'b00100011_10100001 : OUT <= 0;  //35 / 161 = 0
    16'b00100011_10100010 : OUT <= 0;  //35 / 162 = 0
    16'b00100011_10100011 : OUT <= 0;  //35 / 163 = 0
    16'b00100011_10100100 : OUT <= 0;  //35 / 164 = 0
    16'b00100011_10100101 : OUT <= 0;  //35 / 165 = 0
    16'b00100011_10100110 : OUT <= 0;  //35 / 166 = 0
    16'b00100011_10100111 : OUT <= 0;  //35 / 167 = 0
    16'b00100011_10101000 : OUT <= 0;  //35 / 168 = 0
    16'b00100011_10101001 : OUT <= 0;  //35 / 169 = 0
    16'b00100011_10101010 : OUT <= 0;  //35 / 170 = 0
    16'b00100011_10101011 : OUT <= 0;  //35 / 171 = 0
    16'b00100011_10101100 : OUT <= 0;  //35 / 172 = 0
    16'b00100011_10101101 : OUT <= 0;  //35 / 173 = 0
    16'b00100011_10101110 : OUT <= 0;  //35 / 174 = 0
    16'b00100011_10101111 : OUT <= 0;  //35 / 175 = 0
    16'b00100011_10110000 : OUT <= 0;  //35 / 176 = 0
    16'b00100011_10110001 : OUT <= 0;  //35 / 177 = 0
    16'b00100011_10110010 : OUT <= 0;  //35 / 178 = 0
    16'b00100011_10110011 : OUT <= 0;  //35 / 179 = 0
    16'b00100011_10110100 : OUT <= 0;  //35 / 180 = 0
    16'b00100011_10110101 : OUT <= 0;  //35 / 181 = 0
    16'b00100011_10110110 : OUT <= 0;  //35 / 182 = 0
    16'b00100011_10110111 : OUT <= 0;  //35 / 183 = 0
    16'b00100011_10111000 : OUT <= 0;  //35 / 184 = 0
    16'b00100011_10111001 : OUT <= 0;  //35 / 185 = 0
    16'b00100011_10111010 : OUT <= 0;  //35 / 186 = 0
    16'b00100011_10111011 : OUT <= 0;  //35 / 187 = 0
    16'b00100011_10111100 : OUT <= 0;  //35 / 188 = 0
    16'b00100011_10111101 : OUT <= 0;  //35 / 189 = 0
    16'b00100011_10111110 : OUT <= 0;  //35 / 190 = 0
    16'b00100011_10111111 : OUT <= 0;  //35 / 191 = 0
    16'b00100011_11000000 : OUT <= 0;  //35 / 192 = 0
    16'b00100011_11000001 : OUT <= 0;  //35 / 193 = 0
    16'b00100011_11000010 : OUT <= 0;  //35 / 194 = 0
    16'b00100011_11000011 : OUT <= 0;  //35 / 195 = 0
    16'b00100011_11000100 : OUT <= 0;  //35 / 196 = 0
    16'b00100011_11000101 : OUT <= 0;  //35 / 197 = 0
    16'b00100011_11000110 : OUT <= 0;  //35 / 198 = 0
    16'b00100011_11000111 : OUT <= 0;  //35 / 199 = 0
    16'b00100011_11001000 : OUT <= 0;  //35 / 200 = 0
    16'b00100011_11001001 : OUT <= 0;  //35 / 201 = 0
    16'b00100011_11001010 : OUT <= 0;  //35 / 202 = 0
    16'b00100011_11001011 : OUT <= 0;  //35 / 203 = 0
    16'b00100011_11001100 : OUT <= 0;  //35 / 204 = 0
    16'b00100011_11001101 : OUT <= 0;  //35 / 205 = 0
    16'b00100011_11001110 : OUT <= 0;  //35 / 206 = 0
    16'b00100011_11001111 : OUT <= 0;  //35 / 207 = 0
    16'b00100011_11010000 : OUT <= 0;  //35 / 208 = 0
    16'b00100011_11010001 : OUT <= 0;  //35 / 209 = 0
    16'b00100011_11010010 : OUT <= 0;  //35 / 210 = 0
    16'b00100011_11010011 : OUT <= 0;  //35 / 211 = 0
    16'b00100011_11010100 : OUT <= 0;  //35 / 212 = 0
    16'b00100011_11010101 : OUT <= 0;  //35 / 213 = 0
    16'b00100011_11010110 : OUT <= 0;  //35 / 214 = 0
    16'b00100011_11010111 : OUT <= 0;  //35 / 215 = 0
    16'b00100011_11011000 : OUT <= 0;  //35 / 216 = 0
    16'b00100011_11011001 : OUT <= 0;  //35 / 217 = 0
    16'b00100011_11011010 : OUT <= 0;  //35 / 218 = 0
    16'b00100011_11011011 : OUT <= 0;  //35 / 219 = 0
    16'b00100011_11011100 : OUT <= 0;  //35 / 220 = 0
    16'b00100011_11011101 : OUT <= 0;  //35 / 221 = 0
    16'b00100011_11011110 : OUT <= 0;  //35 / 222 = 0
    16'b00100011_11011111 : OUT <= 0;  //35 / 223 = 0
    16'b00100011_11100000 : OUT <= 0;  //35 / 224 = 0
    16'b00100011_11100001 : OUT <= 0;  //35 / 225 = 0
    16'b00100011_11100010 : OUT <= 0;  //35 / 226 = 0
    16'b00100011_11100011 : OUT <= 0;  //35 / 227 = 0
    16'b00100011_11100100 : OUT <= 0;  //35 / 228 = 0
    16'b00100011_11100101 : OUT <= 0;  //35 / 229 = 0
    16'b00100011_11100110 : OUT <= 0;  //35 / 230 = 0
    16'b00100011_11100111 : OUT <= 0;  //35 / 231 = 0
    16'b00100011_11101000 : OUT <= 0;  //35 / 232 = 0
    16'b00100011_11101001 : OUT <= 0;  //35 / 233 = 0
    16'b00100011_11101010 : OUT <= 0;  //35 / 234 = 0
    16'b00100011_11101011 : OUT <= 0;  //35 / 235 = 0
    16'b00100011_11101100 : OUT <= 0;  //35 / 236 = 0
    16'b00100011_11101101 : OUT <= 0;  //35 / 237 = 0
    16'b00100011_11101110 : OUT <= 0;  //35 / 238 = 0
    16'b00100011_11101111 : OUT <= 0;  //35 / 239 = 0
    16'b00100011_11110000 : OUT <= 0;  //35 / 240 = 0
    16'b00100011_11110001 : OUT <= 0;  //35 / 241 = 0
    16'b00100011_11110010 : OUT <= 0;  //35 / 242 = 0
    16'b00100011_11110011 : OUT <= 0;  //35 / 243 = 0
    16'b00100011_11110100 : OUT <= 0;  //35 / 244 = 0
    16'b00100011_11110101 : OUT <= 0;  //35 / 245 = 0
    16'b00100011_11110110 : OUT <= 0;  //35 / 246 = 0
    16'b00100011_11110111 : OUT <= 0;  //35 / 247 = 0
    16'b00100011_11111000 : OUT <= 0;  //35 / 248 = 0
    16'b00100011_11111001 : OUT <= 0;  //35 / 249 = 0
    16'b00100011_11111010 : OUT <= 0;  //35 / 250 = 0
    16'b00100011_11111011 : OUT <= 0;  //35 / 251 = 0
    16'b00100011_11111100 : OUT <= 0;  //35 / 252 = 0
    16'b00100011_11111101 : OUT <= 0;  //35 / 253 = 0
    16'b00100011_11111110 : OUT <= 0;  //35 / 254 = 0
    16'b00100011_11111111 : OUT <= 0;  //35 / 255 = 0
    16'b00100100_00000000 : OUT <= 0;  //36 / 0 = 0
    16'b00100100_00000001 : OUT <= 36;  //36 / 1 = 36
    16'b00100100_00000010 : OUT <= 18;  //36 / 2 = 18
    16'b00100100_00000011 : OUT <= 12;  //36 / 3 = 12
    16'b00100100_00000100 : OUT <= 9;  //36 / 4 = 9
    16'b00100100_00000101 : OUT <= 7;  //36 / 5 = 7
    16'b00100100_00000110 : OUT <= 6;  //36 / 6 = 6
    16'b00100100_00000111 : OUT <= 5;  //36 / 7 = 5
    16'b00100100_00001000 : OUT <= 4;  //36 / 8 = 4
    16'b00100100_00001001 : OUT <= 4;  //36 / 9 = 4
    16'b00100100_00001010 : OUT <= 3;  //36 / 10 = 3
    16'b00100100_00001011 : OUT <= 3;  //36 / 11 = 3
    16'b00100100_00001100 : OUT <= 3;  //36 / 12 = 3
    16'b00100100_00001101 : OUT <= 2;  //36 / 13 = 2
    16'b00100100_00001110 : OUT <= 2;  //36 / 14 = 2
    16'b00100100_00001111 : OUT <= 2;  //36 / 15 = 2
    16'b00100100_00010000 : OUT <= 2;  //36 / 16 = 2
    16'b00100100_00010001 : OUT <= 2;  //36 / 17 = 2
    16'b00100100_00010010 : OUT <= 2;  //36 / 18 = 2
    16'b00100100_00010011 : OUT <= 1;  //36 / 19 = 1
    16'b00100100_00010100 : OUT <= 1;  //36 / 20 = 1
    16'b00100100_00010101 : OUT <= 1;  //36 / 21 = 1
    16'b00100100_00010110 : OUT <= 1;  //36 / 22 = 1
    16'b00100100_00010111 : OUT <= 1;  //36 / 23 = 1
    16'b00100100_00011000 : OUT <= 1;  //36 / 24 = 1
    16'b00100100_00011001 : OUT <= 1;  //36 / 25 = 1
    16'b00100100_00011010 : OUT <= 1;  //36 / 26 = 1
    16'b00100100_00011011 : OUT <= 1;  //36 / 27 = 1
    16'b00100100_00011100 : OUT <= 1;  //36 / 28 = 1
    16'b00100100_00011101 : OUT <= 1;  //36 / 29 = 1
    16'b00100100_00011110 : OUT <= 1;  //36 / 30 = 1
    16'b00100100_00011111 : OUT <= 1;  //36 / 31 = 1
    16'b00100100_00100000 : OUT <= 1;  //36 / 32 = 1
    16'b00100100_00100001 : OUT <= 1;  //36 / 33 = 1
    16'b00100100_00100010 : OUT <= 1;  //36 / 34 = 1
    16'b00100100_00100011 : OUT <= 1;  //36 / 35 = 1
    16'b00100100_00100100 : OUT <= 1;  //36 / 36 = 1
    16'b00100100_00100101 : OUT <= 0;  //36 / 37 = 0
    16'b00100100_00100110 : OUT <= 0;  //36 / 38 = 0
    16'b00100100_00100111 : OUT <= 0;  //36 / 39 = 0
    16'b00100100_00101000 : OUT <= 0;  //36 / 40 = 0
    16'b00100100_00101001 : OUT <= 0;  //36 / 41 = 0
    16'b00100100_00101010 : OUT <= 0;  //36 / 42 = 0
    16'b00100100_00101011 : OUT <= 0;  //36 / 43 = 0
    16'b00100100_00101100 : OUT <= 0;  //36 / 44 = 0
    16'b00100100_00101101 : OUT <= 0;  //36 / 45 = 0
    16'b00100100_00101110 : OUT <= 0;  //36 / 46 = 0
    16'b00100100_00101111 : OUT <= 0;  //36 / 47 = 0
    16'b00100100_00110000 : OUT <= 0;  //36 / 48 = 0
    16'b00100100_00110001 : OUT <= 0;  //36 / 49 = 0
    16'b00100100_00110010 : OUT <= 0;  //36 / 50 = 0
    16'b00100100_00110011 : OUT <= 0;  //36 / 51 = 0
    16'b00100100_00110100 : OUT <= 0;  //36 / 52 = 0
    16'b00100100_00110101 : OUT <= 0;  //36 / 53 = 0
    16'b00100100_00110110 : OUT <= 0;  //36 / 54 = 0
    16'b00100100_00110111 : OUT <= 0;  //36 / 55 = 0
    16'b00100100_00111000 : OUT <= 0;  //36 / 56 = 0
    16'b00100100_00111001 : OUT <= 0;  //36 / 57 = 0
    16'b00100100_00111010 : OUT <= 0;  //36 / 58 = 0
    16'b00100100_00111011 : OUT <= 0;  //36 / 59 = 0
    16'b00100100_00111100 : OUT <= 0;  //36 / 60 = 0
    16'b00100100_00111101 : OUT <= 0;  //36 / 61 = 0
    16'b00100100_00111110 : OUT <= 0;  //36 / 62 = 0
    16'b00100100_00111111 : OUT <= 0;  //36 / 63 = 0
    16'b00100100_01000000 : OUT <= 0;  //36 / 64 = 0
    16'b00100100_01000001 : OUT <= 0;  //36 / 65 = 0
    16'b00100100_01000010 : OUT <= 0;  //36 / 66 = 0
    16'b00100100_01000011 : OUT <= 0;  //36 / 67 = 0
    16'b00100100_01000100 : OUT <= 0;  //36 / 68 = 0
    16'b00100100_01000101 : OUT <= 0;  //36 / 69 = 0
    16'b00100100_01000110 : OUT <= 0;  //36 / 70 = 0
    16'b00100100_01000111 : OUT <= 0;  //36 / 71 = 0
    16'b00100100_01001000 : OUT <= 0;  //36 / 72 = 0
    16'b00100100_01001001 : OUT <= 0;  //36 / 73 = 0
    16'b00100100_01001010 : OUT <= 0;  //36 / 74 = 0
    16'b00100100_01001011 : OUT <= 0;  //36 / 75 = 0
    16'b00100100_01001100 : OUT <= 0;  //36 / 76 = 0
    16'b00100100_01001101 : OUT <= 0;  //36 / 77 = 0
    16'b00100100_01001110 : OUT <= 0;  //36 / 78 = 0
    16'b00100100_01001111 : OUT <= 0;  //36 / 79 = 0
    16'b00100100_01010000 : OUT <= 0;  //36 / 80 = 0
    16'b00100100_01010001 : OUT <= 0;  //36 / 81 = 0
    16'b00100100_01010010 : OUT <= 0;  //36 / 82 = 0
    16'b00100100_01010011 : OUT <= 0;  //36 / 83 = 0
    16'b00100100_01010100 : OUT <= 0;  //36 / 84 = 0
    16'b00100100_01010101 : OUT <= 0;  //36 / 85 = 0
    16'b00100100_01010110 : OUT <= 0;  //36 / 86 = 0
    16'b00100100_01010111 : OUT <= 0;  //36 / 87 = 0
    16'b00100100_01011000 : OUT <= 0;  //36 / 88 = 0
    16'b00100100_01011001 : OUT <= 0;  //36 / 89 = 0
    16'b00100100_01011010 : OUT <= 0;  //36 / 90 = 0
    16'b00100100_01011011 : OUT <= 0;  //36 / 91 = 0
    16'b00100100_01011100 : OUT <= 0;  //36 / 92 = 0
    16'b00100100_01011101 : OUT <= 0;  //36 / 93 = 0
    16'b00100100_01011110 : OUT <= 0;  //36 / 94 = 0
    16'b00100100_01011111 : OUT <= 0;  //36 / 95 = 0
    16'b00100100_01100000 : OUT <= 0;  //36 / 96 = 0
    16'b00100100_01100001 : OUT <= 0;  //36 / 97 = 0
    16'b00100100_01100010 : OUT <= 0;  //36 / 98 = 0
    16'b00100100_01100011 : OUT <= 0;  //36 / 99 = 0
    16'b00100100_01100100 : OUT <= 0;  //36 / 100 = 0
    16'b00100100_01100101 : OUT <= 0;  //36 / 101 = 0
    16'b00100100_01100110 : OUT <= 0;  //36 / 102 = 0
    16'b00100100_01100111 : OUT <= 0;  //36 / 103 = 0
    16'b00100100_01101000 : OUT <= 0;  //36 / 104 = 0
    16'b00100100_01101001 : OUT <= 0;  //36 / 105 = 0
    16'b00100100_01101010 : OUT <= 0;  //36 / 106 = 0
    16'b00100100_01101011 : OUT <= 0;  //36 / 107 = 0
    16'b00100100_01101100 : OUT <= 0;  //36 / 108 = 0
    16'b00100100_01101101 : OUT <= 0;  //36 / 109 = 0
    16'b00100100_01101110 : OUT <= 0;  //36 / 110 = 0
    16'b00100100_01101111 : OUT <= 0;  //36 / 111 = 0
    16'b00100100_01110000 : OUT <= 0;  //36 / 112 = 0
    16'b00100100_01110001 : OUT <= 0;  //36 / 113 = 0
    16'b00100100_01110010 : OUT <= 0;  //36 / 114 = 0
    16'b00100100_01110011 : OUT <= 0;  //36 / 115 = 0
    16'b00100100_01110100 : OUT <= 0;  //36 / 116 = 0
    16'b00100100_01110101 : OUT <= 0;  //36 / 117 = 0
    16'b00100100_01110110 : OUT <= 0;  //36 / 118 = 0
    16'b00100100_01110111 : OUT <= 0;  //36 / 119 = 0
    16'b00100100_01111000 : OUT <= 0;  //36 / 120 = 0
    16'b00100100_01111001 : OUT <= 0;  //36 / 121 = 0
    16'b00100100_01111010 : OUT <= 0;  //36 / 122 = 0
    16'b00100100_01111011 : OUT <= 0;  //36 / 123 = 0
    16'b00100100_01111100 : OUT <= 0;  //36 / 124 = 0
    16'b00100100_01111101 : OUT <= 0;  //36 / 125 = 0
    16'b00100100_01111110 : OUT <= 0;  //36 / 126 = 0
    16'b00100100_01111111 : OUT <= 0;  //36 / 127 = 0
    16'b00100100_10000000 : OUT <= 0;  //36 / 128 = 0
    16'b00100100_10000001 : OUT <= 0;  //36 / 129 = 0
    16'b00100100_10000010 : OUT <= 0;  //36 / 130 = 0
    16'b00100100_10000011 : OUT <= 0;  //36 / 131 = 0
    16'b00100100_10000100 : OUT <= 0;  //36 / 132 = 0
    16'b00100100_10000101 : OUT <= 0;  //36 / 133 = 0
    16'b00100100_10000110 : OUT <= 0;  //36 / 134 = 0
    16'b00100100_10000111 : OUT <= 0;  //36 / 135 = 0
    16'b00100100_10001000 : OUT <= 0;  //36 / 136 = 0
    16'b00100100_10001001 : OUT <= 0;  //36 / 137 = 0
    16'b00100100_10001010 : OUT <= 0;  //36 / 138 = 0
    16'b00100100_10001011 : OUT <= 0;  //36 / 139 = 0
    16'b00100100_10001100 : OUT <= 0;  //36 / 140 = 0
    16'b00100100_10001101 : OUT <= 0;  //36 / 141 = 0
    16'b00100100_10001110 : OUT <= 0;  //36 / 142 = 0
    16'b00100100_10001111 : OUT <= 0;  //36 / 143 = 0
    16'b00100100_10010000 : OUT <= 0;  //36 / 144 = 0
    16'b00100100_10010001 : OUT <= 0;  //36 / 145 = 0
    16'b00100100_10010010 : OUT <= 0;  //36 / 146 = 0
    16'b00100100_10010011 : OUT <= 0;  //36 / 147 = 0
    16'b00100100_10010100 : OUT <= 0;  //36 / 148 = 0
    16'b00100100_10010101 : OUT <= 0;  //36 / 149 = 0
    16'b00100100_10010110 : OUT <= 0;  //36 / 150 = 0
    16'b00100100_10010111 : OUT <= 0;  //36 / 151 = 0
    16'b00100100_10011000 : OUT <= 0;  //36 / 152 = 0
    16'b00100100_10011001 : OUT <= 0;  //36 / 153 = 0
    16'b00100100_10011010 : OUT <= 0;  //36 / 154 = 0
    16'b00100100_10011011 : OUT <= 0;  //36 / 155 = 0
    16'b00100100_10011100 : OUT <= 0;  //36 / 156 = 0
    16'b00100100_10011101 : OUT <= 0;  //36 / 157 = 0
    16'b00100100_10011110 : OUT <= 0;  //36 / 158 = 0
    16'b00100100_10011111 : OUT <= 0;  //36 / 159 = 0
    16'b00100100_10100000 : OUT <= 0;  //36 / 160 = 0
    16'b00100100_10100001 : OUT <= 0;  //36 / 161 = 0
    16'b00100100_10100010 : OUT <= 0;  //36 / 162 = 0
    16'b00100100_10100011 : OUT <= 0;  //36 / 163 = 0
    16'b00100100_10100100 : OUT <= 0;  //36 / 164 = 0
    16'b00100100_10100101 : OUT <= 0;  //36 / 165 = 0
    16'b00100100_10100110 : OUT <= 0;  //36 / 166 = 0
    16'b00100100_10100111 : OUT <= 0;  //36 / 167 = 0
    16'b00100100_10101000 : OUT <= 0;  //36 / 168 = 0
    16'b00100100_10101001 : OUT <= 0;  //36 / 169 = 0
    16'b00100100_10101010 : OUT <= 0;  //36 / 170 = 0
    16'b00100100_10101011 : OUT <= 0;  //36 / 171 = 0
    16'b00100100_10101100 : OUT <= 0;  //36 / 172 = 0
    16'b00100100_10101101 : OUT <= 0;  //36 / 173 = 0
    16'b00100100_10101110 : OUT <= 0;  //36 / 174 = 0
    16'b00100100_10101111 : OUT <= 0;  //36 / 175 = 0
    16'b00100100_10110000 : OUT <= 0;  //36 / 176 = 0
    16'b00100100_10110001 : OUT <= 0;  //36 / 177 = 0
    16'b00100100_10110010 : OUT <= 0;  //36 / 178 = 0
    16'b00100100_10110011 : OUT <= 0;  //36 / 179 = 0
    16'b00100100_10110100 : OUT <= 0;  //36 / 180 = 0
    16'b00100100_10110101 : OUT <= 0;  //36 / 181 = 0
    16'b00100100_10110110 : OUT <= 0;  //36 / 182 = 0
    16'b00100100_10110111 : OUT <= 0;  //36 / 183 = 0
    16'b00100100_10111000 : OUT <= 0;  //36 / 184 = 0
    16'b00100100_10111001 : OUT <= 0;  //36 / 185 = 0
    16'b00100100_10111010 : OUT <= 0;  //36 / 186 = 0
    16'b00100100_10111011 : OUT <= 0;  //36 / 187 = 0
    16'b00100100_10111100 : OUT <= 0;  //36 / 188 = 0
    16'b00100100_10111101 : OUT <= 0;  //36 / 189 = 0
    16'b00100100_10111110 : OUT <= 0;  //36 / 190 = 0
    16'b00100100_10111111 : OUT <= 0;  //36 / 191 = 0
    16'b00100100_11000000 : OUT <= 0;  //36 / 192 = 0
    16'b00100100_11000001 : OUT <= 0;  //36 / 193 = 0
    16'b00100100_11000010 : OUT <= 0;  //36 / 194 = 0
    16'b00100100_11000011 : OUT <= 0;  //36 / 195 = 0
    16'b00100100_11000100 : OUT <= 0;  //36 / 196 = 0
    16'b00100100_11000101 : OUT <= 0;  //36 / 197 = 0
    16'b00100100_11000110 : OUT <= 0;  //36 / 198 = 0
    16'b00100100_11000111 : OUT <= 0;  //36 / 199 = 0
    16'b00100100_11001000 : OUT <= 0;  //36 / 200 = 0
    16'b00100100_11001001 : OUT <= 0;  //36 / 201 = 0
    16'b00100100_11001010 : OUT <= 0;  //36 / 202 = 0
    16'b00100100_11001011 : OUT <= 0;  //36 / 203 = 0
    16'b00100100_11001100 : OUT <= 0;  //36 / 204 = 0
    16'b00100100_11001101 : OUT <= 0;  //36 / 205 = 0
    16'b00100100_11001110 : OUT <= 0;  //36 / 206 = 0
    16'b00100100_11001111 : OUT <= 0;  //36 / 207 = 0
    16'b00100100_11010000 : OUT <= 0;  //36 / 208 = 0
    16'b00100100_11010001 : OUT <= 0;  //36 / 209 = 0
    16'b00100100_11010010 : OUT <= 0;  //36 / 210 = 0
    16'b00100100_11010011 : OUT <= 0;  //36 / 211 = 0
    16'b00100100_11010100 : OUT <= 0;  //36 / 212 = 0
    16'b00100100_11010101 : OUT <= 0;  //36 / 213 = 0
    16'b00100100_11010110 : OUT <= 0;  //36 / 214 = 0
    16'b00100100_11010111 : OUT <= 0;  //36 / 215 = 0
    16'b00100100_11011000 : OUT <= 0;  //36 / 216 = 0
    16'b00100100_11011001 : OUT <= 0;  //36 / 217 = 0
    16'b00100100_11011010 : OUT <= 0;  //36 / 218 = 0
    16'b00100100_11011011 : OUT <= 0;  //36 / 219 = 0
    16'b00100100_11011100 : OUT <= 0;  //36 / 220 = 0
    16'b00100100_11011101 : OUT <= 0;  //36 / 221 = 0
    16'b00100100_11011110 : OUT <= 0;  //36 / 222 = 0
    16'b00100100_11011111 : OUT <= 0;  //36 / 223 = 0
    16'b00100100_11100000 : OUT <= 0;  //36 / 224 = 0
    16'b00100100_11100001 : OUT <= 0;  //36 / 225 = 0
    16'b00100100_11100010 : OUT <= 0;  //36 / 226 = 0
    16'b00100100_11100011 : OUT <= 0;  //36 / 227 = 0
    16'b00100100_11100100 : OUT <= 0;  //36 / 228 = 0
    16'b00100100_11100101 : OUT <= 0;  //36 / 229 = 0
    16'b00100100_11100110 : OUT <= 0;  //36 / 230 = 0
    16'b00100100_11100111 : OUT <= 0;  //36 / 231 = 0
    16'b00100100_11101000 : OUT <= 0;  //36 / 232 = 0
    16'b00100100_11101001 : OUT <= 0;  //36 / 233 = 0
    16'b00100100_11101010 : OUT <= 0;  //36 / 234 = 0
    16'b00100100_11101011 : OUT <= 0;  //36 / 235 = 0
    16'b00100100_11101100 : OUT <= 0;  //36 / 236 = 0
    16'b00100100_11101101 : OUT <= 0;  //36 / 237 = 0
    16'b00100100_11101110 : OUT <= 0;  //36 / 238 = 0
    16'b00100100_11101111 : OUT <= 0;  //36 / 239 = 0
    16'b00100100_11110000 : OUT <= 0;  //36 / 240 = 0
    16'b00100100_11110001 : OUT <= 0;  //36 / 241 = 0
    16'b00100100_11110010 : OUT <= 0;  //36 / 242 = 0
    16'b00100100_11110011 : OUT <= 0;  //36 / 243 = 0
    16'b00100100_11110100 : OUT <= 0;  //36 / 244 = 0
    16'b00100100_11110101 : OUT <= 0;  //36 / 245 = 0
    16'b00100100_11110110 : OUT <= 0;  //36 / 246 = 0
    16'b00100100_11110111 : OUT <= 0;  //36 / 247 = 0
    16'b00100100_11111000 : OUT <= 0;  //36 / 248 = 0
    16'b00100100_11111001 : OUT <= 0;  //36 / 249 = 0
    16'b00100100_11111010 : OUT <= 0;  //36 / 250 = 0
    16'b00100100_11111011 : OUT <= 0;  //36 / 251 = 0
    16'b00100100_11111100 : OUT <= 0;  //36 / 252 = 0
    16'b00100100_11111101 : OUT <= 0;  //36 / 253 = 0
    16'b00100100_11111110 : OUT <= 0;  //36 / 254 = 0
    16'b00100100_11111111 : OUT <= 0;  //36 / 255 = 0
    16'b00100101_00000000 : OUT <= 0;  //37 / 0 = 0
    16'b00100101_00000001 : OUT <= 37;  //37 / 1 = 37
    16'b00100101_00000010 : OUT <= 18;  //37 / 2 = 18
    16'b00100101_00000011 : OUT <= 12;  //37 / 3 = 12
    16'b00100101_00000100 : OUT <= 9;  //37 / 4 = 9
    16'b00100101_00000101 : OUT <= 7;  //37 / 5 = 7
    16'b00100101_00000110 : OUT <= 6;  //37 / 6 = 6
    16'b00100101_00000111 : OUT <= 5;  //37 / 7 = 5
    16'b00100101_00001000 : OUT <= 4;  //37 / 8 = 4
    16'b00100101_00001001 : OUT <= 4;  //37 / 9 = 4
    16'b00100101_00001010 : OUT <= 3;  //37 / 10 = 3
    16'b00100101_00001011 : OUT <= 3;  //37 / 11 = 3
    16'b00100101_00001100 : OUT <= 3;  //37 / 12 = 3
    16'b00100101_00001101 : OUT <= 2;  //37 / 13 = 2
    16'b00100101_00001110 : OUT <= 2;  //37 / 14 = 2
    16'b00100101_00001111 : OUT <= 2;  //37 / 15 = 2
    16'b00100101_00010000 : OUT <= 2;  //37 / 16 = 2
    16'b00100101_00010001 : OUT <= 2;  //37 / 17 = 2
    16'b00100101_00010010 : OUT <= 2;  //37 / 18 = 2
    16'b00100101_00010011 : OUT <= 1;  //37 / 19 = 1
    16'b00100101_00010100 : OUT <= 1;  //37 / 20 = 1
    16'b00100101_00010101 : OUT <= 1;  //37 / 21 = 1
    16'b00100101_00010110 : OUT <= 1;  //37 / 22 = 1
    16'b00100101_00010111 : OUT <= 1;  //37 / 23 = 1
    16'b00100101_00011000 : OUT <= 1;  //37 / 24 = 1
    16'b00100101_00011001 : OUT <= 1;  //37 / 25 = 1
    16'b00100101_00011010 : OUT <= 1;  //37 / 26 = 1
    16'b00100101_00011011 : OUT <= 1;  //37 / 27 = 1
    16'b00100101_00011100 : OUT <= 1;  //37 / 28 = 1
    16'b00100101_00011101 : OUT <= 1;  //37 / 29 = 1
    16'b00100101_00011110 : OUT <= 1;  //37 / 30 = 1
    16'b00100101_00011111 : OUT <= 1;  //37 / 31 = 1
    16'b00100101_00100000 : OUT <= 1;  //37 / 32 = 1
    16'b00100101_00100001 : OUT <= 1;  //37 / 33 = 1
    16'b00100101_00100010 : OUT <= 1;  //37 / 34 = 1
    16'b00100101_00100011 : OUT <= 1;  //37 / 35 = 1
    16'b00100101_00100100 : OUT <= 1;  //37 / 36 = 1
    16'b00100101_00100101 : OUT <= 1;  //37 / 37 = 1
    16'b00100101_00100110 : OUT <= 0;  //37 / 38 = 0
    16'b00100101_00100111 : OUT <= 0;  //37 / 39 = 0
    16'b00100101_00101000 : OUT <= 0;  //37 / 40 = 0
    16'b00100101_00101001 : OUT <= 0;  //37 / 41 = 0
    16'b00100101_00101010 : OUT <= 0;  //37 / 42 = 0
    16'b00100101_00101011 : OUT <= 0;  //37 / 43 = 0
    16'b00100101_00101100 : OUT <= 0;  //37 / 44 = 0
    16'b00100101_00101101 : OUT <= 0;  //37 / 45 = 0
    16'b00100101_00101110 : OUT <= 0;  //37 / 46 = 0
    16'b00100101_00101111 : OUT <= 0;  //37 / 47 = 0
    16'b00100101_00110000 : OUT <= 0;  //37 / 48 = 0
    16'b00100101_00110001 : OUT <= 0;  //37 / 49 = 0
    16'b00100101_00110010 : OUT <= 0;  //37 / 50 = 0
    16'b00100101_00110011 : OUT <= 0;  //37 / 51 = 0
    16'b00100101_00110100 : OUT <= 0;  //37 / 52 = 0
    16'b00100101_00110101 : OUT <= 0;  //37 / 53 = 0
    16'b00100101_00110110 : OUT <= 0;  //37 / 54 = 0
    16'b00100101_00110111 : OUT <= 0;  //37 / 55 = 0
    16'b00100101_00111000 : OUT <= 0;  //37 / 56 = 0
    16'b00100101_00111001 : OUT <= 0;  //37 / 57 = 0
    16'b00100101_00111010 : OUT <= 0;  //37 / 58 = 0
    16'b00100101_00111011 : OUT <= 0;  //37 / 59 = 0
    16'b00100101_00111100 : OUT <= 0;  //37 / 60 = 0
    16'b00100101_00111101 : OUT <= 0;  //37 / 61 = 0
    16'b00100101_00111110 : OUT <= 0;  //37 / 62 = 0
    16'b00100101_00111111 : OUT <= 0;  //37 / 63 = 0
    16'b00100101_01000000 : OUT <= 0;  //37 / 64 = 0
    16'b00100101_01000001 : OUT <= 0;  //37 / 65 = 0
    16'b00100101_01000010 : OUT <= 0;  //37 / 66 = 0
    16'b00100101_01000011 : OUT <= 0;  //37 / 67 = 0
    16'b00100101_01000100 : OUT <= 0;  //37 / 68 = 0
    16'b00100101_01000101 : OUT <= 0;  //37 / 69 = 0
    16'b00100101_01000110 : OUT <= 0;  //37 / 70 = 0
    16'b00100101_01000111 : OUT <= 0;  //37 / 71 = 0
    16'b00100101_01001000 : OUT <= 0;  //37 / 72 = 0
    16'b00100101_01001001 : OUT <= 0;  //37 / 73 = 0
    16'b00100101_01001010 : OUT <= 0;  //37 / 74 = 0
    16'b00100101_01001011 : OUT <= 0;  //37 / 75 = 0
    16'b00100101_01001100 : OUT <= 0;  //37 / 76 = 0
    16'b00100101_01001101 : OUT <= 0;  //37 / 77 = 0
    16'b00100101_01001110 : OUT <= 0;  //37 / 78 = 0
    16'b00100101_01001111 : OUT <= 0;  //37 / 79 = 0
    16'b00100101_01010000 : OUT <= 0;  //37 / 80 = 0
    16'b00100101_01010001 : OUT <= 0;  //37 / 81 = 0
    16'b00100101_01010010 : OUT <= 0;  //37 / 82 = 0
    16'b00100101_01010011 : OUT <= 0;  //37 / 83 = 0
    16'b00100101_01010100 : OUT <= 0;  //37 / 84 = 0
    16'b00100101_01010101 : OUT <= 0;  //37 / 85 = 0
    16'b00100101_01010110 : OUT <= 0;  //37 / 86 = 0
    16'b00100101_01010111 : OUT <= 0;  //37 / 87 = 0
    16'b00100101_01011000 : OUT <= 0;  //37 / 88 = 0
    16'b00100101_01011001 : OUT <= 0;  //37 / 89 = 0
    16'b00100101_01011010 : OUT <= 0;  //37 / 90 = 0
    16'b00100101_01011011 : OUT <= 0;  //37 / 91 = 0
    16'b00100101_01011100 : OUT <= 0;  //37 / 92 = 0
    16'b00100101_01011101 : OUT <= 0;  //37 / 93 = 0
    16'b00100101_01011110 : OUT <= 0;  //37 / 94 = 0
    16'b00100101_01011111 : OUT <= 0;  //37 / 95 = 0
    16'b00100101_01100000 : OUT <= 0;  //37 / 96 = 0
    16'b00100101_01100001 : OUT <= 0;  //37 / 97 = 0
    16'b00100101_01100010 : OUT <= 0;  //37 / 98 = 0
    16'b00100101_01100011 : OUT <= 0;  //37 / 99 = 0
    16'b00100101_01100100 : OUT <= 0;  //37 / 100 = 0
    16'b00100101_01100101 : OUT <= 0;  //37 / 101 = 0
    16'b00100101_01100110 : OUT <= 0;  //37 / 102 = 0
    16'b00100101_01100111 : OUT <= 0;  //37 / 103 = 0
    16'b00100101_01101000 : OUT <= 0;  //37 / 104 = 0
    16'b00100101_01101001 : OUT <= 0;  //37 / 105 = 0
    16'b00100101_01101010 : OUT <= 0;  //37 / 106 = 0
    16'b00100101_01101011 : OUT <= 0;  //37 / 107 = 0
    16'b00100101_01101100 : OUT <= 0;  //37 / 108 = 0
    16'b00100101_01101101 : OUT <= 0;  //37 / 109 = 0
    16'b00100101_01101110 : OUT <= 0;  //37 / 110 = 0
    16'b00100101_01101111 : OUT <= 0;  //37 / 111 = 0
    16'b00100101_01110000 : OUT <= 0;  //37 / 112 = 0
    16'b00100101_01110001 : OUT <= 0;  //37 / 113 = 0
    16'b00100101_01110010 : OUT <= 0;  //37 / 114 = 0
    16'b00100101_01110011 : OUT <= 0;  //37 / 115 = 0
    16'b00100101_01110100 : OUT <= 0;  //37 / 116 = 0
    16'b00100101_01110101 : OUT <= 0;  //37 / 117 = 0
    16'b00100101_01110110 : OUT <= 0;  //37 / 118 = 0
    16'b00100101_01110111 : OUT <= 0;  //37 / 119 = 0
    16'b00100101_01111000 : OUT <= 0;  //37 / 120 = 0
    16'b00100101_01111001 : OUT <= 0;  //37 / 121 = 0
    16'b00100101_01111010 : OUT <= 0;  //37 / 122 = 0
    16'b00100101_01111011 : OUT <= 0;  //37 / 123 = 0
    16'b00100101_01111100 : OUT <= 0;  //37 / 124 = 0
    16'b00100101_01111101 : OUT <= 0;  //37 / 125 = 0
    16'b00100101_01111110 : OUT <= 0;  //37 / 126 = 0
    16'b00100101_01111111 : OUT <= 0;  //37 / 127 = 0
    16'b00100101_10000000 : OUT <= 0;  //37 / 128 = 0
    16'b00100101_10000001 : OUT <= 0;  //37 / 129 = 0
    16'b00100101_10000010 : OUT <= 0;  //37 / 130 = 0
    16'b00100101_10000011 : OUT <= 0;  //37 / 131 = 0
    16'b00100101_10000100 : OUT <= 0;  //37 / 132 = 0
    16'b00100101_10000101 : OUT <= 0;  //37 / 133 = 0
    16'b00100101_10000110 : OUT <= 0;  //37 / 134 = 0
    16'b00100101_10000111 : OUT <= 0;  //37 / 135 = 0
    16'b00100101_10001000 : OUT <= 0;  //37 / 136 = 0
    16'b00100101_10001001 : OUT <= 0;  //37 / 137 = 0
    16'b00100101_10001010 : OUT <= 0;  //37 / 138 = 0
    16'b00100101_10001011 : OUT <= 0;  //37 / 139 = 0
    16'b00100101_10001100 : OUT <= 0;  //37 / 140 = 0
    16'b00100101_10001101 : OUT <= 0;  //37 / 141 = 0
    16'b00100101_10001110 : OUT <= 0;  //37 / 142 = 0
    16'b00100101_10001111 : OUT <= 0;  //37 / 143 = 0
    16'b00100101_10010000 : OUT <= 0;  //37 / 144 = 0
    16'b00100101_10010001 : OUT <= 0;  //37 / 145 = 0
    16'b00100101_10010010 : OUT <= 0;  //37 / 146 = 0
    16'b00100101_10010011 : OUT <= 0;  //37 / 147 = 0
    16'b00100101_10010100 : OUT <= 0;  //37 / 148 = 0
    16'b00100101_10010101 : OUT <= 0;  //37 / 149 = 0
    16'b00100101_10010110 : OUT <= 0;  //37 / 150 = 0
    16'b00100101_10010111 : OUT <= 0;  //37 / 151 = 0
    16'b00100101_10011000 : OUT <= 0;  //37 / 152 = 0
    16'b00100101_10011001 : OUT <= 0;  //37 / 153 = 0
    16'b00100101_10011010 : OUT <= 0;  //37 / 154 = 0
    16'b00100101_10011011 : OUT <= 0;  //37 / 155 = 0
    16'b00100101_10011100 : OUT <= 0;  //37 / 156 = 0
    16'b00100101_10011101 : OUT <= 0;  //37 / 157 = 0
    16'b00100101_10011110 : OUT <= 0;  //37 / 158 = 0
    16'b00100101_10011111 : OUT <= 0;  //37 / 159 = 0
    16'b00100101_10100000 : OUT <= 0;  //37 / 160 = 0
    16'b00100101_10100001 : OUT <= 0;  //37 / 161 = 0
    16'b00100101_10100010 : OUT <= 0;  //37 / 162 = 0
    16'b00100101_10100011 : OUT <= 0;  //37 / 163 = 0
    16'b00100101_10100100 : OUT <= 0;  //37 / 164 = 0
    16'b00100101_10100101 : OUT <= 0;  //37 / 165 = 0
    16'b00100101_10100110 : OUT <= 0;  //37 / 166 = 0
    16'b00100101_10100111 : OUT <= 0;  //37 / 167 = 0
    16'b00100101_10101000 : OUT <= 0;  //37 / 168 = 0
    16'b00100101_10101001 : OUT <= 0;  //37 / 169 = 0
    16'b00100101_10101010 : OUT <= 0;  //37 / 170 = 0
    16'b00100101_10101011 : OUT <= 0;  //37 / 171 = 0
    16'b00100101_10101100 : OUT <= 0;  //37 / 172 = 0
    16'b00100101_10101101 : OUT <= 0;  //37 / 173 = 0
    16'b00100101_10101110 : OUT <= 0;  //37 / 174 = 0
    16'b00100101_10101111 : OUT <= 0;  //37 / 175 = 0
    16'b00100101_10110000 : OUT <= 0;  //37 / 176 = 0
    16'b00100101_10110001 : OUT <= 0;  //37 / 177 = 0
    16'b00100101_10110010 : OUT <= 0;  //37 / 178 = 0
    16'b00100101_10110011 : OUT <= 0;  //37 / 179 = 0
    16'b00100101_10110100 : OUT <= 0;  //37 / 180 = 0
    16'b00100101_10110101 : OUT <= 0;  //37 / 181 = 0
    16'b00100101_10110110 : OUT <= 0;  //37 / 182 = 0
    16'b00100101_10110111 : OUT <= 0;  //37 / 183 = 0
    16'b00100101_10111000 : OUT <= 0;  //37 / 184 = 0
    16'b00100101_10111001 : OUT <= 0;  //37 / 185 = 0
    16'b00100101_10111010 : OUT <= 0;  //37 / 186 = 0
    16'b00100101_10111011 : OUT <= 0;  //37 / 187 = 0
    16'b00100101_10111100 : OUT <= 0;  //37 / 188 = 0
    16'b00100101_10111101 : OUT <= 0;  //37 / 189 = 0
    16'b00100101_10111110 : OUT <= 0;  //37 / 190 = 0
    16'b00100101_10111111 : OUT <= 0;  //37 / 191 = 0
    16'b00100101_11000000 : OUT <= 0;  //37 / 192 = 0
    16'b00100101_11000001 : OUT <= 0;  //37 / 193 = 0
    16'b00100101_11000010 : OUT <= 0;  //37 / 194 = 0
    16'b00100101_11000011 : OUT <= 0;  //37 / 195 = 0
    16'b00100101_11000100 : OUT <= 0;  //37 / 196 = 0
    16'b00100101_11000101 : OUT <= 0;  //37 / 197 = 0
    16'b00100101_11000110 : OUT <= 0;  //37 / 198 = 0
    16'b00100101_11000111 : OUT <= 0;  //37 / 199 = 0
    16'b00100101_11001000 : OUT <= 0;  //37 / 200 = 0
    16'b00100101_11001001 : OUT <= 0;  //37 / 201 = 0
    16'b00100101_11001010 : OUT <= 0;  //37 / 202 = 0
    16'b00100101_11001011 : OUT <= 0;  //37 / 203 = 0
    16'b00100101_11001100 : OUT <= 0;  //37 / 204 = 0
    16'b00100101_11001101 : OUT <= 0;  //37 / 205 = 0
    16'b00100101_11001110 : OUT <= 0;  //37 / 206 = 0
    16'b00100101_11001111 : OUT <= 0;  //37 / 207 = 0
    16'b00100101_11010000 : OUT <= 0;  //37 / 208 = 0
    16'b00100101_11010001 : OUT <= 0;  //37 / 209 = 0
    16'b00100101_11010010 : OUT <= 0;  //37 / 210 = 0
    16'b00100101_11010011 : OUT <= 0;  //37 / 211 = 0
    16'b00100101_11010100 : OUT <= 0;  //37 / 212 = 0
    16'b00100101_11010101 : OUT <= 0;  //37 / 213 = 0
    16'b00100101_11010110 : OUT <= 0;  //37 / 214 = 0
    16'b00100101_11010111 : OUT <= 0;  //37 / 215 = 0
    16'b00100101_11011000 : OUT <= 0;  //37 / 216 = 0
    16'b00100101_11011001 : OUT <= 0;  //37 / 217 = 0
    16'b00100101_11011010 : OUT <= 0;  //37 / 218 = 0
    16'b00100101_11011011 : OUT <= 0;  //37 / 219 = 0
    16'b00100101_11011100 : OUT <= 0;  //37 / 220 = 0
    16'b00100101_11011101 : OUT <= 0;  //37 / 221 = 0
    16'b00100101_11011110 : OUT <= 0;  //37 / 222 = 0
    16'b00100101_11011111 : OUT <= 0;  //37 / 223 = 0
    16'b00100101_11100000 : OUT <= 0;  //37 / 224 = 0
    16'b00100101_11100001 : OUT <= 0;  //37 / 225 = 0
    16'b00100101_11100010 : OUT <= 0;  //37 / 226 = 0
    16'b00100101_11100011 : OUT <= 0;  //37 / 227 = 0
    16'b00100101_11100100 : OUT <= 0;  //37 / 228 = 0
    16'b00100101_11100101 : OUT <= 0;  //37 / 229 = 0
    16'b00100101_11100110 : OUT <= 0;  //37 / 230 = 0
    16'b00100101_11100111 : OUT <= 0;  //37 / 231 = 0
    16'b00100101_11101000 : OUT <= 0;  //37 / 232 = 0
    16'b00100101_11101001 : OUT <= 0;  //37 / 233 = 0
    16'b00100101_11101010 : OUT <= 0;  //37 / 234 = 0
    16'b00100101_11101011 : OUT <= 0;  //37 / 235 = 0
    16'b00100101_11101100 : OUT <= 0;  //37 / 236 = 0
    16'b00100101_11101101 : OUT <= 0;  //37 / 237 = 0
    16'b00100101_11101110 : OUT <= 0;  //37 / 238 = 0
    16'b00100101_11101111 : OUT <= 0;  //37 / 239 = 0
    16'b00100101_11110000 : OUT <= 0;  //37 / 240 = 0
    16'b00100101_11110001 : OUT <= 0;  //37 / 241 = 0
    16'b00100101_11110010 : OUT <= 0;  //37 / 242 = 0
    16'b00100101_11110011 : OUT <= 0;  //37 / 243 = 0
    16'b00100101_11110100 : OUT <= 0;  //37 / 244 = 0
    16'b00100101_11110101 : OUT <= 0;  //37 / 245 = 0
    16'b00100101_11110110 : OUT <= 0;  //37 / 246 = 0
    16'b00100101_11110111 : OUT <= 0;  //37 / 247 = 0
    16'b00100101_11111000 : OUT <= 0;  //37 / 248 = 0
    16'b00100101_11111001 : OUT <= 0;  //37 / 249 = 0
    16'b00100101_11111010 : OUT <= 0;  //37 / 250 = 0
    16'b00100101_11111011 : OUT <= 0;  //37 / 251 = 0
    16'b00100101_11111100 : OUT <= 0;  //37 / 252 = 0
    16'b00100101_11111101 : OUT <= 0;  //37 / 253 = 0
    16'b00100101_11111110 : OUT <= 0;  //37 / 254 = 0
    16'b00100101_11111111 : OUT <= 0;  //37 / 255 = 0
    16'b00100110_00000000 : OUT <= 0;  //38 / 0 = 0
    16'b00100110_00000001 : OUT <= 38;  //38 / 1 = 38
    16'b00100110_00000010 : OUT <= 19;  //38 / 2 = 19
    16'b00100110_00000011 : OUT <= 12;  //38 / 3 = 12
    16'b00100110_00000100 : OUT <= 9;  //38 / 4 = 9
    16'b00100110_00000101 : OUT <= 7;  //38 / 5 = 7
    16'b00100110_00000110 : OUT <= 6;  //38 / 6 = 6
    16'b00100110_00000111 : OUT <= 5;  //38 / 7 = 5
    16'b00100110_00001000 : OUT <= 4;  //38 / 8 = 4
    16'b00100110_00001001 : OUT <= 4;  //38 / 9 = 4
    16'b00100110_00001010 : OUT <= 3;  //38 / 10 = 3
    16'b00100110_00001011 : OUT <= 3;  //38 / 11 = 3
    16'b00100110_00001100 : OUT <= 3;  //38 / 12 = 3
    16'b00100110_00001101 : OUT <= 2;  //38 / 13 = 2
    16'b00100110_00001110 : OUT <= 2;  //38 / 14 = 2
    16'b00100110_00001111 : OUT <= 2;  //38 / 15 = 2
    16'b00100110_00010000 : OUT <= 2;  //38 / 16 = 2
    16'b00100110_00010001 : OUT <= 2;  //38 / 17 = 2
    16'b00100110_00010010 : OUT <= 2;  //38 / 18 = 2
    16'b00100110_00010011 : OUT <= 2;  //38 / 19 = 2
    16'b00100110_00010100 : OUT <= 1;  //38 / 20 = 1
    16'b00100110_00010101 : OUT <= 1;  //38 / 21 = 1
    16'b00100110_00010110 : OUT <= 1;  //38 / 22 = 1
    16'b00100110_00010111 : OUT <= 1;  //38 / 23 = 1
    16'b00100110_00011000 : OUT <= 1;  //38 / 24 = 1
    16'b00100110_00011001 : OUT <= 1;  //38 / 25 = 1
    16'b00100110_00011010 : OUT <= 1;  //38 / 26 = 1
    16'b00100110_00011011 : OUT <= 1;  //38 / 27 = 1
    16'b00100110_00011100 : OUT <= 1;  //38 / 28 = 1
    16'b00100110_00011101 : OUT <= 1;  //38 / 29 = 1
    16'b00100110_00011110 : OUT <= 1;  //38 / 30 = 1
    16'b00100110_00011111 : OUT <= 1;  //38 / 31 = 1
    16'b00100110_00100000 : OUT <= 1;  //38 / 32 = 1
    16'b00100110_00100001 : OUT <= 1;  //38 / 33 = 1
    16'b00100110_00100010 : OUT <= 1;  //38 / 34 = 1
    16'b00100110_00100011 : OUT <= 1;  //38 / 35 = 1
    16'b00100110_00100100 : OUT <= 1;  //38 / 36 = 1
    16'b00100110_00100101 : OUT <= 1;  //38 / 37 = 1
    16'b00100110_00100110 : OUT <= 1;  //38 / 38 = 1
    16'b00100110_00100111 : OUT <= 0;  //38 / 39 = 0
    16'b00100110_00101000 : OUT <= 0;  //38 / 40 = 0
    16'b00100110_00101001 : OUT <= 0;  //38 / 41 = 0
    16'b00100110_00101010 : OUT <= 0;  //38 / 42 = 0
    16'b00100110_00101011 : OUT <= 0;  //38 / 43 = 0
    16'b00100110_00101100 : OUT <= 0;  //38 / 44 = 0
    16'b00100110_00101101 : OUT <= 0;  //38 / 45 = 0
    16'b00100110_00101110 : OUT <= 0;  //38 / 46 = 0
    16'b00100110_00101111 : OUT <= 0;  //38 / 47 = 0
    16'b00100110_00110000 : OUT <= 0;  //38 / 48 = 0
    16'b00100110_00110001 : OUT <= 0;  //38 / 49 = 0
    16'b00100110_00110010 : OUT <= 0;  //38 / 50 = 0
    16'b00100110_00110011 : OUT <= 0;  //38 / 51 = 0
    16'b00100110_00110100 : OUT <= 0;  //38 / 52 = 0
    16'b00100110_00110101 : OUT <= 0;  //38 / 53 = 0
    16'b00100110_00110110 : OUT <= 0;  //38 / 54 = 0
    16'b00100110_00110111 : OUT <= 0;  //38 / 55 = 0
    16'b00100110_00111000 : OUT <= 0;  //38 / 56 = 0
    16'b00100110_00111001 : OUT <= 0;  //38 / 57 = 0
    16'b00100110_00111010 : OUT <= 0;  //38 / 58 = 0
    16'b00100110_00111011 : OUT <= 0;  //38 / 59 = 0
    16'b00100110_00111100 : OUT <= 0;  //38 / 60 = 0
    16'b00100110_00111101 : OUT <= 0;  //38 / 61 = 0
    16'b00100110_00111110 : OUT <= 0;  //38 / 62 = 0
    16'b00100110_00111111 : OUT <= 0;  //38 / 63 = 0
    16'b00100110_01000000 : OUT <= 0;  //38 / 64 = 0
    16'b00100110_01000001 : OUT <= 0;  //38 / 65 = 0
    16'b00100110_01000010 : OUT <= 0;  //38 / 66 = 0
    16'b00100110_01000011 : OUT <= 0;  //38 / 67 = 0
    16'b00100110_01000100 : OUT <= 0;  //38 / 68 = 0
    16'b00100110_01000101 : OUT <= 0;  //38 / 69 = 0
    16'b00100110_01000110 : OUT <= 0;  //38 / 70 = 0
    16'b00100110_01000111 : OUT <= 0;  //38 / 71 = 0
    16'b00100110_01001000 : OUT <= 0;  //38 / 72 = 0
    16'b00100110_01001001 : OUT <= 0;  //38 / 73 = 0
    16'b00100110_01001010 : OUT <= 0;  //38 / 74 = 0
    16'b00100110_01001011 : OUT <= 0;  //38 / 75 = 0
    16'b00100110_01001100 : OUT <= 0;  //38 / 76 = 0
    16'b00100110_01001101 : OUT <= 0;  //38 / 77 = 0
    16'b00100110_01001110 : OUT <= 0;  //38 / 78 = 0
    16'b00100110_01001111 : OUT <= 0;  //38 / 79 = 0
    16'b00100110_01010000 : OUT <= 0;  //38 / 80 = 0
    16'b00100110_01010001 : OUT <= 0;  //38 / 81 = 0
    16'b00100110_01010010 : OUT <= 0;  //38 / 82 = 0
    16'b00100110_01010011 : OUT <= 0;  //38 / 83 = 0
    16'b00100110_01010100 : OUT <= 0;  //38 / 84 = 0
    16'b00100110_01010101 : OUT <= 0;  //38 / 85 = 0
    16'b00100110_01010110 : OUT <= 0;  //38 / 86 = 0
    16'b00100110_01010111 : OUT <= 0;  //38 / 87 = 0
    16'b00100110_01011000 : OUT <= 0;  //38 / 88 = 0
    16'b00100110_01011001 : OUT <= 0;  //38 / 89 = 0
    16'b00100110_01011010 : OUT <= 0;  //38 / 90 = 0
    16'b00100110_01011011 : OUT <= 0;  //38 / 91 = 0
    16'b00100110_01011100 : OUT <= 0;  //38 / 92 = 0
    16'b00100110_01011101 : OUT <= 0;  //38 / 93 = 0
    16'b00100110_01011110 : OUT <= 0;  //38 / 94 = 0
    16'b00100110_01011111 : OUT <= 0;  //38 / 95 = 0
    16'b00100110_01100000 : OUT <= 0;  //38 / 96 = 0
    16'b00100110_01100001 : OUT <= 0;  //38 / 97 = 0
    16'b00100110_01100010 : OUT <= 0;  //38 / 98 = 0
    16'b00100110_01100011 : OUT <= 0;  //38 / 99 = 0
    16'b00100110_01100100 : OUT <= 0;  //38 / 100 = 0
    16'b00100110_01100101 : OUT <= 0;  //38 / 101 = 0
    16'b00100110_01100110 : OUT <= 0;  //38 / 102 = 0
    16'b00100110_01100111 : OUT <= 0;  //38 / 103 = 0
    16'b00100110_01101000 : OUT <= 0;  //38 / 104 = 0
    16'b00100110_01101001 : OUT <= 0;  //38 / 105 = 0
    16'b00100110_01101010 : OUT <= 0;  //38 / 106 = 0
    16'b00100110_01101011 : OUT <= 0;  //38 / 107 = 0
    16'b00100110_01101100 : OUT <= 0;  //38 / 108 = 0
    16'b00100110_01101101 : OUT <= 0;  //38 / 109 = 0
    16'b00100110_01101110 : OUT <= 0;  //38 / 110 = 0
    16'b00100110_01101111 : OUT <= 0;  //38 / 111 = 0
    16'b00100110_01110000 : OUT <= 0;  //38 / 112 = 0
    16'b00100110_01110001 : OUT <= 0;  //38 / 113 = 0
    16'b00100110_01110010 : OUT <= 0;  //38 / 114 = 0
    16'b00100110_01110011 : OUT <= 0;  //38 / 115 = 0
    16'b00100110_01110100 : OUT <= 0;  //38 / 116 = 0
    16'b00100110_01110101 : OUT <= 0;  //38 / 117 = 0
    16'b00100110_01110110 : OUT <= 0;  //38 / 118 = 0
    16'b00100110_01110111 : OUT <= 0;  //38 / 119 = 0
    16'b00100110_01111000 : OUT <= 0;  //38 / 120 = 0
    16'b00100110_01111001 : OUT <= 0;  //38 / 121 = 0
    16'b00100110_01111010 : OUT <= 0;  //38 / 122 = 0
    16'b00100110_01111011 : OUT <= 0;  //38 / 123 = 0
    16'b00100110_01111100 : OUT <= 0;  //38 / 124 = 0
    16'b00100110_01111101 : OUT <= 0;  //38 / 125 = 0
    16'b00100110_01111110 : OUT <= 0;  //38 / 126 = 0
    16'b00100110_01111111 : OUT <= 0;  //38 / 127 = 0
    16'b00100110_10000000 : OUT <= 0;  //38 / 128 = 0
    16'b00100110_10000001 : OUT <= 0;  //38 / 129 = 0
    16'b00100110_10000010 : OUT <= 0;  //38 / 130 = 0
    16'b00100110_10000011 : OUT <= 0;  //38 / 131 = 0
    16'b00100110_10000100 : OUT <= 0;  //38 / 132 = 0
    16'b00100110_10000101 : OUT <= 0;  //38 / 133 = 0
    16'b00100110_10000110 : OUT <= 0;  //38 / 134 = 0
    16'b00100110_10000111 : OUT <= 0;  //38 / 135 = 0
    16'b00100110_10001000 : OUT <= 0;  //38 / 136 = 0
    16'b00100110_10001001 : OUT <= 0;  //38 / 137 = 0
    16'b00100110_10001010 : OUT <= 0;  //38 / 138 = 0
    16'b00100110_10001011 : OUT <= 0;  //38 / 139 = 0
    16'b00100110_10001100 : OUT <= 0;  //38 / 140 = 0
    16'b00100110_10001101 : OUT <= 0;  //38 / 141 = 0
    16'b00100110_10001110 : OUT <= 0;  //38 / 142 = 0
    16'b00100110_10001111 : OUT <= 0;  //38 / 143 = 0
    16'b00100110_10010000 : OUT <= 0;  //38 / 144 = 0
    16'b00100110_10010001 : OUT <= 0;  //38 / 145 = 0
    16'b00100110_10010010 : OUT <= 0;  //38 / 146 = 0
    16'b00100110_10010011 : OUT <= 0;  //38 / 147 = 0
    16'b00100110_10010100 : OUT <= 0;  //38 / 148 = 0
    16'b00100110_10010101 : OUT <= 0;  //38 / 149 = 0
    16'b00100110_10010110 : OUT <= 0;  //38 / 150 = 0
    16'b00100110_10010111 : OUT <= 0;  //38 / 151 = 0
    16'b00100110_10011000 : OUT <= 0;  //38 / 152 = 0
    16'b00100110_10011001 : OUT <= 0;  //38 / 153 = 0
    16'b00100110_10011010 : OUT <= 0;  //38 / 154 = 0
    16'b00100110_10011011 : OUT <= 0;  //38 / 155 = 0
    16'b00100110_10011100 : OUT <= 0;  //38 / 156 = 0
    16'b00100110_10011101 : OUT <= 0;  //38 / 157 = 0
    16'b00100110_10011110 : OUT <= 0;  //38 / 158 = 0
    16'b00100110_10011111 : OUT <= 0;  //38 / 159 = 0
    16'b00100110_10100000 : OUT <= 0;  //38 / 160 = 0
    16'b00100110_10100001 : OUT <= 0;  //38 / 161 = 0
    16'b00100110_10100010 : OUT <= 0;  //38 / 162 = 0
    16'b00100110_10100011 : OUT <= 0;  //38 / 163 = 0
    16'b00100110_10100100 : OUT <= 0;  //38 / 164 = 0
    16'b00100110_10100101 : OUT <= 0;  //38 / 165 = 0
    16'b00100110_10100110 : OUT <= 0;  //38 / 166 = 0
    16'b00100110_10100111 : OUT <= 0;  //38 / 167 = 0
    16'b00100110_10101000 : OUT <= 0;  //38 / 168 = 0
    16'b00100110_10101001 : OUT <= 0;  //38 / 169 = 0
    16'b00100110_10101010 : OUT <= 0;  //38 / 170 = 0
    16'b00100110_10101011 : OUT <= 0;  //38 / 171 = 0
    16'b00100110_10101100 : OUT <= 0;  //38 / 172 = 0
    16'b00100110_10101101 : OUT <= 0;  //38 / 173 = 0
    16'b00100110_10101110 : OUT <= 0;  //38 / 174 = 0
    16'b00100110_10101111 : OUT <= 0;  //38 / 175 = 0
    16'b00100110_10110000 : OUT <= 0;  //38 / 176 = 0
    16'b00100110_10110001 : OUT <= 0;  //38 / 177 = 0
    16'b00100110_10110010 : OUT <= 0;  //38 / 178 = 0
    16'b00100110_10110011 : OUT <= 0;  //38 / 179 = 0
    16'b00100110_10110100 : OUT <= 0;  //38 / 180 = 0
    16'b00100110_10110101 : OUT <= 0;  //38 / 181 = 0
    16'b00100110_10110110 : OUT <= 0;  //38 / 182 = 0
    16'b00100110_10110111 : OUT <= 0;  //38 / 183 = 0
    16'b00100110_10111000 : OUT <= 0;  //38 / 184 = 0
    16'b00100110_10111001 : OUT <= 0;  //38 / 185 = 0
    16'b00100110_10111010 : OUT <= 0;  //38 / 186 = 0
    16'b00100110_10111011 : OUT <= 0;  //38 / 187 = 0
    16'b00100110_10111100 : OUT <= 0;  //38 / 188 = 0
    16'b00100110_10111101 : OUT <= 0;  //38 / 189 = 0
    16'b00100110_10111110 : OUT <= 0;  //38 / 190 = 0
    16'b00100110_10111111 : OUT <= 0;  //38 / 191 = 0
    16'b00100110_11000000 : OUT <= 0;  //38 / 192 = 0
    16'b00100110_11000001 : OUT <= 0;  //38 / 193 = 0
    16'b00100110_11000010 : OUT <= 0;  //38 / 194 = 0
    16'b00100110_11000011 : OUT <= 0;  //38 / 195 = 0
    16'b00100110_11000100 : OUT <= 0;  //38 / 196 = 0
    16'b00100110_11000101 : OUT <= 0;  //38 / 197 = 0
    16'b00100110_11000110 : OUT <= 0;  //38 / 198 = 0
    16'b00100110_11000111 : OUT <= 0;  //38 / 199 = 0
    16'b00100110_11001000 : OUT <= 0;  //38 / 200 = 0
    16'b00100110_11001001 : OUT <= 0;  //38 / 201 = 0
    16'b00100110_11001010 : OUT <= 0;  //38 / 202 = 0
    16'b00100110_11001011 : OUT <= 0;  //38 / 203 = 0
    16'b00100110_11001100 : OUT <= 0;  //38 / 204 = 0
    16'b00100110_11001101 : OUT <= 0;  //38 / 205 = 0
    16'b00100110_11001110 : OUT <= 0;  //38 / 206 = 0
    16'b00100110_11001111 : OUT <= 0;  //38 / 207 = 0
    16'b00100110_11010000 : OUT <= 0;  //38 / 208 = 0
    16'b00100110_11010001 : OUT <= 0;  //38 / 209 = 0
    16'b00100110_11010010 : OUT <= 0;  //38 / 210 = 0
    16'b00100110_11010011 : OUT <= 0;  //38 / 211 = 0
    16'b00100110_11010100 : OUT <= 0;  //38 / 212 = 0
    16'b00100110_11010101 : OUT <= 0;  //38 / 213 = 0
    16'b00100110_11010110 : OUT <= 0;  //38 / 214 = 0
    16'b00100110_11010111 : OUT <= 0;  //38 / 215 = 0
    16'b00100110_11011000 : OUT <= 0;  //38 / 216 = 0
    16'b00100110_11011001 : OUT <= 0;  //38 / 217 = 0
    16'b00100110_11011010 : OUT <= 0;  //38 / 218 = 0
    16'b00100110_11011011 : OUT <= 0;  //38 / 219 = 0
    16'b00100110_11011100 : OUT <= 0;  //38 / 220 = 0
    16'b00100110_11011101 : OUT <= 0;  //38 / 221 = 0
    16'b00100110_11011110 : OUT <= 0;  //38 / 222 = 0
    16'b00100110_11011111 : OUT <= 0;  //38 / 223 = 0
    16'b00100110_11100000 : OUT <= 0;  //38 / 224 = 0
    16'b00100110_11100001 : OUT <= 0;  //38 / 225 = 0
    16'b00100110_11100010 : OUT <= 0;  //38 / 226 = 0
    16'b00100110_11100011 : OUT <= 0;  //38 / 227 = 0
    16'b00100110_11100100 : OUT <= 0;  //38 / 228 = 0
    16'b00100110_11100101 : OUT <= 0;  //38 / 229 = 0
    16'b00100110_11100110 : OUT <= 0;  //38 / 230 = 0
    16'b00100110_11100111 : OUT <= 0;  //38 / 231 = 0
    16'b00100110_11101000 : OUT <= 0;  //38 / 232 = 0
    16'b00100110_11101001 : OUT <= 0;  //38 / 233 = 0
    16'b00100110_11101010 : OUT <= 0;  //38 / 234 = 0
    16'b00100110_11101011 : OUT <= 0;  //38 / 235 = 0
    16'b00100110_11101100 : OUT <= 0;  //38 / 236 = 0
    16'b00100110_11101101 : OUT <= 0;  //38 / 237 = 0
    16'b00100110_11101110 : OUT <= 0;  //38 / 238 = 0
    16'b00100110_11101111 : OUT <= 0;  //38 / 239 = 0
    16'b00100110_11110000 : OUT <= 0;  //38 / 240 = 0
    16'b00100110_11110001 : OUT <= 0;  //38 / 241 = 0
    16'b00100110_11110010 : OUT <= 0;  //38 / 242 = 0
    16'b00100110_11110011 : OUT <= 0;  //38 / 243 = 0
    16'b00100110_11110100 : OUT <= 0;  //38 / 244 = 0
    16'b00100110_11110101 : OUT <= 0;  //38 / 245 = 0
    16'b00100110_11110110 : OUT <= 0;  //38 / 246 = 0
    16'b00100110_11110111 : OUT <= 0;  //38 / 247 = 0
    16'b00100110_11111000 : OUT <= 0;  //38 / 248 = 0
    16'b00100110_11111001 : OUT <= 0;  //38 / 249 = 0
    16'b00100110_11111010 : OUT <= 0;  //38 / 250 = 0
    16'b00100110_11111011 : OUT <= 0;  //38 / 251 = 0
    16'b00100110_11111100 : OUT <= 0;  //38 / 252 = 0
    16'b00100110_11111101 : OUT <= 0;  //38 / 253 = 0
    16'b00100110_11111110 : OUT <= 0;  //38 / 254 = 0
    16'b00100110_11111111 : OUT <= 0;  //38 / 255 = 0
    16'b00100111_00000000 : OUT <= 0;  //39 / 0 = 0
    16'b00100111_00000001 : OUT <= 39;  //39 / 1 = 39
    16'b00100111_00000010 : OUT <= 19;  //39 / 2 = 19
    16'b00100111_00000011 : OUT <= 13;  //39 / 3 = 13
    16'b00100111_00000100 : OUT <= 9;  //39 / 4 = 9
    16'b00100111_00000101 : OUT <= 7;  //39 / 5 = 7
    16'b00100111_00000110 : OUT <= 6;  //39 / 6 = 6
    16'b00100111_00000111 : OUT <= 5;  //39 / 7 = 5
    16'b00100111_00001000 : OUT <= 4;  //39 / 8 = 4
    16'b00100111_00001001 : OUT <= 4;  //39 / 9 = 4
    16'b00100111_00001010 : OUT <= 3;  //39 / 10 = 3
    16'b00100111_00001011 : OUT <= 3;  //39 / 11 = 3
    16'b00100111_00001100 : OUT <= 3;  //39 / 12 = 3
    16'b00100111_00001101 : OUT <= 3;  //39 / 13 = 3
    16'b00100111_00001110 : OUT <= 2;  //39 / 14 = 2
    16'b00100111_00001111 : OUT <= 2;  //39 / 15 = 2
    16'b00100111_00010000 : OUT <= 2;  //39 / 16 = 2
    16'b00100111_00010001 : OUT <= 2;  //39 / 17 = 2
    16'b00100111_00010010 : OUT <= 2;  //39 / 18 = 2
    16'b00100111_00010011 : OUT <= 2;  //39 / 19 = 2
    16'b00100111_00010100 : OUT <= 1;  //39 / 20 = 1
    16'b00100111_00010101 : OUT <= 1;  //39 / 21 = 1
    16'b00100111_00010110 : OUT <= 1;  //39 / 22 = 1
    16'b00100111_00010111 : OUT <= 1;  //39 / 23 = 1
    16'b00100111_00011000 : OUT <= 1;  //39 / 24 = 1
    16'b00100111_00011001 : OUT <= 1;  //39 / 25 = 1
    16'b00100111_00011010 : OUT <= 1;  //39 / 26 = 1
    16'b00100111_00011011 : OUT <= 1;  //39 / 27 = 1
    16'b00100111_00011100 : OUT <= 1;  //39 / 28 = 1
    16'b00100111_00011101 : OUT <= 1;  //39 / 29 = 1
    16'b00100111_00011110 : OUT <= 1;  //39 / 30 = 1
    16'b00100111_00011111 : OUT <= 1;  //39 / 31 = 1
    16'b00100111_00100000 : OUT <= 1;  //39 / 32 = 1
    16'b00100111_00100001 : OUT <= 1;  //39 / 33 = 1
    16'b00100111_00100010 : OUT <= 1;  //39 / 34 = 1
    16'b00100111_00100011 : OUT <= 1;  //39 / 35 = 1
    16'b00100111_00100100 : OUT <= 1;  //39 / 36 = 1
    16'b00100111_00100101 : OUT <= 1;  //39 / 37 = 1
    16'b00100111_00100110 : OUT <= 1;  //39 / 38 = 1
    16'b00100111_00100111 : OUT <= 1;  //39 / 39 = 1
    16'b00100111_00101000 : OUT <= 0;  //39 / 40 = 0
    16'b00100111_00101001 : OUT <= 0;  //39 / 41 = 0
    16'b00100111_00101010 : OUT <= 0;  //39 / 42 = 0
    16'b00100111_00101011 : OUT <= 0;  //39 / 43 = 0
    16'b00100111_00101100 : OUT <= 0;  //39 / 44 = 0
    16'b00100111_00101101 : OUT <= 0;  //39 / 45 = 0
    16'b00100111_00101110 : OUT <= 0;  //39 / 46 = 0
    16'b00100111_00101111 : OUT <= 0;  //39 / 47 = 0
    16'b00100111_00110000 : OUT <= 0;  //39 / 48 = 0
    16'b00100111_00110001 : OUT <= 0;  //39 / 49 = 0
    16'b00100111_00110010 : OUT <= 0;  //39 / 50 = 0
    16'b00100111_00110011 : OUT <= 0;  //39 / 51 = 0
    16'b00100111_00110100 : OUT <= 0;  //39 / 52 = 0
    16'b00100111_00110101 : OUT <= 0;  //39 / 53 = 0
    16'b00100111_00110110 : OUT <= 0;  //39 / 54 = 0
    16'b00100111_00110111 : OUT <= 0;  //39 / 55 = 0
    16'b00100111_00111000 : OUT <= 0;  //39 / 56 = 0
    16'b00100111_00111001 : OUT <= 0;  //39 / 57 = 0
    16'b00100111_00111010 : OUT <= 0;  //39 / 58 = 0
    16'b00100111_00111011 : OUT <= 0;  //39 / 59 = 0
    16'b00100111_00111100 : OUT <= 0;  //39 / 60 = 0
    16'b00100111_00111101 : OUT <= 0;  //39 / 61 = 0
    16'b00100111_00111110 : OUT <= 0;  //39 / 62 = 0
    16'b00100111_00111111 : OUT <= 0;  //39 / 63 = 0
    16'b00100111_01000000 : OUT <= 0;  //39 / 64 = 0
    16'b00100111_01000001 : OUT <= 0;  //39 / 65 = 0
    16'b00100111_01000010 : OUT <= 0;  //39 / 66 = 0
    16'b00100111_01000011 : OUT <= 0;  //39 / 67 = 0
    16'b00100111_01000100 : OUT <= 0;  //39 / 68 = 0
    16'b00100111_01000101 : OUT <= 0;  //39 / 69 = 0
    16'b00100111_01000110 : OUT <= 0;  //39 / 70 = 0
    16'b00100111_01000111 : OUT <= 0;  //39 / 71 = 0
    16'b00100111_01001000 : OUT <= 0;  //39 / 72 = 0
    16'b00100111_01001001 : OUT <= 0;  //39 / 73 = 0
    16'b00100111_01001010 : OUT <= 0;  //39 / 74 = 0
    16'b00100111_01001011 : OUT <= 0;  //39 / 75 = 0
    16'b00100111_01001100 : OUT <= 0;  //39 / 76 = 0
    16'b00100111_01001101 : OUT <= 0;  //39 / 77 = 0
    16'b00100111_01001110 : OUT <= 0;  //39 / 78 = 0
    16'b00100111_01001111 : OUT <= 0;  //39 / 79 = 0
    16'b00100111_01010000 : OUT <= 0;  //39 / 80 = 0
    16'b00100111_01010001 : OUT <= 0;  //39 / 81 = 0
    16'b00100111_01010010 : OUT <= 0;  //39 / 82 = 0
    16'b00100111_01010011 : OUT <= 0;  //39 / 83 = 0
    16'b00100111_01010100 : OUT <= 0;  //39 / 84 = 0
    16'b00100111_01010101 : OUT <= 0;  //39 / 85 = 0
    16'b00100111_01010110 : OUT <= 0;  //39 / 86 = 0
    16'b00100111_01010111 : OUT <= 0;  //39 / 87 = 0
    16'b00100111_01011000 : OUT <= 0;  //39 / 88 = 0
    16'b00100111_01011001 : OUT <= 0;  //39 / 89 = 0
    16'b00100111_01011010 : OUT <= 0;  //39 / 90 = 0
    16'b00100111_01011011 : OUT <= 0;  //39 / 91 = 0
    16'b00100111_01011100 : OUT <= 0;  //39 / 92 = 0
    16'b00100111_01011101 : OUT <= 0;  //39 / 93 = 0
    16'b00100111_01011110 : OUT <= 0;  //39 / 94 = 0
    16'b00100111_01011111 : OUT <= 0;  //39 / 95 = 0
    16'b00100111_01100000 : OUT <= 0;  //39 / 96 = 0
    16'b00100111_01100001 : OUT <= 0;  //39 / 97 = 0
    16'b00100111_01100010 : OUT <= 0;  //39 / 98 = 0
    16'b00100111_01100011 : OUT <= 0;  //39 / 99 = 0
    16'b00100111_01100100 : OUT <= 0;  //39 / 100 = 0
    16'b00100111_01100101 : OUT <= 0;  //39 / 101 = 0
    16'b00100111_01100110 : OUT <= 0;  //39 / 102 = 0
    16'b00100111_01100111 : OUT <= 0;  //39 / 103 = 0
    16'b00100111_01101000 : OUT <= 0;  //39 / 104 = 0
    16'b00100111_01101001 : OUT <= 0;  //39 / 105 = 0
    16'b00100111_01101010 : OUT <= 0;  //39 / 106 = 0
    16'b00100111_01101011 : OUT <= 0;  //39 / 107 = 0
    16'b00100111_01101100 : OUT <= 0;  //39 / 108 = 0
    16'b00100111_01101101 : OUT <= 0;  //39 / 109 = 0
    16'b00100111_01101110 : OUT <= 0;  //39 / 110 = 0
    16'b00100111_01101111 : OUT <= 0;  //39 / 111 = 0
    16'b00100111_01110000 : OUT <= 0;  //39 / 112 = 0
    16'b00100111_01110001 : OUT <= 0;  //39 / 113 = 0
    16'b00100111_01110010 : OUT <= 0;  //39 / 114 = 0
    16'b00100111_01110011 : OUT <= 0;  //39 / 115 = 0
    16'b00100111_01110100 : OUT <= 0;  //39 / 116 = 0
    16'b00100111_01110101 : OUT <= 0;  //39 / 117 = 0
    16'b00100111_01110110 : OUT <= 0;  //39 / 118 = 0
    16'b00100111_01110111 : OUT <= 0;  //39 / 119 = 0
    16'b00100111_01111000 : OUT <= 0;  //39 / 120 = 0
    16'b00100111_01111001 : OUT <= 0;  //39 / 121 = 0
    16'b00100111_01111010 : OUT <= 0;  //39 / 122 = 0
    16'b00100111_01111011 : OUT <= 0;  //39 / 123 = 0
    16'b00100111_01111100 : OUT <= 0;  //39 / 124 = 0
    16'b00100111_01111101 : OUT <= 0;  //39 / 125 = 0
    16'b00100111_01111110 : OUT <= 0;  //39 / 126 = 0
    16'b00100111_01111111 : OUT <= 0;  //39 / 127 = 0
    16'b00100111_10000000 : OUT <= 0;  //39 / 128 = 0
    16'b00100111_10000001 : OUT <= 0;  //39 / 129 = 0
    16'b00100111_10000010 : OUT <= 0;  //39 / 130 = 0
    16'b00100111_10000011 : OUT <= 0;  //39 / 131 = 0
    16'b00100111_10000100 : OUT <= 0;  //39 / 132 = 0
    16'b00100111_10000101 : OUT <= 0;  //39 / 133 = 0
    16'b00100111_10000110 : OUT <= 0;  //39 / 134 = 0
    16'b00100111_10000111 : OUT <= 0;  //39 / 135 = 0
    16'b00100111_10001000 : OUT <= 0;  //39 / 136 = 0
    16'b00100111_10001001 : OUT <= 0;  //39 / 137 = 0
    16'b00100111_10001010 : OUT <= 0;  //39 / 138 = 0
    16'b00100111_10001011 : OUT <= 0;  //39 / 139 = 0
    16'b00100111_10001100 : OUT <= 0;  //39 / 140 = 0
    16'b00100111_10001101 : OUT <= 0;  //39 / 141 = 0
    16'b00100111_10001110 : OUT <= 0;  //39 / 142 = 0
    16'b00100111_10001111 : OUT <= 0;  //39 / 143 = 0
    16'b00100111_10010000 : OUT <= 0;  //39 / 144 = 0
    16'b00100111_10010001 : OUT <= 0;  //39 / 145 = 0
    16'b00100111_10010010 : OUT <= 0;  //39 / 146 = 0
    16'b00100111_10010011 : OUT <= 0;  //39 / 147 = 0
    16'b00100111_10010100 : OUT <= 0;  //39 / 148 = 0
    16'b00100111_10010101 : OUT <= 0;  //39 / 149 = 0
    16'b00100111_10010110 : OUT <= 0;  //39 / 150 = 0
    16'b00100111_10010111 : OUT <= 0;  //39 / 151 = 0
    16'b00100111_10011000 : OUT <= 0;  //39 / 152 = 0
    16'b00100111_10011001 : OUT <= 0;  //39 / 153 = 0
    16'b00100111_10011010 : OUT <= 0;  //39 / 154 = 0
    16'b00100111_10011011 : OUT <= 0;  //39 / 155 = 0
    16'b00100111_10011100 : OUT <= 0;  //39 / 156 = 0
    16'b00100111_10011101 : OUT <= 0;  //39 / 157 = 0
    16'b00100111_10011110 : OUT <= 0;  //39 / 158 = 0
    16'b00100111_10011111 : OUT <= 0;  //39 / 159 = 0
    16'b00100111_10100000 : OUT <= 0;  //39 / 160 = 0
    16'b00100111_10100001 : OUT <= 0;  //39 / 161 = 0
    16'b00100111_10100010 : OUT <= 0;  //39 / 162 = 0
    16'b00100111_10100011 : OUT <= 0;  //39 / 163 = 0
    16'b00100111_10100100 : OUT <= 0;  //39 / 164 = 0
    16'b00100111_10100101 : OUT <= 0;  //39 / 165 = 0
    16'b00100111_10100110 : OUT <= 0;  //39 / 166 = 0
    16'b00100111_10100111 : OUT <= 0;  //39 / 167 = 0
    16'b00100111_10101000 : OUT <= 0;  //39 / 168 = 0
    16'b00100111_10101001 : OUT <= 0;  //39 / 169 = 0
    16'b00100111_10101010 : OUT <= 0;  //39 / 170 = 0
    16'b00100111_10101011 : OUT <= 0;  //39 / 171 = 0
    16'b00100111_10101100 : OUT <= 0;  //39 / 172 = 0
    16'b00100111_10101101 : OUT <= 0;  //39 / 173 = 0
    16'b00100111_10101110 : OUT <= 0;  //39 / 174 = 0
    16'b00100111_10101111 : OUT <= 0;  //39 / 175 = 0
    16'b00100111_10110000 : OUT <= 0;  //39 / 176 = 0
    16'b00100111_10110001 : OUT <= 0;  //39 / 177 = 0
    16'b00100111_10110010 : OUT <= 0;  //39 / 178 = 0
    16'b00100111_10110011 : OUT <= 0;  //39 / 179 = 0
    16'b00100111_10110100 : OUT <= 0;  //39 / 180 = 0
    16'b00100111_10110101 : OUT <= 0;  //39 / 181 = 0
    16'b00100111_10110110 : OUT <= 0;  //39 / 182 = 0
    16'b00100111_10110111 : OUT <= 0;  //39 / 183 = 0
    16'b00100111_10111000 : OUT <= 0;  //39 / 184 = 0
    16'b00100111_10111001 : OUT <= 0;  //39 / 185 = 0
    16'b00100111_10111010 : OUT <= 0;  //39 / 186 = 0
    16'b00100111_10111011 : OUT <= 0;  //39 / 187 = 0
    16'b00100111_10111100 : OUT <= 0;  //39 / 188 = 0
    16'b00100111_10111101 : OUT <= 0;  //39 / 189 = 0
    16'b00100111_10111110 : OUT <= 0;  //39 / 190 = 0
    16'b00100111_10111111 : OUT <= 0;  //39 / 191 = 0
    16'b00100111_11000000 : OUT <= 0;  //39 / 192 = 0
    16'b00100111_11000001 : OUT <= 0;  //39 / 193 = 0
    16'b00100111_11000010 : OUT <= 0;  //39 / 194 = 0
    16'b00100111_11000011 : OUT <= 0;  //39 / 195 = 0
    16'b00100111_11000100 : OUT <= 0;  //39 / 196 = 0
    16'b00100111_11000101 : OUT <= 0;  //39 / 197 = 0
    16'b00100111_11000110 : OUT <= 0;  //39 / 198 = 0
    16'b00100111_11000111 : OUT <= 0;  //39 / 199 = 0
    16'b00100111_11001000 : OUT <= 0;  //39 / 200 = 0
    16'b00100111_11001001 : OUT <= 0;  //39 / 201 = 0
    16'b00100111_11001010 : OUT <= 0;  //39 / 202 = 0
    16'b00100111_11001011 : OUT <= 0;  //39 / 203 = 0
    16'b00100111_11001100 : OUT <= 0;  //39 / 204 = 0
    16'b00100111_11001101 : OUT <= 0;  //39 / 205 = 0
    16'b00100111_11001110 : OUT <= 0;  //39 / 206 = 0
    16'b00100111_11001111 : OUT <= 0;  //39 / 207 = 0
    16'b00100111_11010000 : OUT <= 0;  //39 / 208 = 0
    16'b00100111_11010001 : OUT <= 0;  //39 / 209 = 0
    16'b00100111_11010010 : OUT <= 0;  //39 / 210 = 0
    16'b00100111_11010011 : OUT <= 0;  //39 / 211 = 0
    16'b00100111_11010100 : OUT <= 0;  //39 / 212 = 0
    16'b00100111_11010101 : OUT <= 0;  //39 / 213 = 0
    16'b00100111_11010110 : OUT <= 0;  //39 / 214 = 0
    16'b00100111_11010111 : OUT <= 0;  //39 / 215 = 0
    16'b00100111_11011000 : OUT <= 0;  //39 / 216 = 0
    16'b00100111_11011001 : OUT <= 0;  //39 / 217 = 0
    16'b00100111_11011010 : OUT <= 0;  //39 / 218 = 0
    16'b00100111_11011011 : OUT <= 0;  //39 / 219 = 0
    16'b00100111_11011100 : OUT <= 0;  //39 / 220 = 0
    16'b00100111_11011101 : OUT <= 0;  //39 / 221 = 0
    16'b00100111_11011110 : OUT <= 0;  //39 / 222 = 0
    16'b00100111_11011111 : OUT <= 0;  //39 / 223 = 0
    16'b00100111_11100000 : OUT <= 0;  //39 / 224 = 0
    16'b00100111_11100001 : OUT <= 0;  //39 / 225 = 0
    16'b00100111_11100010 : OUT <= 0;  //39 / 226 = 0
    16'b00100111_11100011 : OUT <= 0;  //39 / 227 = 0
    16'b00100111_11100100 : OUT <= 0;  //39 / 228 = 0
    16'b00100111_11100101 : OUT <= 0;  //39 / 229 = 0
    16'b00100111_11100110 : OUT <= 0;  //39 / 230 = 0
    16'b00100111_11100111 : OUT <= 0;  //39 / 231 = 0
    16'b00100111_11101000 : OUT <= 0;  //39 / 232 = 0
    16'b00100111_11101001 : OUT <= 0;  //39 / 233 = 0
    16'b00100111_11101010 : OUT <= 0;  //39 / 234 = 0
    16'b00100111_11101011 : OUT <= 0;  //39 / 235 = 0
    16'b00100111_11101100 : OUT <= 0;  //39 / 236 = 0
    16'b00100111_11101101 : OUT <= 0;  //39 / 237 = 0
    16'b00100111_11101110 : OUT <= 0;  //39 / 238 = 0
    16'b00100111_11101111 : OUT <= 0;  //39 / 239 = 0
    16'b00100111_11110000 : OUT <= 0;  //39 / 240 = 0
    16'b00100111_11110001 : OUT <= 0;  //39 / 241 = 0
    16'b00100111_11110010 : OUT <= 0;  //39 / 242 = 0
    16'b00100111_11110011 : OUT <= 0;  //39 / 243 = 0
    16'b00100111_11110100 : OUT <= 0;  //39 / 244 = 0
    16'b00100111_11110101 : OUT <= 0;  //39 / 245 = 0
    16'b00100111_11110110 : OUT <= 0;  //39 / 246 = 0
    16'b00100111_11110111 : OUT <= 0;  //39 / 247 = 0
    16'b00100111_11111000 : OUT <= 0;  //39 / 248 = 0
    16'b00100111_11111001 : OUT <= 0;  //39 / 249 = 0
    16'b00100111_11111010 : OUT <= 0;  //39 / 250 = 0
    16'b00100111_11111011 : OUT <= 0;  //39 / 251 = 0
    16'b00100111_11111100 : OUT <= 0;  //39 / 252 = 0
    16'b00100111_11111101 : OUT <= 0;  //39 / 253 = 0
    16'b00100111_11111110 : OUT <= 0;  //39 / 254 = 0
    16'b00100111_11111111 : OUT <= 0;  //39 / 255 = 0
    16'b00101000_00000000 : OUT <= 0;  //40 / 0 = 0
    16'b00101000_00000001 : OUT <= 40;  //40 / 1 = 40
    16'b00101000_00000010 : OUT <= 20;  //40 / 2 = 20
    16'b00101000_00000011 : OUT <= 13;  //40 / 3 = 13
    16'b00101000_00000100 : OUT <= 10;  //40 / 4 = 10
    16'b00101000_00000101 : OUT <= 8;  //40 / 5 = 8
    16'b00101000_00000110 : OUT <= 6;  //40 / 6 = 6
    16'b00101000_00000111 : OUT <= 5;  //40 / 7 = 5
    16'b00101000_00001000 : OUT <= 5;  //40 / 8 = 5
    16'b00101000_00001001 : OUT <= 4;  //40 / 9 = 4
    16'b00101000_00001010 : OUT <= 4;  //40 / 10 = 4
    16'b00101000_00001011 : OUT <= 3;  //40 / 11 = 3
    16'b00101000_00001100 : OUT <= 3;  //40 / 12 = 3
    16'b00101000_00001101 : OUT <= 3;  //40 / 13 = 3
    16'b00101000_00001110 : OUT <= 2;  //40 / 14 = 2
    16'b00101000_00001111 : OUT <= 2;  //40 / 15 = 2
    16'b00101000_00010000 : OUT <= 2;  //40 / 16 = 2
    16'b00101000_00010001 : OUT <= 2;  //40 / 17 = 2
    16'b00101000_00010010 : OUT <= 2;  //40 / 18 = 2
    16'b00101000_00010011 : OUT <= 2;  //40 / 19 = 2
    16'b00101000_00010100 : OUT <= 2;  //40 / 20 = 2
    16'b00101000_00010101 : OUT <= 1;  //40 / 21 = 1
    16'b00101000_00010110 : OUT <= 1;  //40 / 22 = 1
    16'b00101000_00010111 : OUT <= 1;  //40 / 23 = 1
    16'b00101000_00011000 : OUT <= 1;  //40 / 24 = 1
    16'b00101000_00011001 : OUT <= 1;  //40 / 25 = 1
    16'b00101000_00011010 : OUT <= 1;  //40 / 26 = 1
    16'b00101000_00011011 : OUT <= 1;  //40 / 27 = 1
    16'b00101000_00011100 : OUT <= 1;  //40 / 28 = 1
    16'b00101000_00011101 : OUT <= 1;  //40 / 29 = 1
    16'b00101000_00011110 : OUT <= 1;  //40 / 30 = 1
    16'b00101000_00011111 : OUT <= 1;  //40 / 31 = 1
    16'b00101000_00100000 : OUT <= 1;  //40 / 32 = 1
    16'b00101000_00100001 : OUT <= 1;  //40 / 33 = 1
    16'b00101000_00100010 : OUT <= 1;  //40 / 34 = 1
    16'b00101000_00100011 : OUT <= 1;  //40 / 35 = 1
    16'b00101000_00100100 : OUT <= 1;  //40 / 36 = 1
    16'b00101000_00100101 : OUT <= 1;  //40 / 37 = 1
    16'b00101000_00100110 : OUT <= 1;  //40 / 38 = 1
    16'b00101000_00100111 : OUT <= 1;  //40 / 39 = 1
    16'b00101000_00101000 : OUT <= 1;  //40 / 40 = 1
    16'b00101000_00101001 : OUT <= 0;  //40 / 41 = 0
    16'b00101000_00101010 : OUT <= 0;  //40 / 42 = 0
    16'b00101000_00101011 : OUT <= 0;  //40 / 43 = 0
    16'b00101000_00101100 : OUT <= 0;  //40 / 44 = 0
    16'b00101000_00101101 : OUT <= 0;  //40 / 45 = 0
    16'b00101000_00101110 : OUT <= 0;  //40 / 46 = 0
    16'b00101000_00101111 : OUT <= 0;  //40 / 47 = 0
    16'b00101000_00110000 : OUT <= 0;  //40 / 48 = 0
    16'b00101000_00110001 : OUT <= 0;  //40 / 49 = 0
    16'b00101000_00110010 : OUT <= 0;  //40 / 50 = 0
    16'b00101000_00110011 : OUT <= 0;  //40 / 51 = 0
    16'b00101000_00110100 : OUT <= 0;  //40 / 52 = 0
    16'b00101000_00110101 : OUT <= 0;  //40 / 53 = 0
    16'b00101000_00110110 : OUT <= 0;  //40 / 54 = 0
    16'b00101000_00110111 : OUT <= 0;  //40 / 55 = 0
    16'b00101000_00111000 : OUT <= 0;  //40 / 56 = 0
    16'b00101000_00111001 : OUT <= 0;  //40 / 57 = 0
    16'b00101000_00111010 : OUT <= 0;  //40 / 58 = 0
    16'b00101000_00111011 : OUT <= 0;  //40 / 59 = 0
    16'b00101000_00111100 : OUT <= 0;  //40 / 60 = 0
    16'b00101000_00111101 : OUT <= 0;  //40 / 61 = 0
    16'b00101000_00111110 : OUT <= 0;  //40 / 62 = 0
    16'b00101000_00111111 : OUT <= 0;  //40 / 63 = 0
    16'b00101000_01000000 : OUT <= 0;  //40 / 64 = 0
    16'b00101000_01000001 : OUT <= 0;  //40 / 65 = 0
    16'b00101000_01000010 : OUT <= 0;  //40 / 66 = 0
    16'b00101000_01000011 : OUT <= 0;  //40 / 67 = 0
    16'b00101000_01000100 : OUT <= 0;  //40 / 68 = 0
    16'b00101000_01000101 : OUT <= 0;  //40 / 69 = 0
    16'b00101000_01000110 : OUT <= 0;  //40 / 70 = 0
    16'b00101000_01000111 : OUT <= 0;  //40 / 71 = 0
    16'b00101000_01001000 : OUT <= 0;  //40 / 72 = 0
    16'b00101000_01001001 : OUT <= 0;  //40 / 73 = 0
    16'b00101000_01001010 : OUT <= 0;  //40 / 74 = 0
    16'b00101000_01001011 : OUT <= 0;  //40 / 75 = 0
    16'b00101000_01001100 : OUT <= 0;  //40 / 76 = 0
    16'b00101000_01001101 : OUT <= 0;  //40 / 77 = 0
    16'b00101000_01001110 : OUT <= 0;  //40 / 78 = 0
    16'b00101000_01001111 : OUT <= 0;  //40 / 79 = 0
    16'b00101000_01010000 : OUT <= 0;  //40 / 80 = 0
    16'b00101000_01010001 : OUT <= 0;  //40 / 81 = 0
    16'b00101000_01010010 : OUT <= 0;  //40 / 82 = 0
    16'b00101000_01010011 : OUT <= 0;  //40 / 83 = 0
    16'b00101000_01010100 : OUT <= 0;  //40 / 84 = 0
    16'b00101000_01010101 : OUT <= 0;  //40 / 85 = 0
    16'b00101000_01010110 : OUT <= 0;  //40 / 86 = 0
    16'b00101000_01010111 : OUT <= 0;  //40 / 87 = 0
    16'b00101000_01011000 : OUT <= 0;  //40 / 88 = 0
    16'b00101000_01011001 : OUT <= 0;  //40 / 89 = 0
    16'b00101000_01011010 : OUT <= 0;  //40 / 90 = 0
    16'b00101000_01011011 : OUT <= 0;  //40 / 91 = 0
    16'b00101000_01011100 : OUT <= 0;  //40 / 92 = 0
    16'b00101000_01011101 : OUT <= 0;  //40 / 93 = 0
    16'b00101000_01011110 : OUT <= 0;  //40 / 94 = 0
    16'b00101000_01011111 : OUT <= 0;  //40 / 95 = 0
    16'b00101000_01100000 : OUT <= 0;  //40 / 96 = 0
    16'b00101000_01100001 : OUT <= 0;  //40 / 97 = 0
    16'b00101000_01100010 : OUT <= 0;  //40 / 98 = 0
    16'b00101000_01100011 : OUT <= 0;  //40 / 99 = 0
    16'b00101000_01100100 : OUT <= 0;  //40 / 100 = 0
    16'b00101000_01100101 : OUT <= 0;  //40 / 101 = 0
    16'b00101000_01100110 : OUT <= 0;  //40 / 102 = 0
    16'b00101000_01100111 : OUT <= 0;  //40 / 103 = 0
    16'b00101000_01101000 : OUT <= 0;  //40 / 104 = 0
    16'b00101000_01101001 : OUT <= 0;  //40 / 105 = 0
    16'b00101000_01101010 : OUT <= 0;  //40 / 106 = 0
    16'b00101000_01101011 : OUT <= 0;  //40 / 107 = 0
    16'b00101000_01101100 : OUT <= 0;  //40 / 108 = 0
    16'b00101000_01101101 : OUT <= 0;  //40 / 109 = 0
    16'b00101000_01101110 : OUT <= 0;  //40 / 110 = 0
    16'b00101000_01101111 : OUT <= 0;  //40 / 111 = 0
    16'b00101000_01110000 : OUT <= 0;  //40 / 112 = 0
    16'b00101000_01110001 : OUT <= 0;  //40 / 113 = 0
    16'b00101000_01110010 : OUT <= 0;  //40 / 114 = 0
    16'b00101000_01110011 : OUT <= 0;  //40 / 115 = 0
    16'b00101000_01110100 : OUT <= 0;  //40 / 116 = 0
    16'b00101000_01110101 : OUT <= 0;  //40 / 117 = 0
    16'b00101000_01110110 : OUT <= 0;  //40 / 118 = 0
    16'b00101000_01110111 : OUT <= 0;  //40 / 119 = 0
    16'b00101000_01111000 : OUT <= 0;  //40 / 120 = 0
    16'b00101000_01111001 : OUT <= 0;  //40 / 121 = 0
    16'b00101000_01111010 : OUT <= 0;  //40 / 122 = 0
    16'b00101000_01111011 : OUT <= 0;  //40 / 123 = 0
    16'b00101000_01111100 : OUT <= 0;  //40 / 124 = 0
    16'b00101000_01111101 : OUT <= 0;  //40 / 125 = 0
    16'b00101000_01111110 : OUT <= 0;  //40 / 126 = 0
    16'b00101000_01111111 : OUT <= 0;  //40 / 127 = 0
    16'b00101000_10000000 : OUT <= 0;  //40 / 128 = 0
    16'b00101000_10000001 : OUT <= 0;  //40 / 129 = 0
    16'b00101000_10000010 : OUT <= 0;  //40 / 130 = 0
    16'b00101000_10000011 : OUT <= 0;  //40 / 131 = 0
    16'b00101000_10000100 : OUT <= 0;  //40 / 132 = 0
    16'b00101000_10000101 : OUT <= 0;  //40 / 133 = 0
    16'b00101000_10000110 : OUT <= 0;  //40 / 134 = 0
    16'b00101000_10000111 : OUT <= 0;  //40 / 135 = 0
    16'b00101000_10001000 : OUT <= 0;  //40 / 136 = 0
    16'b00101000_10001001 : OUT <= 0;  //40 / 137 = 0
    16'b00101000_10001010 : OUT <= 0;  //40 / 138 = 0
    16'b00101000_10001011 : OUT <= 0;  //40 / 139 = 0
    16'b00101000_10001100 : OUT <= 0;  //40 / 140 = 0
    16'b00101000_10001101 : OUT <= 0;  //40 / 141 = 0
    16'b00101000_10001110 : OUT <= 0;  //40 / 142 = 0
    16'b00101000_10001111 : OUT <= 0;  //40 / 143 = 0
    16'b00101000_10010000 : OUT <= 0;  //40 / 144 = 0
    16'b00101000_10010001 : OUT <= 0;  //40 / 145 = 0
    16'b00101000_10010010 : OUT <= 0;  //40 / 146 = 0
    16'b00101000_10010011 : OUT <= 0;  //40 / 147 = 0
    16'b00101000_10010100 : OUT <= 0;  //40 / 148 = 0
    16'b00101000_10010101 : OUT <= 0;  //40 / 149 = 0
    16'b00101000_10010110 : OUT <= 0;  //40 / 150 = 0
    16'b00101000_10010111 : OUT <= 0;  //40 / 151 = 0
    16'b00101000_10011000 : OUT <= 0;  //40 / 152 = 0
    16'b00101000_10011001 : OUT <= 0;  //40 / 153 = 0
    16'b00101000_10011010 : OUT <= 0;  //40 / 154 = 0
    16'b00101000_10011011 : OUT <= 0;  //40 / 155 = 0
    16'b00101000_10011100 : OUT <= 0;  //40 / 156 = 0
    16'b00101000_10011101 : OUT <= 0;  //40 / 157 = 0
    16'b00101000_10011110 : OUT <= 0;  //40 / 158 = 0
    16'b00101000_10011111 : OUT <= 0;  //40 / 159 = 0
    16'b00101000_10100000 : OUT <= 0;  //40 / 160 = 0
    16'b00101000_10100001 : OUT <= 0;  //40 / 161 = 0
    16'b00101000_10100010 : OUT <= 0;  //40 / 162 = 0
    16'b00101000_10100011 : OUT <= 0;  //40 / 163 = 0
    16'b00101000_10100100 : OUT <= 0;  //40 / 164 = 0
    16'b00101000_10100101 : OUT <= 0;  //40 / 165 = 0
    16'b00101000_10100110 : OUT <= 0;  //40 / 166 = 0
    16'b00101000_10100111 : OUT <= 0;  //40 / 167 = 0
    16'b00101000_10101000 : OUT <= 0;  //40 / 168 = 0
    16'b00101000_10101001 : OUT <= 0;  //40 / 169 = 0
    16'b00101000_10101010 : OUT <= 0;  //40 / 170 = 0
    16'b00101000_10101011 : OUT <= 0;  //40 / 171 = 0
    16'b00101000_10101100 : OUT <= 0;  //40 / 172 = 0
    16'b00101000_10101101 : OUT <= 0;  //40 / 173 = 0
    16'b00101000_10101110 : OUT <= 0;  //40 / 174 = 0
    16'b00101000_10101111 : OUT <= 0;  //40 / 175 = 0
    16'b00101000_10110000 : OUT <= 0;  //40 / 176 = 0
    16'b00101000_10110001 : OUT <= 0;  //40 / 177 = 0
    16'b00101000_10110010 : OUT <= 0;  //40 / 178 = 0
    16'b00101000_10110011 : OUT <= 0;  //40 / 179 = 0
    16'b00101000_10110100 : OUT <= 0;  //40 / 180 = 0
    16'b00101000_10110101 : OUT <= 0;  //40 / 181 = 0
    16'b00101000_10110110 : OUT <= 0;  //40 / 182 = 0
    16'b00101000_10110111 : OUT <= 0;  //40 / 183 = 0
    16'b00101000_10111000 : OUT <= 0;  //40 / 184 = 0
    16'b00101000_10111001 : OUT <= 0;  //40 / 185 = 0
    16'b00101000_10111010 : OUT <= 0;  //40 / 186 = 0
    16'b00101000_10111011 : OUT <= 0;  //40 / 187 = 0
    16'b00101000_10111100 : OUT <= 0;  //40 / 188 = 0
    16'b00101000_10111101 : OUT <= 0;  //40 / 189 = 0
    16'b00101000_10111110 : OUT <= 0;  //40 / 190 = 0
    16'b00101000_10111111 : OUT <= 0;  //40 / 191 = 0
    16'b00101000_11000000 : OUT <= 0;  //40 / 192 = 0
    16'b00101000_11000001 : OUT <= 0;  //40 / 193 = 0
    16'b00101000_11000010 : OUT <= 0;  //40 / 194 = 0
    16'b00101000_11000011 : OUT <= 0;  //40 / 195 = 0
    16'b00101000_11000100 : OUT <= 0;  //40 / 196 = 0
    16'b00101000_11000101 : OUT <= 0;  //40 / 197 = 0
    16'b00101000_11000110 : OUT <= 0;  //40 / 198 = 0
    16'b00101000_11000111 : OUT <= 0;  //40 / 199 = 0
    16'b00101000_11001000 : OUT <= 0;  //40 / 200 = 0
    16'b00101000_11001001 : OUT <= 0;  //40 / 201 = 0
    16'b00101000_11001010 : OUT <= 0;  //40 / 202 = 0
    16'b00101000_11001011 : OUT <= 0;  //40 / 203 = 0
    16'b00101000_11001100 : OUT <= 0;  //40 / 204 = 0
    16'b00101000_11001101 : OUT <= 0;  //40 / 205 = 0
    16'b00101000_11001110 : OUT <= 0;  //40 / 206 = 0
    16'b00101000_11001111 : OUT <= 0;  //40 / 207 = 0
    16'b00101000_11010000 : OUT <= 0;  //40 / 208 = 0
    16'b00101000_11010001 : OUT <= 0;  //40 / 209 = 0
    16'b00101000_11010010 : OUT <= 0;  //40 / 210 = 0
    16'b00101000_11010011 : OUT <= 0;  //40 / 211 = 0
    16'b00101000_11010100 : OUT <= 0;  //40 / 212 = 0
    16'b00101000_11010101 : OUT <= 0;  //40 / 213 = 0
    16'b00101000_11010110 : OUT <= 0;  //40 / 214 = 0
    16'b00101000_11010111 : OUT <= 0;  //40 / 215 = 0
    16'b00101000_11011000 : OUT <= 0;  //40 / 216 = 0
    16'b00101000_11011001 : OUT <= 0;  //40 / 217 = 0
    16'b00101000_11011010 : OUT <= 0;  //40 / 218 = 0
    16'b00101000_11011011 : OUT <= 0;  //40 / 219 = 0
    16'b00101000_11011100 : OUT <= 0;  //40 / 220 = 0
    16'b00101000_11011101 : OUT <= 0;  //40 / 221 = 0
    16'b00101000_11011110 : OUT <= 0;  //40 / 222 = 0
    16'b00101000_11011111 : OUT <= 0;  //40 / 223 = 0
    16'b00101000_11100000 : OUT <= 0;  //40 / 224 = 0
    16'b00101000_11100001 : OUT <= 0;  //40 / 225 = 0
    16'b00101000_11100010 : OUT <= 0;  //40 / 226 = 0
    16'b00101000_11100011 : OUT <= 0;  //40 / 227 = 0
    16'b00101000_11100100 : OUT <= 0;  //40 / 228 = 0
    16'b00101000_11100101 : OUT <= 0;  //40 / 229 = 0
    16'b00101000_11100110 : OUT <= 0;  //40 / 230 = 0
    16'b00101000_11100111 : OUT <= 0;  //40 / 231 = 0
    16'b00101000_11101000 : OUT <= 0;  //40 / 232 = 0
    16'b00101000_11101001 : OUT <= 0;  //40 / 233 = 0
    16'b00101000_11101010 : OUT <= 0;  //40 / 234 = 0
    16'b00101000_11101011 : OUT <= 0;  //40 / 235 = 0
    16'b00101000_11101100 : OUT <= 0;  //40 / 236 = 0
    16'b00101000_11101101 : OUT <= 0;  //40 / 237 = 0
    16'b00101000_11101110 : OUT <= 0;  //40 / 238 = 0
    16'b00101000_11101111 : OUT <= 0;  //40 / 239 = 0
    16'b00101000_11110000 : OUT <= 0;  //40 / 240 = 0
    16'b00101000_11110001 : OUT <= 0;  //40 / 241 = 0
    16'b00101000_11110010 : OUT <= 0;  //40 / 242 = 0
    16'b00101000_11110011 : OUT <= 0;  //40 / 243 = 0
    16'b00101000_11110100 : OUT <= 0;  //40 / 244 = 0
    16'b00101000_11110101 : OUT <= 0;  //40 / 245 = 0
    16'b00101000_11110110 : OUT <= 0;  //40 / 246 = 0
    16'b00101000_11110111 : OUT <= 0;  //40 / 247 = 0
    16'b00101000_11111000 : OUT <= 0;  //40 / 248 = 0
    16'b00101000_11111001 : OUT <= 0;  //40 / 249 = 0
    16'b00101000_11111010 : OUT <= 0;  //40 / 250 = 0
    16'b00101000_11111011 : OUT <= 0;  //40 / 251 = 0
    16'b00101000_11111100 : OUT <= 0;  //40 / 252 = 0
    16'b00101000_11111101 : OUT <= 0;  //40 / 253 = 0
    16'b00101000_11111110 : OUT <= 0;  //40 / 254 = 0
    16'b00101000_11111111 : OUT <= 0;  //40 / 255 = 0
    16'b00101001_00000000 : OUT <= 0;  //41 / 0 = 0
    16'b00101001_00000001 : OUT <= 41;  //41 / 1 = 41
    16'b00101001_00000010 : OUT <= 20;  //41 / 2 = 20
    16'b00101001_00000011 : OUT <= 13;  //41 / 3 = 13
    16'b00101001_00000100 : OUT <= 10;  //41 / 4 = 10
    16'b00101001_00000101 : OUT <= 8;  //41 / 5 = 8
    16'b00101001_00000110 : OUT <= 6;  //41 / 6 = 6
    16'b00101001_00000111 : OUT <= 5;  //41 / 7 = 5
    16'b00101001_00001000 : OUT <= 5;  //41 / 8 = 5
    16'b00101001_00001001 : OUT <= 4;  //41 / 9 = 4
    16'b00101001_00001010 : OUT <= 4;  //41 / 10 = 4
    16'b00101001_00001011 : OUT <= 3;  //41 / 11 = 3
    16'b00101001_00001100 : OUT <= 3;  //41 / 12 = 3
    16'b00101001_00001101 : OUT <= 3;  //41 / 13 = 3
    16'b00101001_00001110 : OUT <= 2;  //41 / 14 = 2
    16'b00101001_00001111 : OUT <= 2;  //41 / 15 = 2
    16'b00101001_00010000 : OUT <= 2;  //41 / 16 = 2
    16'b00101001_00010001 : OUT <= 2;  //41 / 17 = 2
    16'b00101001_00010010 : OUT <= 2;  //41 / 18 = 2
    16'b00101001_00010011 : OUT <= 2;  //41 / 19 = 2
    16'b00101001_00010100 : OUT <= 2;  //41 / 20 = 2
    16'b00101001_00010101 : OUT <= 1;  //41 / 21 = 1
    16'b00101001_00010110 : OUT <= 1;  //41 / 22 = 1
    16'b00101001_00010111 : OUT <= 1;  //41 / 23 = 1
    16'b00101001_00011000 : OUT <= 1;  //41 / 24 = 1
    16'b00101001_00011001 : OUT <= 1;  //41 / 25 = 1
    16'b00101001_00011010 : OUT <= 1;  //41 / 26 = 1
    16'b00101001_00011011 : OUT <= 1;  //41 / 27 = 1
    16'b00101001_00011100 : OUT <= 1;  //41 / 28 = 1
    16'b00101001_00011101 : OUT <= 1;  //41 / 29 = 1
    16'b00101001_00011110 : OUT <= 1;  //41 / 30 = 1
    16'b00101001_00011111 : OUT <= 1;  //41 / 31 = 1
    16'b00101001_00100000 : OUT <= 1;  //41 / 32 = 1
    16'b00101001_00100001 : OUT <= 1;  //41 / 33 = 1
    16'b00101001_00100010 : OUT <= 1;  //41 / 34 = 1
    16'b00101001_00100011 : OUT <= 1;  //41 / 35 = 1
    16'b00101001_00100100 : OUT <= 1;  //41 / 36 = 1
    16'b00101001_00100101 : OUT <= 1;  //41 / 37 = 1
    16'b00101001_00100110 : OUT <= 1;  //41 / 38 = 1
    16'b00101001_00100111 : OUT <= 1;  //41 / 39 = 1
    16'b00101001_00101000 : OUT <= 1;  //41 / 40 = 1
    16'b00101001_00101001 : OUT <= 1;  //41 / 41 = 1
    16'b00101001_00101010 : OUT <= 0;  //41 / 42 = 0
    16'b00101001_00101011 : OUT <= 0;  //41 / 43 = 0
    16'b00101001_00101100 : OUT <= 0;  //41 / 44 = 0
    16'b00101001_00101101 : OUT <= 0;  //41 / 45 = 0
    16'b00101001_00101110 : OUT <= 0;  //41 / 46 = 0
    16'b00101001_00101111 : OUT <= 0;  //41 / 47 = 0
    16'b00101001_00110000 : OUT <= 0;  //41 / 48 = 0
    16'b00101001_00110001 : OUT <= 0;  //41 / 49 = 0
    16'b00101001_00110010 : OUT <= 0;  //41 / 50 = 0
    16'b00101001_00110011 : OUT <= 0;  //41 / 51 = 0
    16'b00101001_00110100 : OUT <= 0;  //41 / 52 = 0
    16'b00101001_00110101 : OUT <= 0;  //41 / 53 = 0
    16'b00101001_00110110 : OUT <= 0;  //41 / 54 = 0
    16'b00101001_00110111 : OUT <= 0;  //41 / 55 = 0
    16'b00101001_00111000 : OUT <= 0;  //41 / 56 = 0
    16'b00101001_00111001 : OUT <= 0;  //41 / 57 = 0
    16'b00101001_00111010 : OUT <= 0;  //41 / 58 = 0
    16'b00101001_00111011 : OUT <= 0;  //41 / 59 = 0
    16'b00101001_00111100 : OUT <= 0;  //41 / 60 = 0
    16'b00101001_00111101 : OUT <= 0;  //41 / 61 = 0
    16'b00101001_00111110 : OUT <= 0;  //41 / 62 = 0
    16'b00101001_00111111 : OUT <= 0;  //41 / 63 = 0
    16'b00101001_01000000 : OUT <= 0;  //41 / 64 = 0
    16'b00101001_01000001 : OUT <= 0;  //41 / 65 = 0
    16'b00101001_01000010 : OUT <= 0;  //41 / 66 = 0
    16'b00101001_01000011 : OUT <= 0;  //41 / 67 = 0
    16'b00101001_01000100 : OUT <= 0;  //41 / 68 = 0
    16'b00101001_01000101 : OUT <= 0;  //41 / 69 = 0
    16'b00101001_01000110 : OUT <= 0;  //41 / 70 = 0
    16'b00101001_01000111 : OUT <= 0;  //41 / 71 = 0
    16'b00101001_01001000 : OUT <= 0;  //41 / 72 = 0
    16'b00101001_01001001 : OUT <= 0;  //41 / 73 = 0
    16'b00101001_01001010 : OUT <= 0;  //41 / 74 = 0
    16'b00101001_01001011 : OUT <= 0;  //41 / 75 = 0
    16'b00101001_01001100 : OUT <= 0;  //41 / 76 = 0
    16'b00101001_01001101 : OUT <= 0;  //41 / 77 = 0
    16'b00101001_01001110 : OUT <= 0;  //41 / 78 = 0
    16'b00101001_01001111 : OUT <= 0;  //41 / 79 = 0
    16'b00101001_01010000 : OUT <= 0;  //41 / 80 = 0
    16'b00101001_01010001 : OUT <= 0;  //41 / 81 = 0
    16'b00101001_01010010 : OUT <= 0;  //41 / 82 = 0
    16'b00101001_01010011 : OUT <= 0;  //41 / 83 = 0
    16'b00101001_01010100 : OUT <= 0;  //41 / 84 = 0
    16'b00101001_01010101 : OUT <= 0;  //41 / 85 = 0
    16'b00101001_01010110 : OUT <= 0;  //41 / 86 = 0
    16'b00101001_01010111 : OUT <= 0;  //41 / 87 = 0
    16'b00101001_01011000 : OUT <= 0;  //41 / 88 = 0
    16'b00101001_01011001 : OUT <= 0;  //41 / 89 = 0
    16'b00101001_01011010 : OUT <= 0;  //41 / 90 = 0
    16'b00101001_01011011 : OUT <= 0;  //41 / 91 = 0
    16'b00101001_01011100 : OUT <= 0;  //41 / 92 = 0
    16'b00101001_01011101 : OUT <= 0;  //41 / 93 = 0
    16'b00101001_01011110 : OUT <= 0;  //41 / 94 = 0
    16'b00101001_01011111 : OUT <= 0;  //41 / 95 = 0
    16'b00101001_01100000 : OUT <= 0;  //41 / 96 = 0
    16'b00101001_01100001 : OUT <= 0;  //41 / 97 = 0
    16'b00101001_01100010 : OUT <= 0;  //41 / 98 = 0
    16'b00101001_01100011 : OUT <= 0;  //41 / 99 = 0
    16'b00101001_01100100 : OUT <= 0;  //41 / 100 = 0
    16'b00101001_01100101 : OUT <= 0;  //41 / 101 = 0
    16'b00101001_01100110 : OUT <= 0;  //41 / 102 = 0
    16'b00101001_01100111 : OUT <= 0;  //41 / 103 = 0
    16'b00101001_01101000 : OUT <= 0;  //41 / 104 = 0
    16'b00101001_01101001 : OUT <= 0;  //41 / 105 = 0
    16'b00101001_01101010 : OUT <= 0;  //41 / 106 = 0
    16'b00101001_01101011 : OUT <= 0;  //41 / 107 = 0
    16'b00101001_01101100 : OUT <= 0;  //41 / 108 = 0
    16'b00101001_01101101 : OUT <= 0;  //41 / 109 = 0
    16'b00101001_01101110 : OUT <= 0;  //41 / 110 = 0
    16'b00101001_01101111 : OUT <= 0;  //41 / 111 = 0
    16'b00101001_01110000 : OUT <= 0;  //41 / 112 = 0
    16'b00101001_01110001 : OUT <= 0;  //41 / 113 = 0
    16'b00101001_01110010 : OUT <= 0;  //41 / 114 = 0
    16'b00101001_01110011 : OUT <= 0;  //41 / 115 = 0
    16'b00101001_01110100 : OUT <= 0;  //41 / 116 = 0
    16'b00101001_01110101 : OUT <= 0;  //41 / 117 = 0
    16'b00101001_01110110 : OUT <= 0;  //41 / 118 = 0
    16'b00101001_01110111 : OUT <= 0;  //41 / 119 = 0
    16'b00101001_01111000 : OUT <= 0;  //41 / 120 = 0
    16'b00101001_01111001 : OUT <= 0;  //41 / 121 = 0
    16'b00101001_01111010 : OUT <= 0;  //41 / 122 = 0
    16'b00101001_01111011 : OUT <= 0;  //41 / 123 = 0
    16'b00101001_01111100 : OUT <= 0;  //41 / 124 = 0
    16'b00101001_01111101 : OUT <= 0;  //41 / 125 = 0
    16'b00101001_01111110 : OUT <= 0;  //41 / 126 = 0
    16'b00101001_01111111 : OUT <= 0;  //41 / 127 = 0
    16'b00101001_10000000 : OUT <= 0;  //41 / 128 = 0
    16'b00101001_10000001 : OUT <= 0;  //41 / 129 = 0
    16'b00101001_10000010 : OUT <= 0;  //41 / 130 = 0
    16'b00101001_10000011 : OUT <= 0;  //41 / 131 = 0
    16'b00101001_10000100 : OUT <= 0;  //41 / 132 = 0
    16'b00101001_10000101 : OUT <= 0;  //41 / 133 = 0
    16'b00101001_10000110 : OUT <= 0;  //41 / 134 = 0
    16'b00101001_10000111 : OUT <= 0;  //41 / 135 = 0
    16'b00101001_10001000 : OUT <= 0;  //41 / 136 = 0
    16'b00101001_10001001 : OUT <= 0;  //41 / 137 = 0
    16'b00101001_10001010 : OUT <= 0;  //41 / 138 = 0
    16'b00101001_10001011 : OUT <= 0;  //41 / 139 = 0
    16'b00101001_10001100 : OUT <= 0;  //41 / 140 = 0
    16'b00101001_10001101 : OUT <= 0;  //41 / 141 = 0
    16'b00101001_10001110 : OUT <= 0;  //41 / 142 = 0
    16'b00101001_10001111 : OUT <= 0;  //41 / 143 = 0
    16'b00101001_10010000 : OUT <= 0;  //41 / 144 = 0
    16'b00101001_10010001 : OUT <= 0;  //41 / 145 = 0
    16'b00101001_10010010 : OUT <= 0;  //41 / 146 = 0
    16'b00101001_10010011 : OUT <= 0;  //41 / 147 = 0
    16'b00101001_10010100 : OUT <= 0;  //41 / 148 = 0
    16'b00101001_10010101 : OUT <= 0;  //41 / 149 = 0
    16'b00101001_10010110 : OUT <= 0;  //41 / 150 = 0
    16'b00101001_10010111 : OUT <= 0;  //41 / 151 = 0
    16'b00101001_10011000 : OUT <= 0;  //41 / 152 = 0
    16'b00101001_10011001 : OUT <= 0;  //41 / 153 = 0
    16'b00101001_10011010 : OUT <= 0;  //41 / 154 = 0
    16'b00101001_10011011 : OUT <= 0;  //41 / 155 = 0
    16'b00101001_10011100 : OUT <= 0;  //41 / 156 = 0
    16'b00101001_10011101 : OUT <= 0;  //41 / 157 = 0
    16'b00101001_10011110 : OUT <= 0;  //41 / 158 = 0
    16'b00101001_10011111 : OUT <= 0;  //41 / 159 = 0
    16'b00101001_10100000 : OUT <= 0;  //41 / 160 = 0
    16'b00101001_10100001 : OUT <= 0;  //41 / 161 = 0
    16'b00101001_10100010 : OUT <= 0;  //41 / 162 = 0
    16'b00101001_10100011 : OUT <= 0;  //41 / 163 = 0
    16'b00101001_10100100 : OUT <= 0;  //41 / 164 = 0
    16'b00101001_10100101 : OUT <= 0;  //41 / 165 = 0
    16'b00101001_10100110 : OUT <= 0;  //41 / 166 = 0
    16'b00101001_10100111 : OUT <= 0;  //41 / 167 = 0
    16'b00101001_10101000 : OUT <= 0;  //41 / 168 = 0
    16'b00101001_10101001 : OUT <= 0;  //41 / 169 = 0
    16'b00101001_10101010 : OUT <= 0;  //41 / 170 = 0
    16'b00101001_10101011 : OUT <= 0;  //41 / 171 = 0
    16'b00101001_10101100 : OUT <= 0;  //41 / 172 = 0
    16'b00101001_10101101 : OUT <= 0;  //41 / 173 = 0
    16'b00101001_10101110 : OUT <= 0;  //41 / 174 = 0
    16'b00101001_10101111 : OUT <= 0;  //41 / 175 = 0
    16'b00101001_10110000 : OUT <= 0;  //41 / 176 = 0
    16'b00101001_10110001 : OUT <= 0;  //41 / 177 = 0
    16'b00101001_10110010 : OUT <= 0;  //41 / 178 = 0
    16'b00101001_10110011 : OUT <= 0;  //41 / 179 = 0
    16'b00101001_10110100 : OUT <= 0;  //41 / 180 = 0
    16'b00101001_10110101 : OUT <= 0;  //41 / 181 = 0
    16'b00101001_10110110 : OUT <= 0;  //41 / 182 = 0
    16'b00101001_10110111 : OUT <= 0;  //41 / 183 = 0
    16'b00101001_10111000 : OUT <= 0;  //41 / 184 = 0
    16'b00101001_10111001 : OUT <= 0;  //41 / 185 = 0
    16'b00101001_10111010 : OUT <= 0;  //41 / 186 = 0
    16'b00101001_10111011 : OUT <= 0;  //41 / 187 = 0
    16'b00101001_10111100 : OUT <= 0;  //41 / 188 = 0
    16'b00101001_10111101 : OUT <= 0;  //41 / 189 = 0
    16'b00101001_10111110 : OUT <= 0;  //41 / 190 = 0
    16'b00101001_10111111 : OUT <= 0;  //41 / 191 = 0
    16'b00101001_11000000 : OUT <= 0;  //41 / 192 = 0
    16'b00101001_11000001 : OUT <= 0;  //41 / 193 = 0
    16'b00101001_11000010 : OUT <= 0;  //41 / 194 = 0
    16'b00101001_11000011 : OUT <= 0;  //41 / 195 = 0
    16'b00101001_11000100 : OUT <= 0;  //41 / 196 = 0
    16'b00101001_11000101 : OUT <= 0;  //41 / 197 = 0
    16'b00101001_11000110 : OUT <= 0;  //41 / 198 = 0
    16'b00101001_11000111 : OUT <= 0;  //41 / 199 = 0
    16'b00101001_11001000 : OUT <= 0;  //41 / 200 = 0
    16'b00101001_11001001 : OUT <= 0;  //41 / 201 = 0
    16'b00101001_11001010 : OUT <= 0;  //41 / 202 = 0
    16'b00101001_11001011 : OUT <= 0;  //41 / 203 = 0
    16'b00101001_11001100 : OUT <= 0;  //41 / 204 = 0
    16'b00101001_11001101 : OUT <= 0;  //41 / 205 = 0
    16'b00101001_11001110 : OUT <= 0;  //41 / 206 = 0
    16'b00101001_11001111 : OUT <= 0;  //41 / 207 = 0
    16'b00101001_11010000 : OUT <= 0;  //41 / 208 = 0
    16'b00101001_11010001 : OUT <= 0;  //41 / 209 = 0
    16'b00101001_11010010 : OUT <= 0;  //41 / 210 = 0
    16'b00101001_11010011 : OUT <= 0;  //41 / 211 = 0
    16'b00101001_11010100 : OUT <= 0;  //41 / 212 = 0
    16'b00101001_11010101 : OUT <= 0;  //41 / 213 = 0
    16'b00101001_11010110 : OUT <= 0;  //41 / 214 = 0
    16'b00101001_11010111 : OUT <= 0;  //41 / 215 = 0
    16'b00101001_11011000 : OUT <= 0;  //41 / 216 = 0
    16'b00101001_11011001 : OUT <= 0;  //41 / 217 = 0
    16'b00101001_11011010 : OUT <= 0;  //41 / 218 = 0
    16'b00101001_11011011 : OUT <= 0;  //41 / 219 = 0
    16'b00101001_11011100 : OUT <= 0;  //41 / 220 = 0
    16'b00101001_11011101 : OUT <= 0;  //41 / 221 = 0
    16'b00101001_11011110 : OUT <= 0;  //41 / 222 = 0
    16'b00101001_11011111 : OUT <= 0;  //41 / 223 = 0
    16'b00101001_11100000 : OUT <= 0;  //41 / 224 = 0
    16'b00101001_11100001 : OUT <= 0;  //41 / 225 = 0
    16'b00101001_11100010 : OUT <= 0;  //41 / 226 = 0
    16'b00101001_11100011 : OUT <= 0;  //41 / 227 = 0
    16'b00101001_11100100 : OUT <= 0;  //41 / 228 = 0
    16'b00101001_11100101 : OUT <= 0;  //41 / 229 = 0
    16'b00101001_11100110 : OUT <= 0;  //41 / 230 = 0
    16'b00101001_11100111 : OUT <= 0;  //41 / 231 = 0
    16'b00101001_11101000 : OUT <= 0;  //41 / 232 = 0
    16'b00101001_11101001 : OUT <= 0;  //41 / 233 = 0
    16'b00101001_11101010 : OUT <= 0;  //41 / 234 = 0
    16'b00101001_11101011 : OUT <= 0;  //41 / 235 = 0
    16'b00101001_11101100 : OUT <= 0;  //41 / 236 = 0
    16'b00101001_11101101 : OUT <= 0;  //41 / 237 = 0
    16'b00101001_11101110 : OUT <= 0;  //41 / 238 = 0
    16'b00101001_11101111 : OUT <= 0;  //41 / 239 = 0
    16'b00101001_11110000 : OUT <= 0;  //41 / 240 = 0
    16'b00101001_11110001 : OUT <= 0;  //41 / 241 = 0
    16'b00101001_11110010 : OUT <= 0;  //41 / 242 = 0
    16'b00101001_11110011 : OUT <= 0;  //41 / 243 = 0
    16'b00101001_11110100 : OUT <= 0;  //41 / 244 = 0
    16'b00101001_11110101 : OUT <= 0;  //41 / 245 = 0
    16'b00101001_11110110 : OUT <= 0;  //41 / 246 = 0
    16'b00101001_11110111 : OUT <= 0;  //41 / 247 = 0
    16'b00101001_11111000 : OUT <= 0;  //41 / 248 = 0
    16'b00101001_11111001 : OUT <= 0;  //41 / 249 = 0
    16'b00101001_11111010 : OUT <= 0;  //41 / 250 = 0
    16'b00101001_11111011 : OUT <= 0;  //41 / 251 = 0
    16'b00101001_11111100 : OUT <= 0;  //41 / 252 = 0
    16'b00101001_11111101 : OUT <= 0;  //41 / 253 = 0
    16'b00101001_11111110 : OUT <= 0;  //41 / 254 = 0
    16'b00101001_11111111 : OUT <= 0;  //41 / 255 = 0
    16'b00101010_00000000 : OUT <= 0;  //42 / 0 = 0
    16'b00101010_00000001 : OUT <= 42;  //42 / 1 = 42
    16'b00101010_00000010 : OUT <= 21;  //42 / 2 = 21
    16'b00101010_00000011 : OUT <= 14;  //42 / 3 = 14
    16'b00101010_00000100 : OUT <= 10;  //42 / 4 = 10
    16'b00101010_00000101 : OUT <= 8;  //42 / 5 = 8
    16'b00101010_00000110 : OUT <= 7;  //42 / 6 = 7
    16'b00101010_00000111 : OUT <= 6;  //42 / 7 = 6
    16'b00101010_00001000 : OUT <= 5;  //42 / 8 = 5
    16'b00101010_00001001 : OUT <= 4;  //42 / 9 = 4
    16'b00101010_00001010 : OUT <= 4;  //42 / 10 = 4
    16'b00101010_00001011 : OUT <= 3;  //42 / 11 = 3
    16'b00101010_00001100 : OUT <= 3;  //42 / 12 = 3
    16'b00101010_00001101 : OUT <= 3;  //42 / 13 = 3
    16'b00101010_00001110 : OUT <= 3;  //42 / 14 = 3
    16'b00101010_00001111 : OUT <= 2;  //42 / 15 = 2
    16'b00101010_00010000 : OUT <= 2;  //42 / 16 = 2
    16'b00101010_00010001 : OUT <= 2;  //42 / 17 = 2
    16'b00101010_00010010 : OUT <= 2;  //42 / 18 = 2
    16'b00101010_00010011 : OUT <= 2;  //42 / 19 = 2
    16'b00101010_00010100 : OUT <= 2;  //42 / 20 = 2
    16'b00101010_00010101 : OUT <= 2;  //42 / 21 = 2
    16'b00101010_00010110 : OUT <= 1;  //42 / 22 = 1
    16'b00101010_00010111 : OUT <= 1;  //42 / 23 = 1
    16'b00101010_00011000 : OUT <= 1;  //42 / 24 = 1
    16'b00101010_00011001 : OUT <= 1;  //42 / 25 = 1
    16'b00101010_00011010 : OUT <= 1;  //42 / 26 = 1
    16'b00101010_00011011 : OUT <= 1;  //42 / 27 = 1
    16'b00101010_00011100 : OUT <= 1;  //42 / 28 = 1
    16'b00101010_00011101 : OUT <= 1;  //42 / 29 = 1
    16'b00101010_00011110 : OUT <= 1;  //42 / 30 = 1
    16'b00101010_00011111 : OUT <= 1;  //42 / 31 = 1
    16'b00101010_00100000 : OUT <= 1;  //42 / 32 = 1
    16'b00101010_00100001 : OUT <= 1;  //42 / 33 = 1
    16'b00101010_00100010 : OUT <= 1;  //42 / 34 = 1
    16'b00101010_00100011 : OUT <= 1;  //42 / 35 = 1
    16'b00101010_00100100 : OUT <= 1;  //42 / 36 = 1
    16'b00101010_00100101 : OUT <= 1;  //42 / 37 = 1
    16'b00101010_00100110 : OUT <= 1;  //42 / 38 = 1
    16'b00101010_00100111 : OUT <= 1;  //42 / 39 = 1
    16'b00101010_00101000 : OUT <= 1;  //42 / 40 = 1
    16'b00101010_00101001 : OUT <= 1;  //42 / 41 = 1
    16'b00101010_00101010 : OUT <= 1;  //42 / 42 = 1
    16'b00101010_00101011 : OUT <= 0;  //42 / 43 = 0
    16'b00101010_00101100 : OUT <= 0;  //42 / 44 = 0
    16'b00101010_00101101 : OUT <= 0;  //42 / 45 = 0
    16'b00101010_00101110 : OUT <= 0;  //42 / 46 = 0
    16'b00101010_00101111 : OUT <= 0;  //42 / 47 = 0
    16'b00101010_00110000 : OUT <= 0;  //42 / 48 = 0
    16'b00101010_00110001 : OUT <= 0;  //42 / 49 = 0
    16'b00101010_00110010 : OUT <= 0;  //42 / 50 = 0
    16'b00101010_00110011 : OUT <= 0;  //42 / 51 = 0
    16'b00101010_00110100 : OUT <= 0;  //42 / 52 = 0
    16'b00101010_00110101 : OUT <= 0;  //42 / 53 = 0
    16'b00101010_00110110 : OUT <= 0;  //42 / 54 = 0
    16'b00101010_00110111 : OUT <= 0;  //42 / 55 = 0
    16'b00101010_00111000 : OUT <= 0;  //42 / 56 = 0
    16'b00101010_00111001 : OUT <= 0;  //42 / 57 = 0
    16'b00101010_00111010 : OUT <= 0;  //42 / 58 = 0
    16'b00101010_00111011 : OUT <= 0;  //42 / 59 = 0
    16'b00101010_00111100 : OUT <= 0;  //42 / 60 = 0
    16'b00101010_00111101 : OUT <= 0;  //42 / 61 = 0
    16'b00101010_00111110 : OUT <= 0;  //42 / 62 = 0
    16'b00101010_00111111 : OUT <= 0;  //42 / 63 = 0
    16'b00101010_01000000 : OUT <= 0;  //42 / 64 = 0
    16'b00101010_01000001 : OUT <= 0;  //42 / 65 = 0
    16'b00101010_01000010 : OUT <= 0;  //42 / 66 = 0
    16'b00101010_01000011 : OUT <= 0;  //42 / 67 = 0
    16'b00101010_01000100 : OUT <= 0;  //42 / 68 = 0
    16'b00101010_01000101 : OUT <= 0;  //42 / 69 = 0
    16'b00101010_01000110 : OUT <= 0;  //42 / 70 = 0
    16'b00101010_01000111 : OUT <= 0;  //42 / 71 = 0
    16'b00101010_01001000 : OUT <= 0;  //42 / 72 = 0
    16'b00101010_01001001 : OUT <= 0;  //42 / 73 = 0
    16'b00101010_01001010 : OUT <= 0;  //42 / 74 = 0
    16'b00101010_01001011 : OUT <= 0;  //42 / 75 = 0
    16'b00101010_01001100 : OUT <= 0;  //42 / 76 = 0
    16'b00101010_01001101 : OUT <= 0;  //42 / 77 = 0
    16'b00101010_01001110 : OUT <= 0;  //42 / 78 = 0
    16'b00101010_01001111 : OUT <= 0;  //42 / 79 = 0
    16'b00101010_01010000 : OUT <= 0;  //42 / 80 = 0
    16'b00101010_01010001 : OUT <= 0;  //42 / 81 = 0
    16'b00101010_01010010 : OUT <= 0;  //42 / 82 = 0
    16'b00101010_01010011 : OUT <= 0;  //42 / 83 = 0
    16'b00101010_01010100 : OUT <= 0;  //42 / 84 = 0
    16'b00101010_01010101 : OUT <= 0;  //42 / 85 = 0
    16'b00101010_01010110 : OUT <= 0;  //42 / 86 = 0
    16'b00101010_01010111 : OUT <= 0;  //42 / 87 = 0
    16'b00101010_01011000 : OUT <= 0;  //42 / 88 = 0
    16'b00101010_01011001 : OUT <= 0;  //42 / 89 = 0
    16'b00101010_01011010 : OUT <= 0;  //42 / 90 = 0
    16'b00101010_01011011 : OUT <= 0;  //42 / 91 = 0
    16'b00101010_01011100 : OUT <= 0;  //42 / 92 = 0
    16'b00101010_01011101 : OUT <= 0;  //42 / 93 = 0
    16'b00101010_01011110 : OUT <= 0;  //42 / 94 = 0
    16'b00101010_01011111 : OUT <= 0;  //42 / 95 = 0
    16'b00101010_01100000 : OUT <= 0;  //42 / 96 = 0
    16'b00101010_01100001 : OUT <= 0;  //42 / 97 = 0
    16'b00101010_01100010 : OUT <= 0;  //42 / 98 = 0
    16'b00101010_01100011 : OUT <= 0;  //42 / 99 = 0
    16'b00101010_01100100 : OUT <= 0;  //42 / 100 = 0
    16'b00101010_01100101 : OUT <= 0;  //42 / 101 = 0
    16'b00101010_01100110 : OUT <= 0;  //42 / 102 = 0
    16'b00101010_01100111 : OUT <= 0;  //42 / 103 = 0
    16'b00101010_01101000 : OUT <= 0;  //42 / 104 = 0
    16'b00101010_01101001 : OUT <= 0;  //42 / 105 = 0
    16'b00101010_01101010 : OUT <= 0;  //42 / 106 = 0
    16'b00101010_01101011 : OUT <= 0;  //42 / 107 = 0
    16'b00101010_01101100 : OUT <= 0;  //42 / 108 = 0
    16'b00101010_01101101 : OUT <= 0;  //42 / 109 = 0
    16'b00101010_01101110 : OUT <= 0;  //42 / 110 = 0
    16'b00101010_01101111 : OUT <= 0;  //42 / 111 = 0
    16'b00101010_01110000 : OUT <= 0;  //42 / 112 = 0
    16'b00101010_01110001 : OUT <= 0;  //42 / 113 = 0
    16'b00101010_01110010 : OUT <= 0;  //42 / 114 = 0
    16'b00101010_01110011 : OUT <= 0;  //42 / 115 = 0
    16'b00101010_01110100 : OUT <= 0;  //42 / 116 = 0
    16'b00101010_01110101 : OUT <= 0;  //42 / 117 = 0
    16'b00101010_01110110 : OUT <= 0;  //42 / 118 = 0
    16'b00101010_01110111 : OUT <= 0;  //42 / 119 = 0
    16'b00101010_01111000 : OUT <= 0;  //42 / 120 = 0
    16'b00101010_01111001 : OUT <= 0;  //42 / 121 = 0
    16'b00101010_01111010 : OUT <= 0;  //42 / 122 = 0
    16'b00101010_01111011 : OUT <= 0;  //42 / 123 = 0
    16'b00101010_01111100 : OUT <= 0;  //42 / 124 = 0
    16'b00101010_01111101 : OUT <= 0;  //42 / 125 = 0
    16'b00101010_01111110 : OUT <= 0;  //42 / 126 = 0
    16'b00101010_01111111 : OUT <= 0;  //42 / 127 = 0
    16'b00101010_10000000 : OUT <= 0;  //42 / 128 = 0
    16'b00101010_10000001 : OUT <= 0;  //42 / 129 = 0
    16'b00101010_10000010 : OUT <= 0;  //42 / 130 = 0
    16'b00101010_10000011 : OUT <= 0;  //42 / 131 = 0
    16'b00101010_10000100 : OUT <= 0;  //42 / 132 = 0
    16'b00101010_10000101 : OUT <= 0;  //42 / 133 = 0
    16'b00101010_10000110 : OUT <= 0;  //42 / 134 = 0
    16'b00101010_10000111 : OUT <= 0;  //42 / 135 = 0
    16'b00101010_10001000 : OUT <= 0;  //42 / 136 = 0
    16'b00101010_10001001 : OUT <= 0;  //42 / 137 = 0
    16'b00101010_10001010 : OUT <= 0;  //42 / 138 = 0
    16'b00101010_10001011 : OUT <= 0;  //42 / 139 = 0
    16'b00101010_10001100 : OUT <= 0;  //42 / 140 = 0
    16'b00101010_10001101 : OUT <= 0;  //42 / 141 = 0
    16'b00101010_10001110 : OUT <= 0;  //42 / 142 = 0
    16'b00101010_10001111 : OUT <= 0;  //42 / 143 = 0
    16'b00101010_10010000 : OUT <= 0;  //42 / 144 = 0
    16'b00101010_10010001 : OUT <= 0;  //42 / 145 = 0
    16'b00101010_10010010 : OUT <= 0;  //42 / 146 = 0
    16'b00101010_10010011 : OUT <= 0;  //42 / 147 = 0
    16'b00101010_10010100 : OUT <= 0;  //42 / 148 = 0
    16'b00101010_10010101 : OUT <= 0;  //42 / 149 = 0
    16'b00101010_10010110 : OUT <= 0;  //42 / 150 = 0
    16'b00101010_10010111 : OUT <= 0;  //42 / 151 = 0
    16'b00101010_10011000 : OUT <= 0;  //42 / 152 = 0
    16'b00101010_10011001 : OUT <= 0;  //42 / 153 = 0
    16'b00101010_10011010 : OUT <= 0;  //42 / 154 = 0
    16'b00101010_10011011 : OUT <= 0;  //42 / 155 = 0
    16'b00101010_10011100 : OUT <= 0;  //42 / 156 = 0
    16'b00101010_10011101 : OUT <= 0;  //42 / 157 = 0
    16'b00101010_10011110 : OUT <= 0;  //42 / 158 = 0
    16'b00101010_10011111 : OUT <= 0;  //42 / 159 = 0
    16'b00101010_10100000 : OUT <= 0;  //42 / 160 = 0
    16'b00101010_10100001 : OUT <= 0;  //42 / 161 = 0
    16'b00101010_10100010 : OUT <= 0;  //42 / 162 = 0
    16'b00101010_10100011 : OUT <= 0;  //42 / 163 = 0
    16'b00101010_10100100 : OUT <= 0;  //42 / 164 = 0
    16'b00101010_10100101 : OUT <= 0;  //42 / 165 = 0
    16'b00101010_10100110 : OUT <= 0;  //42 / 166 = 0
    16'b00101010_10100111 : OUT <= 0;  //42 / 167 = 0
    16'b00101010_10101000 : OUT <= 0;  //42 / 168 = 0
    16'b00101010_10101001 : OUT <= 0;  //42 / 169 = 0
    16'b00101010_10101010 : OUT <= 0;  //42 / 170 = 0
    16'b00101010_10101011 : OUT <= 0;  //42 / 171 = 0
    16'b00101010_10101100 : OUT <= 0;  //42 / 172 = 0
    16'b00101010_10101101 : OUT <= 0;  //42 / 173 = 0
    16'b00101010_10101110 : OUT <= 0;  //42 / 174 = 0
    16'b00101010_10101111 : OUT <= 0;  //42 / 175 = 0
    16'b00101010_10110000 : OUT <= 0;  //42 / 176 = 0
    16'b00101010_10110001 : OUT <= 0;  //42 / 177 = 0
    16'b00101010_10110010 : OUT <= 0;  //42 / 178 = 0
    16'b00101010_10110011 : OUT <= 0;  //42 / 179 = 0
    16'b00101010_10110100 : OUT <= 0;  //42 / 180 = 0
    16'b00101010_10110101 : OUT <= 0;  //42 / 181 = 0
    16'b00101010_10110110 : OUT <= 0;  //42 / 182 = 0
    16'b00101010_10110111 : OUT <= 0;  //42 / 183 = 0
    16'b00101010_10111000 : OUT <= 0;  //42 / 184 = 0
    16'b00101010_10111001 : OUT <= 0;  //42 / 185 = 0
    16'b00101010_10111010 : OUT <= 0;  //42 / 186 = 0
    16'b00101010_10111011 : OUT <= 0;  //42 / 187 = 0
    16'b00101010_10111100 : OUT <= 0;  //42 / 188 = 0
    16'b00101010_10111101 : OUT <= 0;  //42 / 189 = 0
    16'b00101010_10111110 : OUT <= 0;  //42 / 190 = 0
    16'b00101010_10111111 : OUT <= 0;  //42 / 191 = 0
    16'b00101010_11000000 : OUT <= 0;  //42 / 192 = 0
    16'b00101010_11000001 : OUT <= 0;  //42 / 193 = 0
    16'b00101010_11000010 : OUT <= 0;  //42 / 194 = 0
    16'b00101010_11000011 : OUT <= 0;  //42 / 195 = 0
    16'b00101010_11000100 : OUT <= 0;  //42 / 196 = 0
    16'b00101010_11000101 : OUT <= 0;  //42 / 197 = 0
    16'b00101010_11000110 : OUT <= 0;  //42 / 198 = 0
    16'b00101010_11000111 : OUT <= 0;  //42 / 199 = 0
    16'b00101010_11001000 : OUT <= 0;  //42 / 200 = 0
    16'b00101010_11001001 : OUT <= 0;  //42 / 201 = 0
    16'b00101010_11001010 : OUT <= 0;  //42 / 202 = 0
    16'b00101010_11001011 : OUT <= 0;  //42 / 203 = 0
    16'b00101010_11001100 : OUT <= 0;  //42 / 204 = 0
    16'b00101010_11001101 : OUT <= 0;  //42 / 205 = 0
    16'b00101010_11001110 : OUT <= 0;  //42 / 206 = 0
    16'b00101010_11001111 : OUT <= 0;  //42 / 207 = 0
    16'b00101010_11010000 : OUT <= 0;  //42 / 208 = 0
    16'b00101010_11010001 : OUT <= 0;  //42 / 209 = 0
    16'b00101010_11010010 : OUT <= 0;  //42 / 210 = 0
    16'b00101010_11010011 : OUT <= 0;  //42 / 211 = 0
    16'b00101010_11010100 : OUT <= 0;  //42 / 212 = 0
    16'b00101010_11010101 : OUT <= 0;  //42 / 213 = 0
    16'b00101010_11010110 : OUT <= 0;  //42 / 214 = 0
    16'b00101010_11010111 : OUT <= 0;  //42 / 215 = 0
    16'b00101010_11011000 : OUT <= 0;  //42 / 216 = 0
    16'b00101010_11011001 : OUT <= 0;  //42 / 217 = 0
    16'b00101010_11011010 : OUT <= 0;  //42 / 218 = 0
    16'b00101010_11011011 : OUT <= 0;  //42 / 219 = 0
    16'b00101010_11011100 : OUT <= 0;  //42 / 220 = 0
    16'b00101010_11011101 : OUT <= 0;  //42 / 221 = 0
    16'b00101010_11011110 : OUT <= 0;  //42 / 222 = 0
    16'b00101010_11011111 : OUT <= 0;  //42 / 223 = 0
    16'b00101010_11100000 : OUT <= 0;  //42 / 224 = 0
    16'b00101010_11100001 : OUT <= 0;  //42 / 225 = 0
    16'b00101010_11100010 : OUT <= 0;  //42 / 226 = 0
    16'b00101010_11100011 : OUT <= 0;  //42 / 227 = 0
    16'b00101010_11100100 : OUT <= 0;  //42 / 228 = 0
    16'b00101010_11100101 : OUT <= 0;  //42 / 229 = 0
    16'b00101010_11100110 : OUT <= 0;  //42 / 230 = 0
    16'b00101010_11100111 : OUT <= 0;  //42 / 231 = 0
    16'b00101010_11101000 : OUT <= 0;  //42 / 232 = 0
    16'b00101010_11101001 : OUT <= 0;  //42 / 233 = 0
    16'b00101010_11101010 : OUT <= 0;  //42 / 234 = 0
    16'b00101010_11101011 : OUT <= 0;  //42 / 235 = 0
    16'b00101010_11101100 : OUT <= 0;  //42 / 236 = 0
    16'b00101010_11101101 : OUT <= 0;  //42 / 237 = 0
    16'b00101010_11101110 : OUT <= 0;  //42 / 238 = 0
    16'b00101010_11101111 : OUT <= 0;  //42 / 239 = 0
    16'b00101010_11110000 : OUT <= 0;  //42 / 240 = 0
    16'b00101010_11110001 : OUT <= 0;  //42 / 241 = 0
    16'b00101010_11110010 : OUT <= 0;  //42 / 242 = 0
    16'b00101010_11110011 : OUT <= 0;  //42 / 243 = 0
    16'b00101010_11110100 : OUT <= 0;  //42 / 244 = 0
    16'b00101010_11110101 : OUT <= 0;  //42 / 245 = 0
    16'b00101010_11110110 : OUT <= 0;  //42 / 246 = 0
    16'b00101010_11110111 : OUT <= 0;  //42 / 247 = 0
    16'b00101010_11111000 : OUT <= 0;  //42 / 248 = 0
    16'b00101010_11111001 : OUT <= 0;  //42 / 249 = 0
    16'b00101010_11111010 : OUT <= 0;  //42 / 250 = 0
    16'b00101010_11111011 : OUT <= 0;  //42 / 251 = 0
    16'b00101010_11111100 : OUT <= 0;  //42 / 252 = 0
    16'b00101010_11111101 : OUT <= 0;  //42 / 253 = 0
    16'b00101010_11111110 : OUT <= 0;  //42 / 254 = 0
    16'b00101010_11111111 : OUT <= 0;  //42 / 255 = 0
    16'b00101011_00000000 : OUT <= 0;  //43 / 0 = 0
    16'b00101011_00000001 : OUT <= 43;  //43 / 1 = 43
    16'b00101011_00000010 : OUT <= 21;  //43 / 2 = 21
    16'b00101011_00000011 : OUT <= 14;  //43 / 3 = 14
    16'b00101011_00000100 : OUT <= 10;  //43 / 4 = 10
    16'b00101011_00000101 : OUT <= 8;  //43 / 5 = 8
    16'b00101011_00000110 : OUT <= 7;  //43 / 6 = 7
    16'b00101011_00000111 : OUT <= 6;  //43 / 7 = 6
    16'b00101011_00001000 : OUT <= 5;  //43 / 8 = 5
    16'b00101011_00001001 : OUT <= 4;  //43 / 9 = 4
    16'b00101011_00001010 : OUT <= 4;  //43 / 10 = 4
    16'b00101011_00001011 : OUT <= 3;  //43 / 11 = 3
    16'b00101011_00001100 : OUT <= 3;  //43 / 12 = 3
    16'b00101011_00001101 : OUT <= 3;  //43 / 13 = 3
    16'b00101011_00001110 : OUT <= 3;  //43 / 14 = 3
    16'b00101011_00001111 : OUT <= 2;  //43 / 15 = 2
    16'b00101011_00010000 : OUT <= 2;  //43 / 16 = 2
    16'b00101011_00010001 : OUT <= 2;  //43 / 17 = 2
    16'b00101011_00010010 : OUT <= 2;  //43 / 18 = 2
    16'b00101011_00010011 : OUT <= 2;  //43 / 19 = 2
    16'b00101011_00010100 : OUT <= 2;  //43 / 20 = 2
    16'b00101011_00010101 : OUT <= 2;  //43 / 21 = 2
    16'b00101011_00010110 : OUT <= 1;  //43 / 22 = 1
    16'b00101011_00010111 : OUT <= 1;  //43 / 23 = 1
    16'b00101011_00011000 : OUT <= 1;  //43 / 24 = 1
    16'b00101011_00011001 : OUT <= 1;  //43 / 25 = 1
    16'b00101011_00011010 : OUT <= 1;  //43 / 26 = 1
    16'b00101011_00011011 : OUT <= 1;  //43 / 27 = 1
    16'b00101011_00011100 : OUT <= 1;  //43 / 28 = 1
    16'b00101011_00011101 : OUT <= 1;  //43 / 29 = 1
    16'b00101011_00011110 : OUT <= 1;  //43 / 30 = 1
    16'b00101011_00011111 : OUT <= 1;  //43 / 31 = 1
    16'b00101011_00100000 : OUT <= 1;  //43 / 32 = 1
    16'b00101011_00100001 : OUT <= 1;  //43 / 33 = 1
    16'b00101011_00100010 : OUT <= 1;  //43 / 34 = 1
    16'b00101011_00100011 : OUT <= 1;  //43 / 35 = 1
    16'b00101011_00100100 : OUT <= 1;  //43 / 36 = 1
    16'b00101011_00100101 : OUT <= 1;  //43 / 37 = 1
    16'b00101011_00100110 : OUT <= 1;  //43 / 38 = 1
    16'b00101011_00100111 : OUT <= 1;  //43 / 39 = 1
    16'b00101011_00101000 : OUT <= 1;  //43 / 40 = 1
    16'b00101011_00101001 : OUT <= 1;  //43 / 41 = 1
    16'b00101011_00101010 : OUT <= 1;  //43 / 42 = 1
    16'b00101011_00101011 : OUT <= 1;  //43 / 43 = 1
    16'b00101011_00101100 : OUT <= 0;  //43 / 44 = 0
    16'b00101011_00101101 : OUT <= 0;  //43 / 45 = 0
    16'b00101011_00101110 : OUT <= 0;  //43 / 46 = 0
    16'b00101011_00101111 : OUT <= 0;  //43 / 47 = 0
    16'b00101011_00110000 : OUT <= 0;  //43 / 48 = 0
    16'b00101011_00110001 : OUT <= 0;  //43 / 49 = 0
    16'b00101011_00110010 : OUT <= 0;  //43 / 50 = 0
    16'b00101011_00110011 : OUT <= 0;  //43 / 51 = 0
    16'b00101011_00110100 : OUT <= 0;  //43 / 52 = 0
    16'b00101011_00110101 : OUT <= 0;  //43 / 53 = 0
    16'b00101011_00110110 : OUT <= 0;  //43 / 54 = 0
    16'b00101011_00110111 : OUT <= 0;  //43 / 55 = 0
    16'b00101011_00111000 : OUT <= 0;  //43 / 56 = 0
    16'b00101011_00111001 : OUT <= 0;  //43 / 57 = 0
    16'b00101011_00111010 : OUT <= 0;  //43 / 58 = 0
    16'b00101011_00111011 : OUT <= 0;  //43 / 59 = 0
    16'b00101011_00111100 : OUT <= 0;  //43 / 60 = 0
    16'b00101011_00111101 : OUT <= 0;  //43 / 61 = 0
    16'b00101011_00111110 : OUT <= 0;  //43 / 62 = 0
    16'b00101011_00111111 : OUT <= 0;  //43 / 63 = 0
    16'b00101011_01000000 : OUT <= 0;  //43 / 64 = 0
    16'b00101011_01000001 : OUT <= 0;  //43 / 65 = 0
    16'b00101011_01000010 : OUT <= 0;  //43 / 66 = 0
    16'b00101011_01000011 : OUT <= 0;  //43 / 67 = 0
    16'b00101011_01000100 : OUT <= 0;  //43 / 68 = 0
    16'b00101011_01000101 : OUT <= 0;  //43 / 69 = 0
    16'b00101011_01000110 : OUT <= 0;  //43 / 70 = 0
    16'b00101011_01000111 : OUT <= 0;  //43 / 71 = 0
    16'b00101011_01001000 : OUT <= 0;  //43 / 72 = 0
    16'b00101011_01001001 : OUT <= 0;  //43 / 73 = 0
    16'b00101011_01001010 : OUT <= 0;  //43 / 74 = 0
    16'b00101011_01001011 : OUT <= 0;  //43 / 75 = 0
    16'b00101011_01001100 : OUT <= 0;  //43 / 76 = 0
    16'b00101011_01001101 : OUT <= 0;  //43 / 77 = 0
    16'b00101011_01001110 : OUT <= 0;  //43 / 78 = 0
    16'b00101011_01001111 : OUT <= 0;  //43 / 79 = 0
    16'b00101011_01010000 : OUT <= 0;  //43 / 80 = 0
    16'b00101011_01010001 : OUT <= 0;  //43 / 81 = 0
    16'b00101011_01010010 : OUT <= 0;  //43 / 82 = 0
    16'b00101011_01010011 : OUT <= 0;  //43 / 83 = 0
    16'b00101011_01010100 : OUT <= 0;  //43 / 84 = 0
    16'b00101011_01010101 : OUT <= 0;  //43 / 85 = 0
    16'b00101011_01010110 : OUT <= 0;  //43 / 86 = 0
    16'b00101011_01010111 : OUT <= 0;  //43 / 87 = 0
    16'b00101011_01011000 : OUT <= 0;  //43 / 88 = 0
    16'b00101011_01011001 : OUT <= 0;  //43 / 89 = 0
    16'b00101011_01011010 : OUT <= 0;  //43 / 90 = 0
    16'b00101011_01011011 : OUT <= 0;  //43 / 91 = 0
    16'b00101011_01011100 : OUT <= 0;  //43 / 92 = 0
    16'b00101011_01011101 : OUT <= 0;  //43 / 93 = 0
    16'b00101011_01011110 : OUT <= 0;  //43 / 94 = 0
    16'b00101011_01011111 : OUT <= 0;  //43 / 95 = 0
    16'b00101011_01100000 : OUT <= 0;  //43 / 96 = 0
    16'b00101011_01100001 : OUT <= 0;  //43 / 97 = 0
    16'b00101011_01100010 : OUT <= 0;  //43 / 98 = 0
    16'b00101011_01100011 : OUT <= 0;  //43 / 99 = 0
    16'b00101011_01100100 : OUT <= 0;  //43 / 100 = 0
    16'b00101011_01100101 : OUT <= 0;  //43 / 101 = 0
    16'b00101011_01100110 : OUT <= 0;  //43 / 102 = 0
    16'b00101011_01100111 : OUT <= 0;  //43 / 103 = 0
    16'b00101011_01101000 : OUT <= 0;  //43 / 104 = 0
    16'b00101011_01101001 : OUT <= 0;  //43 / 105 = 0
    16'b00101011_01101010 : OUT <= 0;  //43 / 106 = 0
    16'b00101011_01101011 : OUT <= 0;  //43 / 107 = 0
    16'b00101011_01101100 : OUT <= 0;  //43 / 108 = 0
    16'b00101011_01101101 : OUT <= 0;  //43 / 109 = 0
    16'b00101011_01101110 : OUT <= 0;  //43 / 110 = 0
    16'b00101011_01101111 : OUT <= 0;  //43 / 111 = 0
    16'b00101011_01110000 : OUT <= 0;  //43 / 112 = 0
    16'b00101011_01110001 : OUT <= 0;  //43 / 113 = 0
    16'b00101011_01110010 : OUT <= 0;  //43 / 114 = 0
    16'b00101011_01110011 : OUT <= 0;  //43 / 115 = 0
    16'b00101011_01110100 : OUT <= 0;  //43 / 116 = 0
    16'b00101011_01110101 : OUT <= 0;  //43 / 117 = 0
    16'b00101011_01110110 : OUT <= 0;  //43 / 118 = 0
    16'b00101011_01110111 : OUT <= 0;  //43 / 119 = 0
    16'b00101011_01111000 : OUT <= 0;  //43 / 120 = 0
    16'b00101011_01111001 : OUT <= 0;  //43 / 121 = 0
    16'b00101011_01111010 : OUT <= 0;  //43 / 122 = 0
    16'b00101011_01111011 : OUT <= 0;  //43 / 123 = 0
    16'b00101011_01111100 : OUT <= 0;  //43 / 124 = 0
    16'b00101011_01111101 : OUT <= 0;  //43 / 125 = 0
    16'b00101011_01111110 : OUT <= 0;  //43 / 126 = 0
    16'b00101011_01111111 : OUT <= 0;  //43 / 127 = 0
    16'b00101011_10000000 : OUT <= 0;  //43 / 128 = 0
    16'b00101011_10000001 : OUT <= 0;  //43 / 129 = 0
    16'b00101011_10000010 : OUT <= 0;  //43 / 130 = 0
    16'b00101011_10000011 : OUT <= 0;  //43 / 131 = 0
    16'b00101011_10000100 : OUT <= 0;  //43 / 132 = 0
    16'b00101011_10000101 : OUT <= 0;  //43 / 133 = 0
    16'b00101011_10000110 : OUT <= 0;  //43 / 134 = 0
    16'b00101011_10000111 : OUT <= 0;  //43 / 135 = 0
    16'b00101011_10001000 : OUT <= 0;  //43 / 136 = 0
    16'b00101011_10001001 : OUT <= 0;  //43 / 137 = 0
    16'b00101011_10001010 : OUT <= 0;  //43 / 138 = 0
    16'b00101011_10001011 : OUT <= 0;  //43 / 139 = 0
    16'b00101011_10001100 : OUT <= 0;  //43 / 140 = 0
    16'b00101011_10001101 : OUT <= 0;  //43 / 141 = 0
    16'b00101011_10001110 : OUT <= 0;  //43 / 142 = 0
    16'b00101011_10001111 : OUT <= 0;  //43 / 143 = 0
    16'b00101011_10010000 : OUT <= 0;  //43 / 144 = 0
    16'b00101011_10010001 : OUT <= 0;  //43 / 145 = 0
    16'b00101011_10010010 : OUT <= 0;  //43 / 146 = 0
    16'b00101011_10010011 : OUT <= 0;  //43 / 147 = 0
    16'b00101011_10010100 : OUT <= 0;  //43 / 148 = 0
    16'b00101011_10010101 : OUT <= 0;  //43 / 149 = 0
    16'b00101011_10010110 : OUT <= 0;  //43 / 150 = 0
    16'b00101011_10010111 : OUT <= 0;  //43 / 151 = 0
    16'b00101011_10011000 : OUT <= 0;  //43 / 152 = 0
    16'b00101011_10011001 : OUT <= 0;  //43 / 153 = 0
    16'b00101011_10011010 : OUT <= 0;  //43 / 154 = 0
    16'b00101011_10011011 : OUT <= 0;  //43 / 155 = 0
    16'b00101011_10011100 : OUT <= 0;  //43 / 156 = 0
    16'b00101011_10011101 : OUT <= 0;  //43 / 157 = 0
    16'b00101011_10011110 : OUT <= 0;  //43 / 158 = 0
    16'b00101011_10011111 : OUT <= 0;  //43 / 159 = 0
    16'b00101011_10100000 : OUT <= 0;  //43 / 160 = 0
    16'b00101011_10100001 : OUT <= 0;  //43 / 161 = 0
    16'b00101011_10100010 : OUT <= 0;  //43 / 162 = 0
    16'b00101011_10100011 : OUT <= 0;  //43 / 163 = 0
    16'b00101011_10100100 : OUT <= 0;  //43 / 164 = 0
    16'b00101011_10100101 : OUT <= 0;  //43 / 165 = 0
    16'b00101011_10100110 : OUT <= 0;  //43 / 166 = 0
    16'b00101011_10100111 : OUT <= 0;  //43 / 167 = 0
    16'b00101011_10101000 : OUT <= 0;  //43 / 168 = 0
    16'b00101011_10101001 : OUT <= 0;  //43 / 169 = 0
    16'b00101011_10101010 : OUT <= 0;  //43 / 170 = 0
    16'b00101011_10101011 : OUT <= 0;  //43 / 171 = 0
    16'b00101011_10101100 : OUT <= 0;  //43 / 172 = 0
    16'b00101011_10101101 : OUT <= 0;  //43 / 173 = 0
    16'b00101011_10101110 : OUT <= 0;  //43 / 174 = 0
    16'b00101011_10101111 : OUT <= 0;  //43 / 175 = 0
    16'b00101011_10110000 : OUT <= 0;  //43 / 176 = 0
    16'b00101011_10110001 : OUT <= 0;  //43 / 177 = 0
    16'b00101011_10110010 : OUT <= 0;  //43 / 178 = 0
    16'b00101011_10110011 : OUT <= 0;  //43 / 179 = 0
    16'b00101011_10110100 : OUT <= 0;  //43 / 180 = 0
    16'b00101011_10110101 : OUT <= 0;  //43 / 181 = 0
    16'b00101011_10110110 : OUT <= 0;  //43 / 182 = 0
    16'b00101011_10110111 : OUT <= 0;  //43 / 183 = 0
    16'b00101011_10111000 : OUT <= 0;  //43 / 184 = 0
    16'b00101011_10111001 : OUT <= 0;  //43 / 185 = 0
    16'b00101011_10111010 : OUT <= 0;  //43 / 186 = 0
    16'b00101011_10111011 : OUT <= 0;  //43 / 187 = 0
    16'b00101011_10111100 : OUT <= 0;  //43 / 188 = 0
    16'b00101011_10111101 : OUT <= 0;  //43 / 189 = 0
    16'b00101011_10111110 : OUT <= 0;  //43 / 190 = 0
    16'b00101011_10111111 : OUT <= 0;  //43 / 191 = 0
    16'b00101011_11000000 : OUT <= 0;  //43 / 192 = 0
    16'b00101011_11000001 : OUT <= 0;  //43 / 193 = 0
    16'b00101011_11000010 : OUT <= 0;  //43 / 194 = 0
    16'b00101011_11000011 : OUT <= 0;  //43 / 195 = 0
    16'b00101011_11000100 : OUT <= 0;  //43 / 196 = 0
    16'b00101011_11000101 : OUT <= 0;  //43 / 197 = 0
    16'b00101011_11000110 : OUT <= 0;  //43 / 198 = 0
    16'b00101011_11000111 : OUT <= 0;  //43 / 199 = 0
    16'b00101011_11001000 : OUT <= 0;  //43 / 200 = 0
    16'b00101011_11001001 : OUT <= 0;  //43 / 201 = 0
    16'b00101011_11001010 : OUT <= 0;  //43 / 202 = 0
    16'b00101011_11001011 : OUT <= 0;  //43 / 203 = 0
    16'b00101011_11001100 : OUT <= 0;  //43 / 204 = 0
    16'b00101011_11001101 : OUT <= 0;  //43 / 205 = 0
    16'b00101011_11001110 : OUT <= 0;  //43 / 206 = 0
    16'b00101011_11001111 : OUT <= 0;  //43 / 207 = 0
    16'b00101011_11010000 : OUT <= 0;  //43 / 208 = 0
    16'b00101011_11010001 : OUT <= 0;  //43 / 209 = 0
    16'b00101011_11010010 : OUT <= 0;  //43 / 210 = 0
    16'b00101011_11010011 : OUT <= 0;  //43 / 211 = 0
    16'b00101011_11010100 : OUT <= 0;  //43 / 212 = 0
    16'b00101011_11010101 : OUT <= 0;  //43 / 213 = 0
    16'b00101011_11010110 : OUT <= 0;  //43 / 214 = 0
    16'b00101011_11010111 : OUT <= 0;  //43 / 215 = 0
    16'b00101011_11011000 : OUT <= 0;  //43 / 216 = 0
    16'b00101011_11011001 : OUT <= 0;  //43 / 217 = 0
    16'b00101011_11011010 : OUT <= 0;  //43 / 218 = 0
    16'b00101011_11011011 : OUT <= 0;  //43 / 219 = 0
    16'b00101011_11011100 : OUT <= 0;  //43 / 220 = 0
    16'b00101011_11011101 : OUT <= 0;  //43 / 221 = 0
    16'b00101011_11011110 : OUT <= 0;  //43 / 222 = 0
    16'b00101011_11011111 : OUT <= 0;  //43 / 223 = 0
    16'b00101011_11100000 : OUT <= 0;  //43 / 224 = 0
    16'b00101011_11100001 : OUT <= 0;  //43 / 225 = 0
    16'b00101011_11100010 : OUT <= 0;  //43 / 226 = 0
    16'b00101011_11100011 : OUT <= 0;  //43 / 227 = 0
    16'b00101011_11100100 : OUT <= 0;  //43 / 228 = 0
    16'b00101011_11100101 : OUT <= 0;  //43 / 229 = 0
    16'b00101011_11100110 : OUT <= 0;  //43 / 230 = 0
    16'b00101011_11100111 : OUT <= 0;  //43 / 231 = 0
    16'b00101011_11101000 : OUT <= 0;  //43 / 232 = 0
    16'b00101011_11101001 : OUT <= 0;  //43 / 233 = 0
    16'b00101011_11101010 : OUT <= 0;  //43 / 234 = 0
    16'b00101011_11101011 : OUT <= 0;  //43 / 235 = 0
    16'b00101011_11101100 : OUT <= 0;  //43 / 236 = 0
    16'b00101011_11101101 : OUT <= 0;  //43 / 237 = 0
    16'b00101011_11101110 : OUT <= 0;  //43 / 238 = 0
    16'b00101011_11101111 : OUT <= 0;  //43 / 239 = 0
    16'b00101011_11110000 : OUT <= 0;  //43 / 240 = 0
    16'b00101011_11110001 : OUT <= 0;  //43 / 241 = 0
    16'b00101011_11110010 : OUT <= 0;  //43 / 242 = 0
    16'b00101011_11110011 : OUT <= 0;  //43 / 243 = 0
    16'b00101011_11110100 : OUT <= 0;  //43 / 244 = 0
    16'b00101011_11110101 : OUT <= 0;  //43 / 245 = 0
    16'b00101011_11110110 : OUT <= 0;  //43 / 246 = 0
    16'b00101011_11110111 : OUT <= 0;  //43 / 247 = 0
    16'b00101011_11111000 : OUT <= 0;  //43 / 248 = 0
    16'b00101011_11111001 : OUT <= 0;  //43 / 249 = 0
    16'b00101011_11111010 : OUT <= 0;  //43 / 250 = 0
    16'b00101011_11111011 : OUT <= 0;  //43 / 251 = 0
    16'b00101011_11111100 : OUT <= 0;  //43 / 252 = 0
    16'b00101011_11111101 : OUT <= 0;  //43 / 253 = 0
    16'b00101011_11111110 : OUT <= 0;  //43 / 254 = 0
    16'b00101011_11111111 : OUT <= 0;  //43 / 255 = 0
    16'b00101100_00000000 : OUT <= 0;  //44 / 0 = 0
    16'b00101100_00000001 : OUT <= 44;  //44 / 1 = 44
    16'b00101100_00000010 : OUT <= 22;  //44 / 2 = 22
    16'b00101100_00000011 : OUT <= 14;  //44 / 3 = 14
    16'b00101100_00000100 : OUT <= 11;  //44 / 4 = 11
    16'b00101100_00000101 : OUT <= 8;  //44 / 5 = 8
    16'b00101100_00000110 : OUT <= 7;  //44 / 6 = 7
    16'b00101100_00000111 : OUT <= 6;  //44 / 7 = 6
    16'b00101100_00001000 : OUT <= 5;  //44 / 8 = 5
    16'b00101100_00001001 : OUT <= 4;  //44 / 9 = 4
    16'b00101100_00001010 : OUT <= 4;  //44 / 10 = 4
    16'b00101100_00001011 : OUT <= 4;  //44 / 11 = 4
    16'b00101100_00001100 : OUT <= 3;  //44 / 12 = 3
    16'b00101100_00001101 : OUT <= 3;  //44 / 13 = 3
    16'b00101100_00001110 : OUT <= 3;  //44 / 14 = 3
    16'b00101100_00001111 : OUT <= 2;  //44 / 15 = 2
    16'b00101100_00010000 : OUT <= 2;  //44 / 16 = 2
    16'b00101100_00010001 : OUT <= 2;  //44 / 17 = 2
    16'b00101100_00010010 : OUT <= 2;  //44 / 18 = 2
    16'b00101100_00010011 : OUT <= 2;  //44 / 19 = 2
    16'b00101100_00010100 : OUT <= 2;  //44 / 20 = 2
    16'b00101100_00010101 : OUT <= 2;  //44 / 21 = 2
    16'b00101100_00010110 : OUT <= 2;  //44 / 22 = 2
    16'b00101100_00010111 : OUT <= 1;  //44 / 23 = 1
    16'b00101100_00011000 : OUT <= 1;  //44 / 24 = 1
    16'b00101100_00011001 : OUT <= 1;  //44 / 25 = 1
    16'b00101100_00011010 : OUT <= 1;  //44 / 26 = 1
    16'b00101100_00011011 : OUT <= 1;  //44 / 27 = 1
    16'b00101100_00011100 : OUT <= 1;  //44 / 28 = 1
    16'b00101100_00011101 : OUT <= 1;  //44 / 29 = 1
    16'b00101100_00011110 : OUT <= 1;  //44 / 30 = 1
    16'b00101100_00011111 : OUT <= 1;  //44 / 31 = 1
    16'b00101100_00100000 : OUT <= 1;  //44 / 32 = 1
    16'b00101100_00100001 : OUT <= 1;  //44 / 33 = 1
    16'b00101100_00100010 : OUT <= 1;  //44 / 34 = 1
    16'b00101100_00100011 : OUT <= 1;  //44 / 35 = 1
    16'b00101100_00100100 : OUT <= 1;  //44 / 36 = 1
    16'b00101100_00100101 : OUT <= 1;  //44 / 37 = 1
    16'b00101100_00100110 : OUT <= 1;  //44 / 38 = 1
    16'b00101100_00100111 : OUT <= 1;  //44 / 39 = 1
    16'b00101100_00101000 : OUT <= 1;  //44 / 40 = 1
    16'b00101100_00101001 : OUT <= 1;  //44 / 41 = 1
    16'b00101100_00101010 : OUT <= 1;  //44 / 42 = 1
    16'b00101100_00101011 : OUT <= 1;  //44 / 43 = 1
    16'b00101100_00101100 : OUT <= 1;  //44 / 44 = 1
    16'b00101100_00101101 : OUT <= 0;  //44 / 45 = 0
    16'b00101100_00101110 : OUT <= 0;  //44 / 46 = 0
    16'b00101100_00101111 : OUT <= 0;  //44 / 47 = 0
    16'b00101100_00110000 : OUT <= 0;  //44 / 48 = 0
    16'b00101100_00110001 : OUT <= 0;  //44 / 49 = 0
    16'b00101100_00110010 : OUT <= 0;  //44 / 50 = 0
    16'b00101100_00110011 : OUT <= 0;  //44 / 51 = 0
    16'b00101100_00110100 : OUT <= 0;  //44 / 52 = 0
    16'b00101100_00110101 : OUT <= 0;  //44 / 53 = 0
    16'b00101100_00110110 : OUT <= 0;  //44 / 54 = 0
    16'b00101100_00110111 : OUT <= 0;  //44 / 55 = 0
    16'b00101100_00111000 : OUT <= 0;  //44 / 56 = 0
    16'b00101100_00111001 : OUT <= 0;  //44 / 57 = 0
    16'b00101100_00111010 : OUT <= 0;  //44 / 58 = 0
    16'b00101100_00111011 : OUT <= 0;  //44 / 59 = 0
    16'b00101100_00111100 : OUT <= 0;  //44 / 60 = 0
    16'b00101100_00111101 : OUT <= 0;  //44 / 61 = 0
    16'b00101100_00111110 : OUT <= 0;  //44 / 62 = 0
    16'b00101100_00111111 : OUT <= 0;  //44 / 63 = 0
    16'b00101100_01000000 : OUT <= 0;  //44 / 64 = 0
    16'b00101100_01000001 : OUT <= 0;  //44 / 65 = 0
    16'b00101100_01000010 : OUT <= 0;  //44 / 66 = 0
    16'b00101100_01000011 : OUT <= 0;  //44 / 67 = 0
    16'b00101100_01000100 : OUT <= 0;  //44 / 68 = 0
    16'b00101100_01000101 : OUT <= 0;  //44 / 69 = 0
    16'b00101100_01000110 : OUT <= 0;  //44 / 70 = 0
    16'b00101100_01000111 : OUT <= 0;  //44 / 71 = 0
    16'b00101100_01001000 : OUT <= 0;  //44 / 72 = 0
    16'b00101100_01001001 : OUT <= 0;  //44 / 73 = 0
    16'b00101100_01001010 : OUT <= 0;  //44 / 74 = 0
    16'b00101100_01001011 : OUT <= 0;  //44 / 75 = 0
    16'b00101100_01001100 : OUT <= 0;  //44 / 76 = 0
    16'b00101100_01001101 : OUT <= 0;  //44 / 77 = 0
    16'b00101100_01001110 : OUT <= 0;  //44 / 78 = 0
    16'b00101100_01001111 : OUT <= 0;  //44 / 79 = 0
    16'b00101100_01010000 : OUT <= 0;  //44 / 80 = 0
    16'b00101100_01010001 : OUT <= 0;  //44 / 81 = 0
    16'b00101100_01010010 : OUT <= 0;  //44 / 82 = 0
    16'b00101100_01010011 : OUT <= 0;  //44 / 83 = 0
    16'b00101100_01010100 : OUT <= 0;  //44 / 84 = 0
    16'b00101100_01010101 : OUT <= 0;  //44 / 85 = 0
    16'b00101100_01010110 : OUT <= 0;  //44 / 86 = 0
    16'b00101100_01010111 : OUT <= 0;  //44 / 87 = 0
    16'b00101100_01011000 : OUT <= 0;  //44 / 88 = 0
    16'b00101100_01011001 : OUT <= 0;  //44 / 89 = 0
    16'b00101100_01011010 : OUT <= 0;  //44 / 90 = 0
    16'b00101100_01011011 : OUT <= 0;  //44 / 91 = 0
    16'b00101100_01011100 : OUT <= 0;  //44 / 92 = 0
    16'b00101100_01011101 : OUT <= 0;  //44 / 93 = 0
    16'b00101100_01011110 : OUT <= 0;  //44 / 94 = 0
    16'b00101100_01011111 : OUT <= 0;  //44 / 95 = 0
    16'b00101100_01100000 : OUT <= 0;  //44 / 96 = 0
    16'b00101100_01100001 : OUT <= 0;  //44 / 97 = 0
    16'b00101100_01100010 : OUT <= 0;  //44 / 98 = 0
    16'b00101100_01100011 : OUT <= 0;  //44 / 99 = 0
    16'b00101100_01100100 : OUT <= 0;  //44 / 100 = 0
    16'b00101100_01100101 : OUT <= 0;  //44 / 101 = 0
    16'b00101100_01100110 : OUT <= 0;  //44 / 102 = 0
    16'b00101100_01100111 : OUT <= 0;  //44 / 103 = 0
    16'b00101100_01101000 : OUT <= 0;  //44 / 104 = 0
    16'b00101100_01101001 : OUT <= 0;  //44 / 105 = 0
    16'b00101100_01101010 : OUT <= 0;  //44 / 106 = 0
    16'b00101100_01101011 : OUT <= 0;  //44 / 107 = 0
    16'b00101100_01101100 : OUT <= 0;  //44 / 108 = 0
    16'b00101100_01101101 : OUT <= 0;  //44 / 109 = 0
    16'b00101100_01101110 : OUT <= 0;  //44 / 110 = 0
    16'b00101100_01101111 : OUT <= 0;  //44 / 111 = 0
    16'b00101100_01110000 : OUT <= 0;  //44 / 112 = 0
    16'b00101100_01110001 : OUT <= 0;  //44 / 113 = 0
    16'b00101100_01110010 : OUT <= 0;  //44 / 114 = 0
    16'b00101100_01110011 : OUT <= 0;  //44 / 115 = 0
    16'b00101100_01110100 : OUT <= 0;  //44 / 116 = 0
    16'b00101100_01110101 : OUT <= 0;  //44 / 117 = 0
    16'b00101100_01110110 : OUT <= 0;  //44 / 118 = 0
    16'b00101100_01110111 : OUT <= 0;  //44 / 119 = 0
    16'b00101100_01111000 : OUT <= 0;  //44 / 120 = 0
    16'b00101100_01111001 : OUT <= 0;  //44 / 121 = 0
    16'b00101100_01111010 : OUT <= 0;  //44 / 122 = 0
    16'b00101100_01111011 : OUT <= 0;  //44 / 123 = 0
    16'b00101100_01111100 : OUT <= 0;  //44 / 124 = 0
    16'b00101100_01111101 : OUT <= 0;  //44 / 125 = 0
    16'b00101100_01111110 : OUT <= 0;  //44 / 126 = 0
    16'b00101100_01111111 : OUT <= 0;  //44 / 127 = 0
    16'b00101100_10000000 : OUT <= 0;  //44 / 128 = 0
    16'b00101100_10000001 : OUT <= 0;  //44 / 129 = 0
    16'b00101100_10000010 : OUT <= 0;  //44 / 130 = 0
    16'b00101100_10000011 : OUT <= 0;  //44 / 131 = 0
    16'b00101100_10000100 : OUT <= 0;  //44 / 132 = 0
    16'b00101100_10000101 : OUT <= 0;  //44 / 133 = 0
    16'b00101100_10000110 : OUT <= 0;  //44 / 134 = 0
    16'b00101100_10000111 : OUT <= 0;  //44 / 135 = 0
    16'b00101100_10001000 : OUT <= 0;  //44 / 136 = 0
    16'b00101100_10001001 : OUT <= 0;  //44 / 137 = 0
    16'b00101100_10001010 : OUT <= 0;  //44 / 138 = 0
    16'b00101100_10001011 : OUT <= 0;  //44 / 139 = 0
    16'b00101100_10001100 : OUT <= 0;  //44 / 140 = 0
    16'b00101100_10001101 : OUT <= 0;  //44 / 141 = 0
    16'b00101100_10001110 : OUT <= 0;  //44 / 142 = 0
    16'b00101100_10001111 : OUT <= 0;  //44 / 143 = 0
    16'b00101100_10010000 : OUT <= 0;  //44 / 144 = 0
    16'b00101100_10010001 : OUT <= 0;  //44 / 145 = 0
    16'b00101100_10010010 : OUT <= 0;  //44 / 146 = 0
    16'b00101100_10010011 : OUT <= 0;  //44 / 147 = 0
    16'b00101100_10010100 : OUT <= 0;  //44 / 148 = 0
    16'b00101100_10010101 : OUT <= 0;  //44 / 149 = 0
    16'b00101100_10010110 : OUT <= 0;  //44 / 150 = 0
    16'b00101100_10010111 : OUT <= 0;  //44 / 151 = 0
    16'b00101100_10011000 : OUT <= 0;  //44 / 152 = 0
    16'b00101100_10011001 : OUT <= 0;  //44 / 153 = 0
    16'b00101100_10011010 : OUT <= 0;  //44 / 154 = 0
    16'b00101100_10011011 : OUT <= 0;  //44 / 155 = 0
    16'b00101100_10011100 : OUT <= 0;  //44 / 156 = 0
    16'b00101100_10011101 : OUT <= 0;  //44 / 157 = 0
    16'b00101100_10011110 : OUT <= 0;  //44 / 158 = 0
    16'b00101100_10011111 : OUT <= 0;  //44 / 159 = 0
    16'b00101100_10100000 : OUT <= 0;  //44 / 160 = 0
    16'b00101100_10100001 : OUT <= 0;  //44 / 161 = 0
    16'b00101100_10100010 : OUT <= 0;  //44 / 162 = 0
    16'b00101100_10100011 : OUT <= 0;  //44 / 163 = 0
    16'b00101100_10100100 : OUT <= 0;  //44 / 164 = 0
    16'b00101100_10100101 : OUT <= 0;  //44 / 165 = 0
    16'b00101100_10100110 : OUT <= 0;  //44 / 166 = 0
    16'b00101100_10100111 : OUT <= 0;  //44 / 167 = 0
    16'b00101100_10101000 : OUT <= 0;  //44 / 168 = 0
    16'b00101100_10101001 : OUT <= 0;  //44 / 169 = 0
    16'b00101100_10101010 : OUT <= 0;  //44 / 170 = 0
    16'b00101100_10101011 : OUT <= 0;  //44 / 171 = 0
    16'b00101100_10101100 : OUT <= 0;  //44 / 172 = 0
    16'b00101100_10101101 : OUT <= 0;  //44 / 173 = 0
    16'b00101100_10101110 : OUT <= 0;  //44 / 174 = 0
    16'b00101100_10101111 : OUT <= 0;  //44 / 175 = 0
    16'b00101100_10110000 : OUT <= 0;  //44 / 176 = 0
    16'b00101100_10110001 : OUT <= 0;  //44 / 177 = 0
    16'b00101100_10110010 : OUT <= 0;  //44 / 178 = 0
    16'b00101100_10110011 : OUT <= 0;  //44 / 179 = 0
    16'b00101100_10110100 : OUT <= 0;  //44 / 180 = 0
    16'b00101100_10110101 : OUT <= 0;  //44 / 181 = 0
    16'b00101100_10110110 : OUT <= 0;  //44 / 182 = 0
    16'b00101100_10110111 : OUT <= 0;  //44 / 183 = 0
    16'b00101100_10111000 : OUT <= 0;  //44 / 184 = 0
    16'b00101100_10111001 : OUT <= 0;  //44 / 185 = 0
    16'b00101100_10111010 : OUT <= 0;  //44 / 186 = 0
    16'b00101100_10111011 : OUT <= 0;  //44 / 187 = 0
    16'b00101100_10111100 : OUT <= 0;  //44 / 188 = 0
    16'b00101100_10111101 : OUT <= 0;  //44 / 189 = 0
    16'b00101100_10111110 : OUT <= 0;  //44 / 190 = 0
    16'b00101100_10111111 : OUT <= 0;  //44 / 191 = 0
    16'b00101100_11000000 : OUT <= 0;  //44 / 192 = 0
    16'b00101100_11000001 : OUT <= 0;  //44 / 193 = 0
    16'b00101100_11000010 : OUT <= 0;  //44 / 194 = 0
    16'b00101100_11000011 : OUT <= 0;  //44 / 195 = 0
    16'b00101100_11000100 : OUT <= 0;  //44 / 196 = 0
    16'b00101100_11000101 : OUT <= 0;  //44 / 197 = 0
    16'b00101100_11000110 : OUT <= 0;  //44 / 198 = 0
    16'b00101100_11000111 : OUT <= 0;  //44 / 199 = 0
    16'b00101100_11001000 : OUT <= 0;  //44 / 200 = 0
    16'b00101100_11001001 : OUT <= 0;  //44 / 201 = 0
    16'b00101100_11001010 : OUT <= 0;  //44 / 202 = 0
    16'b00101100_11001011 : OUT <= 0;  //44 / 203 = 0
    16'b00101100_11001100 : OUT <= 0;  //44 / 204 = 0
    16'b00101100_11001101 : OUT <= 0;  //44 / 205 = 0
    16'b00101100_11001110 : OUT <= 0;  //44 / 206 = 0
    16'b00101100_11001111 : OUT <= 0;  //44 / 207 = 0
    16'b00101100_11010000 : OUT <= 0;  //44 / 208 = 0
    16'b00101100_11010001 : OUT <= 0;  //44 / 209 = 0
    16'b00101100_11010010 : OUT <= 0;  //44 / 210 = 0
    16'b00101100_11010011 : OUT <= 0;  //44 / 211 = 0
    16'b00101100_11010100 : OUT <= 0;  //44 / 212 = 0
    16'b00101100_11010101 : OUT <= 0;  //44 / 213 = 0
    16'b00101100_11010110 : OUT <= 0;  //44 / 214 = 0
    16'b00101100_11010111 : OUT <= 0;  //44 / 215 = 0
    16'b00101100_11011000 : OUT <= 0;  //44 / 216 = 0
    16'b00101100_11011001 : OUT <= 0;  //44 / 217 = 0
    16'b00101100_11011010 : OUT <= 0;  //44 / 218 = 0
    16'b00101100_11011011 : OUT <= 0;  //44 / 219 = 0
    16'b00101100_11011100 : OUT <= 0;  //44 / 220 = 0
    16'b00101100_11011101 : OUT <= 0;  //44 / 221 = 0
    16'b00101100_11011110 : OUT <= 0;  //44 / 222 = 0
    16'b00101100_11011111 : OUT <= 0;  //44 / 223 = 0
    16'b00101100_11100000 : OUT <= 0;  //44 / 224 = 0
    16'b00101100_11100001 : OUT <= 0;  //44 / 225 = 0
    16'b00101100_11100010 : OUT <= 0;  //44 / 226 = 0
    16'b00101100_11100011 : OUT <= 0;  //44 / 227 = 0
    16'b00101100_11100100 : OUT <= 0;  //44 / 228 = 0
    16'b00101100_11100101 : OUT <= 0;  //44 / 229 = 0
    16'b00101100_11100110 : OUT <= 0;  //44 / 230 = 0
    16'b00101100_11100111 : OUT <= 0;  //44 / 231 = 0
    16'b00101100_11101000 : OUT <= 0;  //44 / 232 = 0
    16'b00101100_11101001 : OUT <= 0;  //44 / 233 = 0
    16'b00101100_11101010 : OUT <= 0;  //44 / 234 = 0
    16'b00101100_11101011 : OUT <= 0;  //44 / 235 = 0
    16'b00101100_11101100 : OUT <= 0;  //44 / 236 = 0
    16'b00101100_11101101 : OUT <= 0;  //44 / 237 = 0
    16'b00101100_11101110 : OUT <= 0;  //44 / 238 = 0
    16'b00101100_11101111 : OUT <= 0;  //44 / 239 = 0
    16'b00101100_11110000 : OUT <= 0;  //44 / 240 = 0
    16'b00101100_11110001 : OUT <= 0;  //44 / 241 = 0
    16'b00101100_11110010 : OUT <= 0;  //44 / 242 = 0
    16'b00101100_11110011 : OUT <= 0;  //44 / 243 = 0
    16'b00101100_11110100 : OUT <= 0;  //44 / 244 = 0
    16'b00101100_11110101 : OUT <= 0;  //44 / 245 = 0
    16'b00101100_11110110 : OUT <= 0;  //44 / 246 = 0
    16'b00101100_11110111 : OUT <= 0;  //44 / 247 = 0
    16'b00101100_11111000 : OUT <= 0;  //44 / 248 = 0
    16'b00101100_11111001 : OUT <= 0;  //44 / 249 = 0
    16'b00101100_11111010 : OUT <= 0;  //44 / 250 = 0
    16'b00101100_11111011 : OUT <= 0;  //44 / 251 = 0
    16'b00101100_11111100 : OUT <= 0;  //44 / 252 = 0
    16'b00101100_11111101 : OUT <= 0;  //44 / 253 = 0
    16'b00101100_11111110 : OUT <= 0;  //44 / 254 = 0
    16'b00101100_11111111 : OUT <= 0;  //44 / 255 = 0
    16'b00101101_00000000 : OUT <= 0;  //45 / 0 = 0
    16'b00101101_00000001 : OUT <= 45;  //45 / 1 = 45
    16'b00101101_00000010 : OUT <= 22;  //45 / 2 = 22
    16'b00101101_00000011 : OUT <= 15;  //45 / 3 = 15
    16'b00101101_00000100 : OUT <= 11;  //45 / 4 = 11
    16'b00101101_00000101 : OUT <= 9;  //45 / 5 = 9
    16'b00101101_00000110 : OUT <= 7;  //45 / 6 = 7
    16'b00101101_00000111 : OUT <= 6;  //45 / 7 = 6
    16'b00101101_00001000 : OUT <= 5;  //45 / 8 = 5
    16'b00101101_00001001 : OUT <= 5;  //45 / 9 = 5
    16'b00101101_00001010 : OUT <= 4;  //45 / 10 = 4
    16'b00101101_00001011 : OUT <= 4;  //45 / 11 = 4
    16'b00101101_00001100 : OUT <= 3;  //45 / 12 = 3
    16'b00101101_00001101 : OUT <= 3;  //45 / 13 = 3
    16'b00101101_00001110 : OUT <= 3;  //45 / 14 = 3
    16'b00101101_00001111 : OUT <= 3;  //45 / 15 = 3
    16'b00101101_00010000 : OUT <= 2;  //45 / 16 = 2
    16'b00101101_00010001 : OUT <= 2;  //45 / 17 = 2
    16'b00101101_00010010 : OUT <= 2;  //45 / 18 = 2
    16'b00101101_00010011 : OUT <= 2;  //45 / 19 = 2
    16'b00101101_00010100 : OUT <= 2;  //45 / 20 = 2
    16'b00101101_00010101 : OUT <= 2;  //45 / 21 = 2
    16'b00101101_00010110 : OUT <= 2;  //45 / 22 = 2
    16'b00101101_00010111 : OUT <= 1;  //45 / 23 = 1
    16'b00101101_00011000 : OUT <= 1;  //45 / 24 = 1
    16'b00101101_00011001 : OUT <= 1;  //45 / 25 = 1
    16'b00101101_00011010 : OUT <= 1;  //45 / 26 = 1
    16'b00101101_00011011 : OUT <= 1;  //45 / 27 = 1
    16'b00101101_00011100 : OUT <= 1;  //45 / 28 = 1
    16'b00101101_00011101 : OUT <= 1;  //45 / 29 = 1
    16'b00101101_00011110 : OUT <= 1;  //45 / 30 = 1
    16'b00101101_00011111 : OUT <= 1;  //45 / 31 = 1
    16'b00101101_00100000 : OUT <= 1;  //45 / 32 = 1
    16'b00101101_00100001 : OUT <= 1;  //45 / 33 = 1
    16'b00101101_00100010 : OUT <= 1;  //45 / 34 = 1
    16'b00101101_00100011 : OUT <= 1;  //45 / 35 = 1
    16'b00101101_00100100 : OUT <= 1;  //45 / 36 = 1
    16'b00101101_00100101 : OUT <= 1;  //45 / 37 = 1
    16'b00101101_00100110 : OUT <= 1;  //45 / 38 = 1
    16'b00101101_00100111 : OUT <= 1;  //45 / 39 = 1
    16'b00101101_00101000 : OUT <= 1;  //45 / 40 = 1
    16'b00101101_00101001 : OUT <= 1;  //45 / 41 = 1
    16'b00101101_00101010 : OUT <= 1;  //45 / 42 = 1
    16'b00101101_00101011 : OUT <= 1;  //45 / 43 = 1
    16'b00101101_00101100 : OUT <= 1;  //45 / 44 = 1
    16'b00101101_00101101 : OUT <= 1;  //45 / 45 = 1
    16'b00101101_00101110 : OUT <= 0;  //45 / 46 = 0
    16'b00101101_00101111 : OUT <= 0;  //45 / 47 = 0
    16'b00101101_00110000 : OUT <= 0;  //45 / 48 = 0
    16'b00101101_00110001 : OUT <= 0;  //45 / 49 = 0
    16'b00101101_00110010 : OUT <= 0;  //45 / 50 = 0
    16'b00101101_00110011 : OUT <= 0;  //45 / 51 = 0
    16'b00101101_00110100 : OUT <= 0;  //45 / 52 = 0
    16'b00101101_00110101 : OUT <= 0;  //45 / 53 = 0
    16'b00101101_00110110 : OUT <= 0;  //45 / 54 = 0
    16'b00101101_00110111 : OUT <= 0;  //45 / 55 = 0
    16'b00101101_00111000 : OUT <= 0;  //45 / 56 = 0
    16'b00101101_00111001 : OUT <= 0;  //45 / 57 = 0
    16'b00101101_00111010 : OUT <= 0;  //45 / 58 = 0
    16'b00101101_00111011 : OUT <= 0;  //45 / 59 = 0
    16'b00101101_00111100 : OUT <= 0;  //45 / 60 = 0
    16'b00101101_00111101 : OUT <= 0;  //45 / 61 = 0
    16'b00101101_00111110 : OUT <= 0;  //45 / 62 = 0
    16'b00101101_00111111 : OUT <= 0;  //45 / 63 = 0
    16'b00101101_01000000 : OUT <= 0;  //45 / 64 = 0
    16'b00101101_01000001 : OUT <= 0;  //45 / 65 = 0
    16'b00101101_01000010 : OUT <= 0;  //45 / 66 = 0
    16'b00101101_01000011 : OUT <= 0;  //45 / 67 = 0
    16'b00101101_01000100 : OUT <= 0;  //45 / 68 = 0
    16'b00101101_01000101 : OUT <= 0;  //45 / 69 = 0
    16'b00101101_01000110 : OUT <= 0;  //45 / 70 = 0
    16'b00101101_01000111 : OUT <= 0;  //45 / 71 = 0
    16'b00101101_01001000 : OUT <= 0;  //45 / 72 = 0
    16'b00101101_01001001 : OUT <= 0;  //45 / 73 = 0
    16'b00101101_01001010 : OUT <= 0;  //45 / 74 = 0
    16'b00101101_01001011 : OUT <= 0;  //45 / 75 = 0
    16'b00101101_01001100 : OUT <= 0;  //45 / 76 = 0
    16'b00101101_01001101 : OUT <= 0;  //45 / 77 = 0
    16'b00101101_01001110 : OUT <= 0;  //45 / 78 = 0
    16'b00101101_01001111 : OUT <= 0;  //45 / 79 = 0
    16'b00101101_01010000 : OUT <= 0;  //45 / 80 = 0
    16'b00101101_01010001 : OUT <= 0;  //45 / 81 = 0
    16'b00101101_01010010 : OUT <= 0;  //45 / 82 = 0
    16'b00101101_01010011 : OUT <= 0;  //45 / 83 = 0
    16'b00101101_01010100 : OUT <= 0;  //45 / 84 = 0
    16'b00101101_01010101 : OUT <= 0;  //45 / 85 = 0
    16'b00101101_01010110 : OUT <= 0;  //45 / 86 = 0
    16'b00101101_01010111 : OUT <= 0;  //45 / 87 = 0
    16'b00101101_01011000 : OUT <= 0;  //45 / 88 = 0
    16'b00101101_01011001 : OUT <= 0;  //45 / 89 = 0
    16'b00101101_01011010 : OUT <= 0;  //45 / 90 = 0
    16'b00101101_01011011 : OUT <= 0;  //45 / 91 = 0
    16'b00101101_01011100 : OUT <= 0;  //45 / 92 = 0
    16'b00101101_01011101 : OUT <= 0;  //45 / 93 = 0
    16'b00101101_01011110 : OUT <= 0;  //45 / 94 = 0
    16'b00101101_01011111 : OUT <= 0;  //45 / 95 = 0
    16'b00101101_01100000 : OUT <= 0;  //45 / 96 = 0
    16'b00101101_01100001 : OUT <= 0;  //45 / 97 = 0
    16'b00101101_01100010 : OUT <= 0;  //45 / 98 = 0
    16'b00101101_01100011 : OUT <= 0;  //45 / 99 = 0
    16'b00101101_01100100 : OUT <= 0;  //45 / 100 = 0
    16'b00101101_01100101 : OUT <= 0;  //45 / 101 = 0
    16'b00101101_01100110 : OUT <= 0;  //45 / 102 = 0
    16'b00101101_01100111 : OUT <= 0;  //45 / 103 = 0
    16'b00101101_01101000 : OUT <= 0;  //45 / 104 = 0
    16'b00101101_01101001 : OUT <= 0;  //45 / 105 = 0
    16'b00101101_01101010 : OUT <= 0;  //45 / 106 = 0
    16'b00101101_01101011 : OUT <= 0;  //45 / 107 = 0
    16'b00101101_01101100 : OUT <= 0;  //45 / 108 = 0
    16'b00101101_01101101 : OUT <= 0;  //45 / 109 = 0
    16'b00101101_01101110 : OUT <= 0;  //45 / 110 = 0
    16'b00101101_01101111 : OUT <= 0;  //45 / 111 = 0
    16'b00101101_01110000 : OUT <= 0;  //45 / 112 = 0
    16'b00101101_01110001 : OUT <= 0;  //45 / 113 = 0
    16'b00101101_01110010 : OUT <= 0;  //45 / 114 = 0
    16'b00101101_01110011 : OUT <= 0;  //45 / 115 = 0
    16'b00101101_01110100 : OUT <= 0;  //45 / 116 = 0
    16'b00101101_01110101 : OUT <= 0;  //45 / 117 = 0
    16'b00101101_01110110 : OUT <= 0;  //45 / 118 = 0
    16'b00101101_01110111 : OUT <= 0;  //45 / 119 = 0
    16'b00101101_01111000 : OUT <= 0;  //45 / 120 = 0
    16'b00101101_01111001 : OUT <= 0;  //45 / 121 = 0
    16'b00101101_01111010 : OUT <= 0;  //45 / 122 = 0
    16'b00101101_01111011 : OUT <= 0;  //45 / 123 = 0
    16'b00101101_01111100 : OUT <= 0;  //45 / 124 = 0
    16'b00101101_01111101 : OUT <= 0;  //45 / 125 = 0
    16'b00101101_01111110 : OUT <= 0;  //45 / 126 = 0
    16'b00101101_01111111 : OUT <= 0;  //45 / 127 = 0
    16'b00101101_10000000 : OUT <= 0;  //45 / 128 = 0
    16'b00101101_10000001 : OUT <= 0;  //45 / 129 = 0
    16'b00101101_10000010 : OUT <= 0;  //45 / 130 = 0
    16'b00101101_10000011 : OUT <= 0;  //45 / 131 = 0
    16'b00101101_10000100 : OUT <= 0;  //45 / 132 = 0
    16'b00101101_10000101 : OUT <= 0;  //45 / 133 = 0
    16'b00101101_10000110 : OUT <= 0;  //45 / 134 = 0
    16'b00101101_10000111 : OUT <= 0;  //45 / 135 = 0
    16'b00101101_10001000 : OUT <= 0;  //45 / 136 = 0
    16'b00101101_10001001 : OUT <= 0;  //45 / 137 = 0
    16'b00101101_10001010 : OUT <= 0;  //45 / 138 = 0
    16'b00101101_10001011 : OUT <= 0;  //45 / 139 = 0
    16'b00101101_10001100 : OUT <= 0;  //45 / 140 = 0
    16'b00101101_10001101 : OUT <= 0;  //45 / 141 = 0
    16'b00101101_10001110 : OUT <= 0;  //45 / 142 = 0
    16'b00101101_10001111 : OUT <= 0;  //45 / 143 = 0
    16'b00101101_10010000 : OUT <= 0;  //45 / 144 = 0
    16'b00101101_10010001 : OUT <= 0;  //45 / 145 = 0
    16'b00101101_10010010 : OUT <= 0;  //45 / 146 = 0
    16'b00101101_10010011 : OUT <= 0;  //45 / 147 = 0
    16'b00101101_10010100 : OUT <= 0;  //45 / 148 = 0
    16'b00101101_10010101 : OUT <= 0;  //45 / 149 = 0
    16'b00101101_10010110 : OUT <= 0;  //45 / 150 = 0
    16'b00101101_10010111 : OUT <= 0;  //45 / 151 = 0
    16'b00101101_10011000 : OUT <= 0;  //45 / 152 = 0
    16'b00101101_10011001 : OUT <= 0;  //45 / 153 = 0
    16'b00101101_10011010 : OUT <= 0;  //45 / 154 = 0
    16'b00101101_10011011 : OUT <= 0;  //45 / 155 = 0
    16'b00101101_10011100 : OUT <= 0;  //45 / 156 = 0
    16'b00101101_10011101 : OUT <= 0;  //45 / 157 = 0
    16'b00101101_10011110 : OUT <= 0;  //45 / 158 = 0
    16'b00101101_10011111 : OUT <= 0;  //45 / 159 = 0
    16'b00101101_10100000 : OUT <= 0;  //45 / 160 = 0
    16'b00101101_10100001 : OUT <= 0;  //45 / 161 = 0
    16'b00101101_10100010 : OUT <= 0;  //45 / 162 = 0
    16'b00101101_10100011 : OUT <= 0;  //45 / 163 = 0
    16'b00101101_10100100 : OUT <= 0;  //45 / 164 = 0
    16'b00101101_10100101 : OUT <= 0;  //45 / 165 = 0
    16'b00101101_10100110 : OUT <= 0;  //45 / 166 = 0
    16'b00101101_10100111 : OUT <= 0;  //45 / 167 = 0
    16'b00101101_10101000 : OUT <= 0;  //45 / 168 = 0
    16'b00101101_10101001 : OUT <= 0;  //45 / 169 = 0
    16'b00101101_10101010 : OUT <= 0;  //45 / 170 = 0
    16'b00101101_10101011 : OUT <= 0;  //45 / 171 = 0
    16'b00101101_10101100 : OUT <= 0;  //45 / 172 = 0
    16'b00101101_10101101 : OUT <= 0;  //45 / 173 = 0
    16'b00101101_10101110 : OUT <= 0;  //45 / 174 = 0
    16'b00101101_10101111 : OUT <= 0;  //45 / 175 = 0
    16'b00101101_10110000 : OUT <= 0;  //45 / 176 = 0
    16'b00101101_10110001 : OUT <= 0;  //45 / 177 = 0
    16'b00101101_10110010 : OUT <= 0;  //45 / 178 = 0
    16'b00101101_10110011 : OUT <= 0;  //45 / 179 = 0
    16'b00101101_10110100 : OUT <= 0;  //45 / 180 = 0
    16'b00101101_10110101 : OUT <= 0;  //45 / 181 = 0
    16'b00101101_10110110 : OUT <= 0;  //45 / 182 = 0
    16'b00101101_10110111 : OUT <= 0;  //45 / 183 = 0
    16'b00101101_10111000 : OUT <= 0;  //45 / 184 = 0
    16'b00101101_10111001 : OUT <= 0;  //45 / 185 = 0
    16'b00101101_10111010 : OUT <= 0;  //45 / 186 = 0
    16'b00101101_10111011 : OUT <= 0;  //45 / 187 = 0
    16'b00101101_10111100 : OUT <= 0;  //45 / 188 = 0
    16'b00101101_10111101 : OUT <= 0;  //45 / 189 = 0
    16'b00101101_10111110 : OUT <= 0;  //45 / 190 = 0
    16'b00101101_10111111 : OUT <= 0;  //45 / 191 = 0
    16'b00101101_11000000 : OUT <= 0;  //45 / 192 = 0
    16'b00101101_11000001 : OUT <= 0;  //45 / 193 = 0
    16'b00101101_11000010 : OUT <= 0;  //45 / 194 = 0
    16'b00101101_11000011 : OUT <= 0;  //45 / 195 = 0
    16'b00101101_11000100 : OUT <= 0;  //45 / 196 = 0
    16'b00101101_11000101 : OUT <= 0;  //45 / 197 = 0
    16'b00101101_11000110 : OUT <= 0;  //45 / 198 = 0
    16'b00101101_11000111 : OUT <= 0;  //45 / 199 = 0
    16'b00101101_11001000 : OUT <= 0;  //45 / 200 = 0
    16'b00101101_11001001 : OUT <= 0;  //45 / 201 = 0
    16'b00101101_11001010 : OUT <= 0;  //45 / 202 = 0
    16'b00101101_11001011 : OUT <= 0;  //45 / 203 = 0
    16'b00101101_11001100 : OUT <= 0;  //45 / 204 = 0
    16'b00101101_11001101 : OUT <= 0;  //45 / 205 = 0
    16'b00101101_11001110 : OUT <= 0;  //45 / 206 = 0
    16'b00101101_11001111 : OUT <= 0;  //45 / 207 = 0
    16'b00101101_11010000 : OUT <= 0;  //45 / 208 = 0
    16'b00101101_11010001 : OUT <= 0;  //45 / 209 = 0
    16'b00101101_11010010 : OUT <= 0;  //45 / 210 = 0
    16'b00101101_11010011 : OUT <= 0;  //45 / 211 = 0
    16'b00101101_11010100 : OUT <= 0;  //45 / 212 = 0
    16'b00101101_11010101 : OUT <= 0;  //45 / 213 = 0
    16'b00101101_11010110 : OUT <= 0;  //45 / 214 = 0
    16'b00101101_11010111 : OUT <= 0;  //45 / 215 = 0
    16'b00101101_11011000 : OUT <= 0;  //45 / 216 = 0
    16'b00101101_11011001 : OUT <= 0;  //45 / 217 = 0
    16'b00101101_11011010 : OUT <= 0;  //45 / 218 = 0
    16'b00101101_11011011 : OUT <= 0;  //45 / 219 = 0
    16'b00101101_11011100 : OUT <= 0;  //45 / 220 = 0
    16'b00101101_11011101 : OUT <= 0;  //45 / 221 = 0
    16'b00101101_11011110 : OUT <= 0;  //45 / 222 = 0
    16'b00101101_11011111 : OUT <= 0;  //45 / 223 = 0
    16'b00101101_11100000 : OUT <= 0;  //45 / 224 = 0
    16'b00101101_11100001 : OUT <= 0;  //45 / 225 = 0
    16'b00101101_11100010 : OUT <= 0;  //45 / 226 = 0
    16'b00101101_11100011 : OUT <= 0;  //45 / 227 = 0
    16'b00101101_11100100 : OUT <= 0;  //45 / 228 = 0
    16'b00101101_11100101 : OUT <= 0;  //45 / 229 = 0
    16'b00101101_11100110 : OUT <= 0;  //45 / 230 = 0
    16'b00101101_11100111 : OUT <= 0;  //45 / 231 = 0
    16'b00101101_11101000 : OUT <= 0;  //45 / 232 = 0
    16'b00101101_11101001 : OUT <= 0;  //45 / 233 = 0
    16'b00101101_11101010 : OUT <= 0;  //45 / 234 = 0
    16'b00101101_11101011 : OUT <= 0;  //45 / 235 = 0
    16'b00101101_11101100 : OUT <= 0;  //45 / 236 = 0
    16'b00101101_11101101 : OUT <= 0;  //45 / 237 = 0
    16'b00101101_11101110 : OUT <= 0;  //45 / 238 = 0
    16'b00101101_11101111 : OUT <= 0;  //45 / 239 = 0
    16'b00101101_11110000 : OUT <= 0;  //45 / 240 = 0
    16'b00101101_11110001 : OUT <= 0;  //45 / 241 = 0
    16'b00101101_11110010 : OUT <= 0;  //45 / 242 = 0
    16'b00101101_11110011 : OUT <= 0;  //45 / 243 = 0
    16'b00101101_11110100 : OUT <= 0;  //45 / 244 = 0
    16'b00101101_11110101 : OUT <= 0;  //45 / 245 = 0
    16'b00101101_11110110 : OUT <= 0;  //45 / 246 = 0
    16'b00101101_11110111 : OUT <= 0;  //45 / 247 = 0
    16'b00101101_11111000 : OUT <= 0;  //45 / 248 = 0
    16'b00101101_11111001 : OUT <= 0;  //45 / 249 = 0
    16'b00101101_11111010 : OUT <= 0;  //45 / 250 = 0
    16'b00101101_11111011 : OUT <= 0;  //45 / 251 = 0
    16'b00101101_11111100 : OUT <= 0;  //45 / 252 = 0
    16'b00101101_11111101 : OUT <= 0;  //45 / 253 = 0
    16'b00101101_11111110 : OUT <= 0;  //45 / 254 = 0
    16'b00101101_11111111 : OUT <= 0;  //45 / 255 = 0
    16'b00101110_00000000 : OUT <= 0;  //46 / 0 = 0
    16'b00101110_00000001 : OUT <= 46;  //46 / 1 = 46
    16'b00101110_00000010 : OUT <= 23;  //46 / 2 = 23
    16'b00101110_00000011 : OUT <= 15;  //46 / 3 = 15
    16'b00101110_00000100 : OUT <= 11;  //46 / 4 = 11
    16'b00101110_00000101 : OUT <= 9;  //46 / 5 = 9
    16'b00101110_00000110 : OUT <= 7;  //46 / 6 = 7
    16'b00101110_00000111 : OUT <= 6;  //46 / 7 = 6
    16'b00101110_00001000 : OUT <= 5;  //46 / 8 = 5
    16'b00101110_00001001 : OUT <= 5;  //46 / 9 = 5
    16'b00101110_00001010 : OUT <= 4;  //46 / 10 = 4
    16'b00101110_00001011 : OUT <= 4;  //46 / 11 = 4
    16'b00101110_00001100 : OUT <= 3;  //46 / 12 = 3
    16'b00101110_00001101 : OUT <= 3;  //46 / 13 = 3
    16'b00101110_00001110 : OUT <= 3;  //46 / 14 = 3
    16'b00101110_00001111 : OUT <= 3;  //46 / 15 = 3
    16'b00101110_00010000 : OUT <= 2;  //46 / 16 = 2
    16'b00101110_00010001 : OUT <= 2;  //46 / 17 = 2
    16'b00101110_00010010 : OUT <= 2;  //46 / 18 = 2
    16'b00101110_00010011 : OUT <= 2;  //46 / 19 = 2
    16'b00101110_00010100 : OUT <= 2;  //46 / 20 = 2
    16'b00101110_00010101 : OUT <= 2;  //46 / 21 = 2
    16'b00101110_00010110 : OUT <= 2;  //46 / 22 = 2
    16'b00101110_00010111 : OUT <= 2;  //46 / 23 = 2
    16'b00101110_00011000 : OUT <= 1;  //46 / 24 = 1
    16'b00101110_00011001 : OUT <= 1;  //46 / 25 = 1
    16'b00101110_00011010 : OUT <= 1;  //46 / 26 = 1
    16'b00101110_00011011 : OUT <= 1;  //46 / 27 = 1
    16'b00101110_00011100 : OUT <= 1;  //46 / 28 = 1
    16'b00101110_00011101 : OUT <= 1;  //46 / 29 = 1
    16'b00101110_00011110 : OUT <= 1;  //46 / 30 = 1
    16'b00101110_00011111 : OUT <= 1;  //46 / 31 = 1
    16'b00101110_00100000 : OUT <= 1;  //46 / 32 = 1
    16'b00101110_00100001 : OUT <= 1;  //46 / 33 = 1
    16'b00101110_00100010 : OUT <= 1;  //46 / 34 = 1
    16'b00101110_00100011 : OUT <= 1;  //46 / 35 = 1
    16'b00101110_00100100 : OUT <= 1;  //46 / 36 = 1
    16'b00101110_00100101 : OUT <= 1;  //46 / 37 = 1
    16'b00101110_00100110 : OUT <= 1;  //46 / 38 = 1
    16'b00101110_00100111 : OUT <= 1;  //46 / 39 = 1
    16'b00101110_00101000 : OUT <= 1;  //46 / 40 = 1
    16'b00101110_00101001 : OUT <= 1;  //46 / 41 = 1
    16'b00101110_00101010 : OUT <= 1;  //46 / 42 = 1
    16'b00101110_00101011 : OUT <= 1;  //46 / 43 = 1
    16'b00101110_00101100 : OUT <= 1;  //46 / 44 = 1
    16'b00101110_00101101 : OUT <= 1;  //46 / 45 = 1
    16'b00101110_00101110 : OUT <= 1;  //46 / 46 = 1
    16'b00101110_00101111 : OUT <= 0;  //46 / 47 = 0
    16'b00101110_00110000 : OUT <= 0;  //46 / 48 = 0
    16'b00101110_00110001 : OUT <= 0;  //46 / 49 = 0
    16'b00101110_00110010 : OUT <= 0;  //46 / 50 = 0
    16'b00101110_00110011 : OUT <= 0;  //46 / 51 = 0
    16'b00101110_00110100 : OUT <= 0;  //46 / 52 = 0
    16'b00101110_00110101 : OUT <= 0;  //46 / 53 = 0
    16'b00101110_00110110 : OUT <= 0;  //46 / 54 = 0
    16'b00101110_00110111 : OUT <= 0;  //46 / 55 = 0
    16'b00101110_00111000 : OUT <= 0;  //46 / 56 = 0
    16'b00101110_00111001 : OUT <= 0;  //46 / 57 = 0
    16'b00101110_00111010 : OUT <= 0;  //46 / 58 = 0
    16'b00101110_00111011 : OUT <= 0;  //46 / 59 = 0
    16'b00101110_00111100 : OUT <= 0;  //46 / 60 = 0
    16'b00101110_00111101 : OUT <= 0;  //46 / 61 = 0
    16'b00101110_00111110 : OUT <= 0;  //46 / 62 = 0
    16'b00101110_00111111 : OUT <= 0;  //46 / 63 = 0
    16'b00101110_01000000 : OUT <= 0;  //46 / 64 = 0
    16'b00101110_01000001 : OUT <= 0;  //46 / 65 = 0
    16'b00101110_01000010 : OUT <= 0;  //46 / 66 = 0
    16'b00101110_01000011 : OUT <= 0;  //46 / 67 = 0
    16'b00101110_01000100 : OUT <= 0;  //46 / 68 = 0
    16'b00101110_01000101 : OUT <= 0;  //46 / 69 = 0
    16'b00101110_01000110 : OUT <= 0;  //46 / 70 = 0
    16'b00101110_01000111 : OUT <= 0;  //46 / 71 = 0
    16'b00101110_01001000 : OUT <= 0;  //46 / 72 = 0
    16'b00101110_01001001 : OUT <= 0;  //46 / 73 = 0
    16'b00101110_01001010 : OUT <= 0;  //46 / 74 = 0
    16'b00101110_01001011 : OUT <= 0;  //46 / 75 = 0
    16'b00101110_01001100 : OUT <= 0;  //46 / 76 = 0
    16'b00101110_01001101 : OUT <= 0;  //46 / 77 = 0
    16'b00101110_01001110 : OUT <= 0;  //46 / 78 = 0
    16'b00101110_01001111 : OUT <= 0;  //46 / 79 = 0
    16'b00101110_01010000 : OUT <= 0;  //46 / 80 = 0
    16'b00101110_01010001 : OUT <= 0;  //46 / 81 = 0
    16'b00101110_01010010 : OUT <= 0;  //46 / 82 = 0
    16'b00101110_01010011 : OUT <= 0;  //46 / 83 = 0
    16'b00101110_01010100 : OUT <= 0;  //46 / 84 = 0
    16'b00101110_01010101 : OUT <= 0;  //46 / 85 = 0
    16'b00101110_01010110 : OUT <= 0;  //46 / 86 = 0
    16'b00101110_01010111 : OUT <= 0;  //46 / 87 = 0
    16'b00101110_01011000 : OUT <= 0;  //46 / 88 = 0
    16'b00101110_01011001 : OUT <= 0;  //46 / 89 = 0
    16'b00101110_01011010 : OUT <= 0;  //46 / 90 = 0
    16'b00101110_01011011 : OUT <= 0;  //46 / 91 = 0
    16'b00101110_01011100 : OUT <= 0;  //46 / 92 = 0
    16'b00101110_01011101 : OUT <= 0;  //46 / 93 = 0
    16'b00101110_01011110 : OUT <= 0;  //46 / 94 = 0
    16'b00101110_01011111 : OUT <= 0;  //46 / 95 = 0
    16'b00101110_01100000 : OUT <= 0;  //46 / 96 = 0
    16'b00101110_01100001 : OUT <= 0;  //46 / 97 = 0
    16'b00101110_01100010 : OUT <= 0;  //46 / 98 = 0
    16'b00101110_01100011 : OUT <= 0;  //46 / 99 = 0
    16'b00101110_01100100 : OUT <= 0;  //46 / 100 = 0
    16'b00101110_01100101 : OUT <= 0;  //46 / 101 = 0
    16'b00101110_01100110 : OUT <= 0;  //46 / 102 = 0
    16'b00101110_01100111 : OUT <= 0;  //46 / 103 = 0
    16'b00101110_01101000 : OUT <= 0;  //46 / 104 = 0
    16'b00101110_01101001 : OUT <= 0;  //46 / 105 = 0
    16'b00101110_01101010 : OUT <= 0;  //46 / 106 = 0
    16'b00101110_01101011 : OUT <= 0;  //46 / 107 = 0
    16'b00101110_01101100 : OUT <= 0;  //46 / 108 = 0
    16'b00101110_01101101 : OUT <= 0;  //46 / 109 = 0
    16'b00101110_01101110 : OUT <= 0;  //46 / 110 = 0
    16'b00101110_01101111 : OUT <= 0;  //46 / 111 = 0
    16'b00101110_01110000 : OUT <= 0;  //46 / 112 = 0
    16'b00101110_01110001 : OUT <= 0;  //46 / 113 = 0
    16'b00101110_01110010 : OUT <= 0;  //46 / 114 = 0
    16'b00101110_01110011 : OUT <= 0;  //46 / 115 = 0
    16'b00101110_01110100 : OUT <= 0;  //46 / 116 = 0
    16'b00101110_01110101 : OUT <= 0;  //46 / 117 = 0
    16'b00101110_01110110 : OUT <= 0;  //46 / 118 = 0
    16'b00101110_01110111 : OUT <= 0;  //46 / 119 = 0
    16'b00101110_01111000 : OUT <= 0;  //46 / 120 = 0
    16'b00101110_01111001 : OUT <= 0;  //46 / 121 = 0
    16'b00101110_01111010 : OUT <= 0;  //46 / 122 = 0
    16'b00101110_01111011 : OUT <= 0;  //46 / 123 = 0
    16'b00101110_01111100 : OUT <= 0;  //46 / 124 = 0
    16'b00101110_01111101 : OUT <= 0;  //46 / 125 = 0
    16'b00101110_01111110 : OUT <= 0;  //46 / 126 = 0
    16'b00101110_01111111 : OUT <= 0;  //46 / 127 = 0
    16'b00101110_10000000 : OUT <= 0;  //46 / 128 = 0
    16'b00101110_10000001 : OUT <= 0;  //46 / 129 = 0
    16'b00101110_10000010 : OUT <= 0;  //46 / 130 = 0
    16'b00101110_10000011 : OUT <= 0;  //46 / 131 = 0
    16'b00101110_10000100 : OUT <= 0;  //46 / 132 = 0
    16'b00101110_10000101 : OUT <= 0;  //46 / 133 = 0
    16'b00101110_10000110 : OUT <= 0;  //46 / 134 = 0
    16'b00101110_10000111 : OUT <= 0;  //46 / 135 = 0
    16'b00101110_10001000 : OUT <= 0;  //46 / 136 = 0
    16'b00101110_10001001 : OUT <= 0;  //46 / 137 = 0
    16'b00101110_10001010 : OUT <= 0;  //46 / 138 = 0
    16'b00101110_10001011 : OUT <= 0;  //46 / 139 = 0
    16'b00101110_10001100 : OUT <= 0;  //46 / 140 = 0
    16'b00101110_10001101 : OUT <= 0;  //46 / 141 = 0
    16'b00101110_10001110 : OUT <= 0;  //46 / 142 = 0
    16'b00101110_10001111 : OUT <= 0;  //46 / 143 = 0
    16'b00101110_10010000 : OUT <= 0;  //46 / 144 = 0
    16'b00101110_10010001 : OUT <= 0;  //46 / 145 = 0
    16'b00101110_10010010 : OUT <= 0;  //46 / 146 = 0
    16'b00101110_10010011 : OUT <= 0;  //46 / 147 = 0
    16'b00101110_10010100 : OUT <= 0;  //46 / 148 = 0
    16'b00101110_10010101 : OUT <= 0;  //46 / 149 = 0
    16'b00101110_10010110 : OUT <= 0;  //46 / 150 = 0
    16'b00101110_10010111 : OUT <= 0;  //46 / 151 = 0
    16'b00101110_10011000 : OUT <= 0;  //46 / 152 = 0
    16'b00101110_10011001 : OUT <= 0;  //46 / 153 = 0
    16'b00101110_10011010 : OUT <= 0;  //46 / 154 = 0
    16'b00101110_10011011 : OUT <= 0;  //46 / 155 = 0
    16'b00101110_10011100 : OUT <= 0;  //46 / 156 = 0
    16'b00101110_10011101 : OUT <= 0;  //46 / 157 = 0
    16'b00101110_10011110 : OUT <= 0;  //46 / 158 = 0
    16'b00101110_10011111 : OUT <= 0;  //46 / 159 = 0
    16'b00101110_10100000 : OUT <= 0;  //46 / 160 = 0
    16'b00101110_10100001 : OUT <= 0;  //46 / 161 = 0
    16'b00101110_10100010 : OUT <= 0;  //46 / 162 = 0
    16'b00101110_10100011 : OUT <= 0;  //46 / 163 = 0
    16'b00101110_10100100 : OUT <= 0;  //46 / 164 = 0
    16'b00101110_10100101 : OUT <= 0;  //46 / 165 = 0
    16'b00101110_10100110 : OUT <= 0;  //46 / 166 = 0
    16'b00101110_10100111 : OUT <= 0;  //46 / 167 = 0
    16'b00101110_10101000 : OUT <= 0;  //46 / 168 = 0
    16'b00101110_10101001 : OUT <= 0;  //46 / 169 = 0
    16'b00101110_10101010 : OUT <= 0;  //46 / 170 = 0
    16'b00101110_10101011 : OUT <= 0;  //46 / 171 = 0
    16'b00101110_10101100 : OUT <= 0;  //46 / 172 = 0
    16'b00101110_10101101 : OUT <= 0;  //46 / 173 = 0
    16'b00101110_10101110 : OUT <= 0;  //46 / 174 = 0
    16'b00101110_10101111 : OUT <= 0;  //46 / 175 = 0
    16'b00101110_10110000 : OUT <= 0;  //46 / 176 = 0
    16'b00101110_10110001 : OUT <= 0;  //46 / 177 = 0
    16'b00101110_10110010 : OUT <= 0;  //46 / 178 = 0
    16'b00101110_10110011 : OUT <= 0;  //46 / 179 = 0
    16'b00101110_10110100 : OUT <= 0;  //46 / 180 = 0
    16'b00101110_10110101 : OUT <= 0;  //46 / 181 = 0
    16'b00101110_10110110 : OUT <= 0;  //46 / 182 = 0
    16'b00101110_10110111 : OUT <= 0;  //46 / 183 = 0
    16'b00101110_10111000 : OUT <= 0;  //46 / 184 = 0
    16'b00101110_10111001 : OUT <= 0;  //46 / 185 = 0
    16'b00101110_10111010 : OUT <= 0;  //46 / 186 = 0
    16'b00101110_10111011 : OUT <= 0;  //46 / 187 = 0
    16'b00101110_10111100 : OUT <= 0;  //46 / 188 = 0
    16'b00101110_10111101 : OUT <= 0;  //46 / 189 = 0
    16'b00101110_10111110 : OUT <= 0;  //46 / 190 = 0
    16'b00101110_10111111 : OUT <= 0;  //46 / 191 = 0
    16'b00101110_11000000 : OUT <= 0;  //46 / 192 = 0
    16'b00101110_11000001 : OUT <= 0;  //46 / 193 = 0
    16'b00101110_11000010 : OUT <= 0;  //46 / 194 = 0
    16'b00101110_11000011 : OUT <= 0;  //46 / 195 = 0
    16'b00101110_11000100 : OUT <= 0;  //46 / 196 = 0
    16'b00101110_11000101 : OUT <= 0;  //46 / 197 = 0
    16'b00101110_11000110 : OUT <= 0;  //46 / 198 = 0
    16'b00101110_11000111 : OUT <= 0;  //46 / 199 = 0
    16'b00101110_11001000 : OUT <= 0;  //46 / 200 = 0
    16'b00101110_11001001 : OUT <= 0;  //46 / 201 = 0
    16'b00101110_11001010 : OUT <= 0;  //46 / 202 = 0
    16'b00101110_11001011 : OUT <= 0;  //46 / 203 = 0
    16'b00101110_11001100 : OUT <= 0;  //46 / 204 = 0
    16'b00101110_11001101 : OUT <= 0;  //46 / 205 = 0
    16'b00101110_11001110 : OUT <= 0;  //46 / 206 = 0
    16'b00101110_11001111 : OUT <= 0;  //46 / 207 = 0
    16'b00101110_11010000 : OUT <= 0;  //46 / 208 = 0
    16'b00101110_11010001 : OUT <= 0;  //46 / 209 = 0
    16'b00101110_11010010 : OUT <= 0;  //46 / 210 = 0
    16'b00101110_11010011 : OUT <= 0;  //46 / 211 = 0
    16'b00101110_11010100 : OUT <= 0;  //46 / 212 = 0
    16'b00101110_11010101 : OUT <= 0;  //46 / 213 = 0
    16'b00101110_11010110 : OUT <= 0;  //46 / 214 = 0
    16'b00101110_11010111 : OUT <= 0;  //46 / 215 = 0
    16'b00101110_11011000 : OUT <= 0;  //46 / 216 = 0
    16'b00101110_11011001 : OUT <= 0;  //46 / 217 = 0
    16'b00101110_11011010 : OUT <= 0;  //46 / 218 = 0
    16'b00101110_11011011 : OUT <= 0;  //46 / 219 = 0
    16'b00101110_11011100 : OUT <= 0;  //46 / 220 = 0
    16'b00101110_11011101 : OUT <= 0;  //46 / 221 = 0
    16'b00101110_11011110 : OUT <= 0;  //46 / 222 = 0
    16'b00101110_11011111 : OUT <= 0;  //46 / 223 = 0
    16'b00101110_11100000 : OUT <= 0;  //46 / 224 = 0
    16'b00101110_11100001 : OUT <= 0;  //46 / 225 = 0
    16'b00101110_11100010 : OUT <= 0;  //46 / 226 = 0
    16'b00101110_11100011 : OUT <= 0;  //46 / 227 = 0
    16'b00101110_11100100 : OUT <= 0;  //46 / 228 = 0
    16'b00101110_11100101 : OUT <= 0;  //46 / 229 = 0
    16'b00101110_11100110 : OUT <= 0;  //46 / 230 = 0
    16'b00101110_11100111 : OUT <= 0;  //46 / 231 = 0
    16'b00101110_11101000 : OUT <= 0;  //46 / 232 = 0
    16'b00101110_11101001 : OUT <= 0;  //46 / 233 = 0
    16'b00101110_11101010 : OUT <= 0;  //46 / 234 = 0
    16'b00101110_11101011 : OUT <= 0;  //46 / 235 = 0
    16'b00101110_11101100 : OUT <= 0;  //46 / 236 = 0
    16'b00101110_11101101 : OUT <= 0;  //46 / 237 = 0
    16'b00101110_11101110 : OUT <= 0;  //46 / 238 = 0
    16'b00101110_11101111 : OUT <= 0;  //46 / 239 = 0
    16'b00101110_11110000 : OUT <= 0;  //46 / 240 = 0
    16'b00101110_11110001 : OUT <= 0;  //46 / 241 = 0
    16'b00101110_11110010 : OUT <= 0;  //46 / 242 = 0
    16'b00101110_11110011 : OUT <= 0;  //46 / 243 = 0
    16'b00101110_11110100 : OUT <= 0;  //46 / 244 = 0
    16'b00101110_11110101 : OUT <= 0;  //46 / 245 = 0
    16'b00101110_11110110 : OUT <= 0;  //46 / 246 = 0
    16'b00101110_11110111 : OUT <= 0;  //46 / 247 = 0
    16'b00101110_11111000 : OUT <= 0;  //46 / 248 = 0
    16'b00101110_11111001 : OUT <= 0;  //46 / 249 = 0
    16'b00101110_11111010 : OUT <= 0;  //46 / 250 = 0
    16'b00101110_11111011 : OUT <= 0;  //46 / 251 = 0
    16'b00101110_11111100 : OUT <= 0;  //46 / 252 = 0
    16'b00101110_11111101 : OUT <= 0;  //46 / 253 = 0
    16'b00101110_11111110 : OUT <= 0;  //46 / 254 = 0
    16'b00101110_11111111 : OUT <= 0;  //46 / 255 = 0
    16'b00101111_00000000 : OUT <= 0;  //47 / 0 = 0
    16'b00101111_00000001 : OUT <= 47;  //47 / 1 = 47
    16'b00101111_00000010 : OUT <= 23;  //47 / 2 = 23
    16'b00101111_00000011 : OUT <= 15;  //47 / 3 = 15
    16'b00101111_00000100 : OUT <= 11;  //47 / 4 = 11
    16'b00101111_00000101 : OUT <= 9;  //47 / 5 = 9
    16'b00101111_00000110 : OUT <= 7;  //47 / 6 = 7
    16'b00101111_00000111 : OUT <= 6;  //47 / 7 = 6
    16'b00101111_00001000 : OUT <= 5;  //47 / 8 = 5
    16'b00101111_00001001 : OUT <= 5;  //47 / 9 = 5
    16'b00101111_00001010 : OUT <= 4;  //47 / 10 = 4
    16'b00101111_00001011 : OUT <= 4;  //47 / 11 = 4
    16'b00101111_00001100 : OUT <= 3;  //47 / 12 = 3
    16'b00101111_00001101 : OUT <= 3;  //47 / 13 = 3
    16'b00101111_00001110 : OUT <= 3;  //47 / 14 = 3
    16'b00101111_00001111 : OUT <= 3;  //47 / 15 = 3
    16'b00101111_00010000 : OUT <= 2;  //47 / 16 = 2
    16'b00101111_00010001 : OUT <= 2;  //47 / 17 = 2
    16'b00101111_00010010 : OUT <= 2;  //47 / 18 = 2
    16'b00101111_00010011 : OUT <= 2;  //47 / 19 = 2
    16'b00101111_00010100 : OUT <= 2;  //47 / 20 = 2
    16'b00101111_00010101 : OUT <= 2;  //47 / 21 = 2
    16'b00101111_00010110 : OUT <= 2;  //47 / 22 = 2
    16'b00101111_00010111 : OUT <= 2;  //47 / 23 = 2
    16'b00101111_00011000 : OUT <= 1;  //47 / 24 = 1
    16'b00101111_00011001 : OUT <= 1;  //47 / 25 = 1
    16'b00101111_00011010 : OUT <= 1;  //47 / 26 = 1
    16'b00101111_00011011 : OUT <= 1;  //47 / 27 = 1
    16'b00101111_00011100 : OUT <= 1;  //47 / 28 = 1
    16'b00101111_00011101 : OUT <= 1;  //47 / 29 = 1
    16'b00101111_00011110 : OUT <= 1;  //47 / 30 = 1
    16'b00101111_00011111 : OUT <= 1;  //47 / 31 = 1
    16'b00101111_00100000 : OUT <= 1;  //47 / 32 = 1
    16'b00101111_00100001 : OUT <= 1;  //47 / 33 = 1
    16'b00101111_00100010 : OUT <= 1;  //47 / 34 = 1
    16'b00101111_00100011 : OUT <= 1;  //47 / 35 = 1
    16'b00101111_00100100 : OUT <= 1;  //47 / 36 = 1
    16'b00101111_00100101 : OUT <= 1;  //47 / 37 = 1
    16'b00101111_00100110 : OUT <= 1;  //47 / 38 = 1
    16'b00101111_00100111 : OUT <= 1;  //47 / 39 = 1
    16'b00101111_00101000 : OUT <= 1;  //47 / 40 = 1
    16'b00101111_00101001 : OUT <= 1;  //47 / 41 = 1
    16'b00101111_00101010 : OUT <= 1;  //47 / 42 = 1
    16'b00101111_00101011 : OUT <= 1;  //47 / 43 = 1
    16'b00101111_00101100 : OUT <= 1;  //47 / 44 = 1
    16'b00101111_00101101 : OUT <= 1;  //47 / 45 = 1
    16'b00101111_00101110 : OUT <= 1;  //47 / 46 = 1
    16'b00101111_00101111 : OUT <= 1;  //47 / 47 = 1
    16'b00101111_00110000 : OUT <= 0;  //47 / 48 = 0
    16'b00101111_00110001 : OUT <= 0;  //47 / 49 = 0
    16'b00101111_00110010 : OUT <= 0;  //47 / 50 = 0
    16'b00101111_00110011 : OUT <= 0;  //47 / 51 = 0
    16'b00101111_00110100 : OUT <= 0;  //47 / 52 = 0
    16'b00101111_00110101 : OUT <= 0;  //47 / 53 = 0
    16'b00101111_00110110 : OUT <= 0;  //47 / 54 = 0
    16'b00101111_00110111 : OUT <= 0;  //47 / 55 = 0
    16'b00101111_00111000 : OUT <= 0;  //47 / 56 = 0
    16'b00101111_00111001 : OUT <= 0;  //47 / 57 = 0
    16'b00101111_00111010 : OUT <= 0;  //47 / 58 = 0
    16'b00101111_00111011 : OUT <= 0;  //47 / 59 = 0
    16'b00101111_00111100 : OUT <= 0;  //47 / 60 = 0
    16'b00101111_00111101 : OUT <= 0;  //47 / 61 = 0
    16'b00101111_00111110 : OUT <= 0;  //47 / 62 = 0
    16'b00101111_00111111 : OUT <= 0;  //47 / 63 = 0
    16'b00101111_01000000 : OUT <= 0;  //47 / 64 = 0
    16'b00101111_01000001 : OUT <= 0;  //47 / 65 = 0
    16'b00101111_01000010 : OUT <= 0;  //47 / 66 = 0
    16'b00101111_01000011 : OUT <= 0;  //47 / 67 = 0
    16'b00101111_01000100 : OUT <= 0;  //47 / 68 = 0
    16'b00101111_01000101 : OUT <= 0;  //47 / 69 = 0
    16'b00101111_01000110 : OUT <= 0;  //47 / 70 = 0
    16'b00101111_01000111 : OUT <= 0;  //47 / 71 = 0
    16'b00101111_01001000 : OUT <= 0;  //47 / 72 = 0
    16'b00101111_01001001 : OUT <= 0;  //47 / 73 = 0
    16'b00101111_01001010 : OUT <= 0;  //47 / 74 = 0
    16'b00101111_01001011 : OUT <= 0;  //47 / 75 = 0
    16'b00101111_01001100 : OUT <= 0;  //47 / 76 = 0
    16'b00101111_01001101 : OUT <= 0;  //47 / 77 = 0
    16'b00101111_01001110 : OUT <= 0;  //47 / 78 = 0
    16'b00101111_01001111 : OUT <= 0;  //47 / 79 = 0
    16'b00101111_01010000 : OUT <= 0;  //47 / 80 = 0
    16'b00101111_01010001 : OUT <= 0;  //47 / 81 = 0
    16'b00101111_01010010 : OUT <= 0;  //47 / 82 = 0
    16'b00101111_01010011 : OUT <= 0;  //47 / 83 = 0
    16'b00101111_01010100 : OUT <= 0;  //47 / 84 = 0
    16'b00101111_01010101 : OUT <= 0;  //47 / 85 = 0
    16'b00101111_01010110 : OUT <= 0;  //47 / 86 = 0
    16'b00101111_01010111 : OUT <= 0;  //47 / 87 = 0
    16'b00101111_01011000 : OUT <= 0;  //47 / 88 = 0
    16'b00101111_01011001 : OUT <= 0;  //47 / 89 = 0
    16'b00101111_01011010 : OUT <= 0;  //47 / 90 = 0
    16'b00101111_01011011 : OUT <= 0;  //47 / 91 = 0
    16'b00101111_01011100 : OUT <= 0;  //47 / 92 = 0
    16'b00101111_01011101 : OUT <= 0;  //47 / 93 = 0
    16'b00101111_01011110 : OUT <= 0;  //47 / 94 = 0
    16'b00101111_01011111 : OUT <= 0;  //47 / 95 = 0
    16'b00101111_01100000 : OUT <= 0;  //47 / 96 = 0
    16'b00101111_01100001 : OUT <= 0;  //47 / 97 = 0
    16'b00101111_01100010 : OUT <= 0;  //47 / 98 = 0
    16'b00101111_01100011 : OUT <= 0;  //47 / 99 = 0
    16'b00101111_01100100 : OUT <= 0;  //47 / 100 = 0
    16'b00101111_01100101 : OUT <= 0;  //47 / 101 = 0
    16'b00101111_01100110 : OUT <= 0;  //47 / 102 = 0
    16'b00101111_01100111 : OUT <= 0;  //47 / 103 = 0
    16'b00101111_01101000 : OUT <= 0;  //47 / 104 = 0
    16'b00101111_01101001 : OUT <= 0;  //47 / 105 = 0
    16'b00101111_01101010 : OUT <= 0;  //47 / 106 = 0
    16'b00101111_01101011 : OUT <= 0;  //47 / 107 = 0
    16'b00101111_01101100 : OUT <= 0;  //47 / 108 = 0
    16'b00101111_01101101 : OUT <= 0;  //47 / 109 = 0
    16'b00101111_01101110 : OUT <= 0;  //47 / 110 = 0
    16'b00101111_01101111 : OUT <= 0;  //47 / 111 = 0
    16'b00101111_01110000 : OUT <= 0;  //47 / 112 = 0
    16'b00101111_01110001 : OUT <= 0;  //47 / 113 = 0
    16'b00101111_01110010 : OUT <= 0;  //47 / 114 = 0
    16'b00101111_01110011 : OUT <= 0;  //47 / 115 = 0
    16'b00101111_01110100 : OUT <= 0;  //47 / 116 = 0
    16'b00101111_01110101 : OUT <= 0;  //47 / 117 = 0
    16'b00101111_01110110 : OUT <= 0;  //47 / 118 = 0
    16'b00101111_01110111 : OUT <= 0;  //47 / 119 = 0
    16'b00101111_01111000 : OUT <= 0;  //47 / 120 = 0
    16'b00101111_01111001 : OUT <= 0;  //47 / 121 = 0
    16'b00101111_01111010 : OUT <= 0;  //47 / 122 = 0
    16'b00101111_01111011 : OUT <= 0;  //47 / 123 = 0
    16'b00101111_01111100 : OUT <= 0;  //47 / 124 = 0
    16'b00101111_01111101 : OUT <= 0;  //47 / 125 = 0
    16'b00101111_01111110 : OUT <= 0;  //47 / 126 = 0
    16'b00101111_01111111 : OUT <= 0;  //47 / 127 = 0
    16'b00101111_10000000 : OUT <= 0;  //47 / 128 = 0
    16'b00101111_10000001 : OUT <= 0;  //47 / 129 = 0
    16'b00101111_10000010 : OUT <= 0;  //47 / 130 = 0
    16'b00101111_10000011 : OUT <= 0;  //47 / 131 = 0
    16'b00101111_10000100 : OUT <= 0;  //47 / 132 = 0
    16'b00101111_10000101 : OUT <= 0;  //47 / 133 = 0
    16'b00101111_10000110 : OUT <= 0;  //47 / 134 = 0
    16'b00101111_10000111 : OUT <= 0;  //47 / 135 = 0
    16'b00101111_10001000 : OUT <= 0;  //47 / 136 = 0
    16'b00101111_10001001 : OUT <= 0;  //47 / 137 = 0
    16'b00101111_10001010 : OUT <= 0;  //47 / 138 = 0
    16'b00101111_10001011 : OUT <= 0;  //47 / 139 = 0
    16'b00101111_10001100 : OUT <= 0;  //47 / 140 = 0
    16'b00101111_10001101 : OUT <= 0;  //47 / 141 = 0
    16'b00101111_10001110 : OUT <= 0;  //47 / 142 = 0
    16'b00101111_10001111 : OUT <= 0;  //47 / 143 = 0
    16'b00101111_10010000 : OUT <= 0;  //47 / 144 = 0
    16'b00101111_10010001 : OUT <= 0;  //47 / 145 = 0
    16'b00101111_10010010 : OUT <= 0;  //47 / 146 = 0
    16'b00101111_10010011 : OUT <= 0;  //47 / 147 = 0
    16'b00101111_10010100 : OUT <= 0;  //47 / 148 = 0
    16'b00101111_10010101 : OUT <= 0;  //47 / 149 = 0
    16'b00101111_10010110 : OUT <= 0;  //47 / 150 = 0
    16'b00101111_10010111 : OUT <= 0;  //47 / 151 = 0
    16'b00101111_10011000 : OUT <= 0;  //47 / 152 = 0
    16'b00101111_10011001 : OUT <= 0;  //47 / 153 = 0
    16'b00101111_10011010 : OUT <= 0;  //47 / 154 = 0
    16'b00101111_10011011 : OUT <= 0;  //47 / 155 = 0
    16'b00101111_10011100 : OUT <= 0;  //47 / 156 = 0
    16'b00101111_10011101 : OUT <= 0;  //47 / 157 = 0
    16'b00101111_10011110 : OUT <= 0;  //47 / 158 = 0
    16'b00101111_10011111 : OUT <= 0;  //47 / 159 = 0
    16'b00101111_10100000 : OUT <= 0;  //47 / 160 = 0
    16'b00101111_10100001 : OUT <= 0;  //47 / 161 = 0
    16'b00101111_10100010 : OUT <= 0;  //47 / 162 = 0
    16'b00101111_10100011 : OUT <= 0;  //47 / 163 = 0
    16'b00101111_10100100 : OUT <= 0;  //47 / 164 = 0
    16'b00101111_10100101 : OUT <= 0;  //47 / 165 = 0
    16'b00101111_10100110 : OUT <= 0;  //47 / 166 = 0
    16'b00101111_10100111 : OUT <= 0;  //47 / 167 = 0
    16'b00101111_10101000 : OUT <= 0;  //47 / 168 = 0
    16'b00101111_10101001 : OUT <= 0;  //47 / 169 = 0
    16'b00101111_10101010 : OUT <= 0;  //47 / 170 = 0
    16'b00101111_10101011 : OUT <= 0;  //47 / 171 = 0
    16'b00101111_10101100 : OUT <= 0;  //47 / 172 = 0
    16'b00101111_10101101 : OUT <= 0;  //47 / 173 = 0
    16'b00101111_10101110 : OUT <= 0;  //47 / 174 = 0
    16'b00101111_10101111 : OUT <= 0;  //47 / 175 = 0
    16'b00101111_10110000 : OUT <= 0;  //47 / 176 = 0
    16'b00101111_10110001 : OUT <= 0;  //47 / 177 = 0
    16'b00101111_10110010 : OUT <= 0;  //47 / 178 = 0
    16'b00101111_10110011 : OUT <= 0;  //47 / 179 = 0
    16'b00101111_10110100 : OUT <= 0;  //47 / 180 = 0
    16'b00101111_10110101 : OUT <= 0;  //47 / 181 = 0
    16'b00101111_10110110 : OUT <= 0;  //47 / 182 = 0
    16'b00101111_10110111 : OUT <= 0;  //47 / 183 = 0
    16'b00101111_10111000 : OUT <= 0;  //47 / 184 = 0
    16'b00101111_10111001 : OUT <= 0;  //47 / 185 = 0
    16'b00101111_10111010 : OUT <= 0;  //47 / 186 = 0
    16'b00101111_10111011 : OUT <= 0;  //47 / 187 = 0
    16'b00101111_10111100 : OUT <= 0;  //47 / 188 = 0
    16'b00101111_10111101 : OUT <= 0;  //47 / 189 = 0
    16'b00101111_10111110 : OUT <= 0;  //47 / 190 = 0
    16'b00101111_10111111 : OUT <= 0;  //47 / 191 = 0
    16'b00101111_11000000 : OUT <= 0;  //47 / 192 = 0
    16'b00101111_11000001 : OUT <= 0;  //47 / 193 = 0
    16'b00101111_11000010 : OUT <= 0;  //47 / 194 = 0
    16'b00101111_11000011 : OUT <= 0;  //47 / 195 = 0
    16'b00101111_11000100 : OUT <= 0;  //47 / 196 = 0
    16'b00101111_11000101 : OUT <= 0;  //47 / 197 = 0
    16'b00101111_11000110 : OUT <= 0;  //47 / 198 = 0
    16'b00101111_11000111 : OUT <= 0;  //47 / 199 = 0
    16'b00101111_11001000 : OUT <= 0;  //47 / 200 = 0
    16'b00101111_11001001 : OUT <= 0;  //47 / 201 = 0
    16'b00101111_11001010 : OUT <= 0;  //47 / 202 = 0
    16'b00101111_11001011 : OUT <= 0;  //47 / 203 = 0
    16'b00101111_11001100 : OUT <= 0;  //47 / 204 = 0
    16'b00101111_11001101 : OUT <= 0;  //47 / 205 = 0
    16'b00101111_11001110 : OUT <= 0;  //47 / 206 = 0
    16'b00101111_11001111 : OUT <= 0;  //47 / 207 = 0
    16'b00101111_11010000 : OUT <= 0;  //47 / 208 = 0
    16'b00101111_11010001 : OUT <= 0;  //47 / 209 = 0
    16'b00101111_11010010 : OUT <= 0;  //47 / 210 = 0
    16'b00101111_11010011 : OUT <= 0;  //47 / 211 = 0
    16'b00101111_11010100 : OUT <= 0;  //47 / 212 = 0
    16'b00101111_11010101 : OUT <= 0;  //47 / 213 = 0
    16'b00101111_11010110 : OUT <= 0;  //47 / 214 = 0
    16'b00101111_11010111 : OUT <= 0;  //47 / 215 = 0
    16'b00101111_11011000 : OUT <= 0;  //47 / 216 = 0
    16'b00101111_11011001 : OUT <= 0;  //47 / 217 = 0
    16'b00101111_11011010 : OUT <= 0;  //47 / 218 = 0
    16'b00101111_11011011 : OUT <= 0;  //47 / 219 = 0
    16'b00101111_11011100 : OUT <= 0;  //47 / 220 = 0
    16'b00101111_11011101 : OUT <= 0;  //47 / 221 = 0
    16'b00101111_11011110 : OUT <= 0;  //47 / 222 = 0
    16'b00101111_11011111 : OUT <= 0;  //47 / 223 = 0
    16'b00101111_11100000 : OUT <= 0;  //47 / 224 = 0
    16'b00101111_11100001 : OUT <= 0;  //47 / 225 = 0
    16'b00101111_11100010 : OUT <= 0;  //47 / 226 = 0
    16'b00101111_11100011 : OUT <= 0;  //47 / 227 = 0
    16'b00101111_11100100 : OUT <= 0;  //47 / 228 = 0
    16'b00101111_11100101 : OUT <= 0;  //47 / 229 = 0
    16'b00101111_11100110 : OUT <= 0;  //47 / 230 = 0
    16'b00101111_11100111 : OUT <= 0;  //47 / 231 = 0
    16'b00101111_11101000 : OUT <= 0;  //47 / 232 = 0
    16'b00101111_11101001 : OUT <= 0;  //47 / 233 = 0
    16'b00101111_11101010 : OUT <= 0;  //47 / 234 = 0
    16'b00101111_11101011 : OUT <= 0;  //47 / 235 = 0
    16'b00101111_11101100 : OUT <= 0;  //47 / 236 = 0
    16'b00101111_11101101 : OUT <= 0;  //47 / 237 = 0
    16'b00101111_11101110 : OUT <= 0;  //47 / 238 = 0
    16'b00101111_11101111 : OUT <= 0;  //47 / 239 = 0
    16'b00101111_11110000 : OUT <= 0;  //47 / 240 = 0
    16'b00101111_11110001 : OUT <= 0;  //47 / 241 = 0
    16'b00101111_11110010 : OUT <= 0;  //47 / 242 = 0
    16'b00101111_11110011 : OUT <= 0;  //47 / 243 = 0
    16'b00101111_11110100 : OUT <= 0;  //47 / 244 = 0
    16'b00101111_11110101 : OUT <= 0;  //47 / 245 = 0
    16'b00101111_11110110 : OUT <= 0;  //47 / 246 = 0
    16'b00101111_11110111 : OUT <= 0;  //47 / 247 = 0
    16'b00101111_11111000 : OUT <= 0;  //47 / 248 = 0
    16'b00101111_11111001 : OUT <= 0;  //47 / 249 = 0
    16'b00101111_11111010 : OUT <= 0;  //47 / 250 = 0
    16'b00101111_11111011 : OUT <= 0;  //47 / 251 = 0
    16'b00101111_11111100 : OUT <= 0;  //47 / 252 = 0
    16'b00101111_11111101 : OUT <= 0;  //47 / 253 = 0
    16'b00101111_11111110 : OUT <= 0;  //47 / 254 = 0
    16'b00101111_11111111 : OUT <= 0;  //47 / 255 = 0
    16'b00110000_00000000 : OUT <= 0;  //48 / 0 = 0
    16'b00110000_00000001 : OUT <= 48;  //48 / 1 = 48
    16'b00110000_00000010 : OUT <= 24;  //48 / 2 = 24
    16'b00110000_00000011 : OUT <= 16;  //48 / 3 = 16
    16'b00110000_00000100 : OUT <= 12;  //48 / 4 = 12
    16'b00110000_00000101 : OUT <= 9;  //48 / 5 = 9
    16'b00110000_00000110 : OUT <= 8;  //48 / 6 = 8
    16'b00110000_00000111 : OUT <= 6;  //48 / 7 = 6
    16'b00110000_00001000 : OUT <= 6;  //48 / 8 = 6
    16'b00110000_00001001 : OUT <= 5;  //48 / 9 = 5
    16'b00110000_00001010 : OUT <= 4;  //48 / 10 = 4
    16'b00110000_00001011 : OUT <= 4;  //48 / 11 = 4
    16'b00110000_00001100 : OUT <= 4;  //48 / 12 = 4
    16'b00110000_00001101 : OUT <= 3;  //48 / 13 = 3
    16'b00110000_00001110 : OUT <= 3;  //48 / 14 = 3
    16'b00110000_00001111 : OUT <= 3;  //48 / 15 = 3
    16'b00110000_00010000 : OUT <= 3;  //48 / 16 = 3
    16'b00110000_00010001 : OUT <= 2;  //48 / 17 = 2
    16'b00110000_00010010 : OUT <= 2;  //48 / 18 = 2
    16'b00110000_00010011 : OUT <= 2;  //48 / 19 = 2
    16'b00110000_00010100 : OUT <= 2;  //48 / 20 = 2
    16'b00110000_00010101 : OUT <= 2;  //48 / 21 = 2
    16'b00110000_00010110 : OUT <= 2;  //48 / 22 = 2
    16'b00110000_00010111 : OUT <= 2;  //48 / 23 = 2
    16'b00110000_00011000 : OUT <= 2;  //48 / 24 = 2
    16'b00110000_00011001 : OUT <= 1;  //48 / 25 = 1
    16'b00110000_00011010 : OUT <= 1;  //48 / 26 = 1
    16'b00110000_00011011 : OUT <= 1;  //48 / 27 = 1
    16'b00110000_00011100 : OUT <= 1;  //48 / 28 = 1
    16'b00110000_00011101 : OUT <= 1;  //48 / 29 = 1
    16'b00110000_00011110 : OUT <= 1;  //48 / 30 = 1
    16'b00110000_00011111 : OUT <= 1;  //48 / 31 = 1
    16'b00110000_00100000 : OUT <= 1;  //48 / 32 = 1
    16'b00110000_00100001 : OUT <= 1;  //48 / 33 = 1
    16'b00110000_00100010 : OUT <= 1;  //48 / 34 = 1
    16'b00110000_00100011 : OUT <= 1;  //48 / 35 = 1
    16'b00110000_00100100 : OUT <= 1;  //48 / 36 = 1
    16'b00110000_00100101 : OUT <= 1;  //48 / 37 = 1
    16'b00110000_00100110 : OUT <= 1;  //48 / 38 = 1
    16'b00110000_00100111 : OUT <= 1;  //48 / 39 = 1
    16'b00110000_00101000 : OUT <= 1;  //48 / 40 = 1
    16'b00110000_00101001 : OUT <= 1;  //48 / 41 = 1
    16'b00110000_00101010 : OUT <= 1;  //48 / 42 = 1
    16'b00110000_00101011 : OUT <= 1;  //48 / 43 = 1
    16'b00110000_00101100 : OUT <= 1;  //48 / 44 = 1
    16'b00110000_00101101 : OUT <= 1;  //48 / 45 = 1
    16'b00110000_00101110 : OUT <= 1;  //48 / 46 = 1
    16'b00110000_00101111 : OUT <= 1;  //48 / 47 = 1
    16'b00110000_00110000 : OUT <= 1;  //48 / 48 = 1
    16'b00110000_00110001 : OUT <= 0;  //48 / 49 = 0
    16'b00110000_00110010 : OUT <= 0;  //48 / 50 = 0
    16'b00110000_00110011 : OUT <= 0;  //48 / 51 = 0
    16'b00110000_00110100 : OUT <= 0;  //48 / 52 = 0
    16'b00110000_00110101 : OUT <= 0;  //48 / 53 = 0
    16'b00110000_00110110 : OUT <= 0;  //48 / 54 = 0
    16'b00110000_00110111 : OUT <= 0;  //48 / 55 = 0
    16'b00110000_00111000 : OUT <= 0;  //48 / 56 = 0
    16'b00110000_00111001 : OUT <= 0;  //48 / 57 = 0
    16'b00110000_00111010 : OUT <= 0;  //48 / 58 = 0
    16'b00110000_00111011 : OUT <= 0;  //48 / 59 = 0
    16'b00110000_00111100 : OUT <= 0;  //48 / 60 = 0
    16'b00110000_00111101 : OUT <= 0;  //48 / 61 = 0
    16'b00110000_00111110 : OUT <= 0;  //48 / 62 = 0
    16'b00110000_00111111 : OUT <= 0;  //48 / 63 = 0
    16'b00110000_01000000 : OUT <= 0;  //48 / 64 = 0
    16'b00110000_01000001 : OUT <= 0;  //48 / 65 = 0
    16'b00110000_01000010 : OUT <= 0;  //48 / 66 = 0
    16'b00110000_01000011 : OUT <= 0;  //48 / 67 = 0
    16'b00110000_01000100 : OUT <= 0;  //48 / 68 = 0
    16'b00110000_01000101 : OUT <= 0;  //48 / 69 = 0
    16'b00110000_01000110 : OUT <= 0;  //48 / 70 = 0
    16'b00110000_01000111 : OUT <= 0;  //48 / 71 = 0
    16'b00110000_01001000 : OUT <= 0;  //48 / 72 = 0
    16'b00110000_01001001 : OUT <= 0;  //48 / 73 = 0
    16'b00110000_01001010 : OUT <= 0;  //48 / 74 = 0
    16'b00110000_01001011 : OUT <= 0;  //48 / 75 = 0
    16'b00110000_01001100 : OUT <= 0;  //48 / 76 = 0
    16'b00110000_01001101 : OUT <= 0;  //48 / 77 = 0
    16'b00110000_01001110 : OUT <= 0;  //48 / 78 = 0
    16'b00110000_01001111 : OUT <= 0;  //48 / 79 = 0
    16'b00110000_01010000 : OUT <= 0;  //48 / 80 = 0
    16'b00110000_01010001 : OUT <= 0;  //48 / 81 = 0
    16'b00110000_01010010 : OUT <= 0;  //48 / 82 = 0
    16'b00110000_01010011 : OUT <= 0;  //48 / 83 = 0
    16'b00110000_01010100 : OUT <= 0;  //48 / 84 = 0
    16'b00110000_01010101 : OUT <= 0;  //48 / 85 = 0
    16'b00110000_01010110 : OUT <= 0;  //48 / 86 = 0
    16'b00110000_01010111 : OUT <= 0;  //48 / 87 = 0
    16'b00110000_01011000 : OUT <= 0;  //48 / 88 = 0
    16'b00110000_01011001 : OUT <= 0;  //48 / 89 = 0
    16'b00110000_01011010 : OUT <= 0;  //48 / 90 = 0
    16'b00110000_01011011 : OUT <= 0;  //48 / 91 = 0
    16'b00110000_01011100 : OUT <= 0;  //48 / 92 = 0
    16'b00110000_01011101 : OUT <= 0;  //48 / 93 = 0
    16'b00110000_01011110 : OUT <= 0;  //48 / 94 = 0
    16'b00110000_01011111 : OUT <= 0;  //48 / 95 = 0
    16'b00110000_01100000 : OUT <= 0;  //48 / 96 = 0
    16'b00110000_01100001 : OUT <= 0;  //48 / 97 = 0
    16'b00110000_01100010 : OUT <= 0;  //48 / 98 = 0
    16'b00110000_01100011 : OUT <= 0;  //48 / 99 = 0
    16'b00110000_01100100 : OUT <= 0;  //48 / 100 = 0
    16'b00110000_01100101 : OUT <= 0;  //48 / 101 = 0
    16'b00110000_01100110 : OUT <= 0;  //48 / 102 = 0
    16'b00110000_01100111 : OUT <= 0;  //48 / 103 = 0
    16'b00110000_01101000 : OUT <= 0;  //48 / 104 = 0
    16'b00110000_01101001 : OUT <= 0;  //48 / 105 = 0
    16'b00110000_01101010 : OUT <= 0;  //48 / 106 = 0
    16'b00110000_01101011 : OUT <= 0;  //48 / 107 = 0
    16'b00110000_01101100 : OUT <= 0;  //48 / 108 = 0
    16'b00110000_01101101 : OUT <= 0;  //48 / 109 = 0
    16'b00110000_01101110 : OUT <= 0;  //48 / 110 = 0
    16'b00110000_01101111 : OUT <= 0;  //48 / 111 = 0
    16'b00110000_01110000 : OUT <= 0;  //48 / 112 = 0
    16'b00110000_01110001 : OUT <= 0;  //48 / 113 = 0
    16'b00110000_01110010 : OUT <= 0;  //48 / 114 = 0
    16'b00110000_01110011 : OUT <= 0;  //48 / 115 = 0
    16'b00110000_01110100 : OUT <= 0;  //48 / 116 = 0
    16'b00110000_01110101 : OUT <= 0;  //48 / 117 = 0
    16'b00110000_01110110 : OUT <= 0;  //48 / 118 = 0
    16'b00110000_01110111 : OUT <= 0;  //48 / 119 = 0
    16'b00110000_01111000 : OUT <= 0;  //48 / 120 = 0
    16'b00110000_01111001 : OUT <= 0;  //48 / 121 = 0
    16'b00110000_01111010 : OUT <= 0;  //48 / 122 = 0
    16'b00110000_01111011 : OUT <= 0;  //48 / 123 = 0
    16'b00110000_01111100 : OUT <= 0;  //48 / 124 = 0
    16'b00110000_01111101 : OUT <= 0;  //48 / 125 = 0
    16'b00110000_01111110 : OUT <= 0;  //48 / 126 = 0
    16'b00110000_01111111 : OUT <= 0;  //48 / 127 = 0
    16'b00110000_10000000 : OUT <= 0;  //48 / 128 = 0
    16'b00110000_10000001 : OUT <= 0;  //48 / 129 = 0
    16'b00110000_10000010 : OUT <= 0;  //48 / 130 = 0
    16'b00110000_10000011 : OUT <= 0;  //48 / 131 = 0
    16'b00110000_10000100 : OUT <= 0;  //48 / 132 = 0
    16'b00110000_10000101 : OUT <= 0;  //48 / 133 = 0
    16'b00110000_10000110 : OUT <= 0;  //48 / 134 = 0
    16'b00110000_10000111 : OUT <= 0;  //48 / 135 = 0
    16'b00110000_10001000 : OUT <= 0;  //48 / 136 = 0
    16'b00110000_10001001 : OUT <= 0;  //48 / 137 = 0
    16'b00110000_10001010 : OUT <= 0;  //48 / 138 = 0
    16'b00110000_10001011 : OUT <= 0;  //48 / 139 = 0
    16'b00110000_10001100 : OUT <= 0;  //48 / 140 = 0
    16'b00110000_10001101 : OUT <= 0;  //48 / 141 = 0
    16'b00110000_10001110 : OUT <= 0;  //48 / 142 = 0
    16'b00110000_10001111 : OUT <= 0;  //48 / 143 = 0
    16'b00110000_10010000 : OUT <= 0;  //48 / 144 = 0
    16'b00110000_10010001 : OUT <= 0;  //48 / 145 = 0
    16'b00110000_10010010 : OUT <= 0;  //48 / 146 = 0
    16'b00110000_10010011 : OUT <= 0;  //48 / 147 = 0
    16'b00110000_10010100 : OUT <= 0;  //48 / 148 = 0
    16'b00110000_10010101 : OUT <= 0;  //48 / 149 = 0
    16'b00110000_10010110 : OUT <= 0;  //48 / 150 = 0
    16'b00110000_10010111 : OUT <= 0;  //48 / 151 = 0
    16'b00110000_10011000 : OUT <= 0;  //48 / 152 = 0
    16'b00110000_10011001 : OUT <= 0;  //48 / 153 = 0
    16'b00110000_10011010 : OUT <= 0;  //48 / 154 = 0
    16'b00110000_10011011 : OUT <= 0;  //48 / 155 = 0
    16'b00110000_10011100 : OUT <= 0;  //48 / 156 = 0
    16'b00110000_10011101 : OUT <= 0;  //48 / 157 = 0
    16'b00110000_10011110 : OUT <= 0;  //48 / 158 = 0
    16'b00110000_10011111 : OUT <= 0;  //48 / 159 = 0
    16'b00110000_10100000 : OUT <= 0;  //48 / 160 = 0
    16'b00110000_10100001 : OUT <= 0;  //48 / 161 = 0
    16'b00110000_10100010 : OUT <= 0;  //48 / 162 = 0
    16'b00110000_10100011 : OUT <= 0;  //48 / 163 = 0
    16'b00110000_10100100 : OUT <= 0;  //48 / 164 = 0
    16'b00110000_10100101 : OUT <= 0;  //48 / 165 = 0
    16'b00110000_10100110 : OUT <= 0;  //48 / 166 = 0
    16'b00110000_10100111 : OUT <= 0;  //48 / 167 = 0
    16'b00110000_10101000 : OUT <= 0;  //48 / 168 = 0
    16'b00110000_10101001 : OUT <= 0;  //48 / 169 = 0
    16'b00110000_10101010 : OUT <= 0;  //48 / 170 = 0
    16'b00110000_10101011 : OUT <= 0;  //48 / 171 = 0
    16'b00110000_10101100 : OUT <= 0;  //48 / 172 = 0
    16'b00110000_10101101 : OUT <= 0;  //48 / 173 = 0
    16'b00110000_10101110 : OUT <= 0;  //48 / 174 = 0
    16'b00110000_10101111 : OUT <= 0;  //48 / 175 = 0
    16'b00110000_10110000 : OUT <= 0;  //48 / 176 = 0
    16'b00110000_10110001 : OUT <= 0;  //48 / 177 = 0
    16'b00110000_10110010 : OUT <= 0;  //48 / 178 = 0
    16'b00110000_10110011 : OUT <= 0;  //48 / 179 = 0
    16'b00110000_10110100 : OUT <= 0;  //48 / 180 = 0
    16'b00110000_10110101 : OUT <= 0;  //48 / 181 = 0
    16'b00110000_10110110 : OUT <= 0;  //48 / 182 = 0
    16'b00110000_10110111 : OUT <= 0;  //48 / 183 = 0
    16'b00110000_10111000 : OUT <= 0;  //48 / 184 = 0
    16'b00110000_10111001 : OUT <= 0;  //48 / 185 = 0
    16'b00110000_10111010 : OUT <= 0;  //48 / 186 = 0
    16'b00110000_10111011 : OUT <= 0;  //48 / 187 = 0
    16'b00110000_10111100 : OUT <= 0;  //48 / 188 = 0
    16'b00110000_10111101 : OUT <= 0;  //48 / 189 = 0
    16'b00110000_10111110 : OUT <= 0;  //48 / 190 = 0
    16'b00110000_10111111 : OUT <= 0;  //48 / 191 = 0
    16'b00110000_11000000 : OUT <= 0;  //48 / 192 = 0
    16'b00110000_11000001 : OUT <= 0;  //48 / 193 = 0
    16'b00110000_11000010 : OUT <= 0;  //48 / 194 = 0
    16'b00110000_11000011 : OUT <= 0;  //48 / 195 = 0
    16'b00110000_11000100 : OUT <= 0;  //48 / 196 = 0
    16'b00110000_11000101 : OUT <= 0;  //48 / 197 = 0
    16'b00110000_11000110 : OUT <= 0;  //48 / 198 = 0
    16'b00110000_11000111 : OUT <= 0;  //48 / 199 = 0
    16'b00110000_11001000 : OUT <= 0;  //48 / 200 = 0
    16'b00110000_11001001 : OUT <= 0;  //48 / 201 = 0
    16'b00110000_11001010 : OUT <= 0;  //48 / 202 = 0
    16'b00110000_11001011 : OUT <= 0;  //48 / 203 = 0
    16'b00110000_11001100 : OUT <= 0;  //48 / 204 = 0
    16'b00110000_11001101 : OUT <= 0;  //48 / 205 = 0
    16'b00110000_11001110 : OUT <= 0;  //48 / 206 = 0
    16'b00110000_11001111 : OUT <= 0;  //48 / 207 = 0
    16'b00110000_11010000 : OUT <= 0;  //48 / 208 = 0
    16'b00110000_11010001 : OUT <= 0;  //48 / 209 = 0
    16'b00110000_11010010 : OUT <= 0;  //48 / 210 = 0
    16'b00110000_11010011 : OUT <= 0;  //48 / 211 = 0
    16'b00110000_11010100 : OUT <= 0;  //48 / 212 = 0
    16'b00110000_11010101 : OUT <= 0;  //48 / 213 = 0
    16'b00110000_11010110 : OUT <= 0;  //48 / 214 = 0
    16'b00110000_11010111 : OUT <= 0;  //48 / 215 = 0
    16'b00110000_11011000 : OUT <= 0;  //48 / 216 = 0
    16'b00110000_11011001 : OUT <= 0;  //48 / 217 = 0
    16'b00110000_11011010 : OUT <= 0;  //48 / 218 = 0
    16'b00110000_11011011 : OUT <= 0;  //48 / 219 = 0
    16'b00110000_11011100 : OUT <= 0;  //48 / 220 = 0
    16'b00110000_11011101 : OUT <= 0;  //48 / 221 = 0
    16'b00110000_11011110 : OUT <= 0;  //48 / 222 = 0
    16'b00110000_11011111 : OUT <= 0;  //48 / 223 = 0
    16'b00110000_11100000 : OUT <= 0;  //48 / 224 = 0
    16'b00110000_11100001 : OUT <= 0;  //48 / 225 = 0
    16'b00110000_11100010 : OUT <= 0;  //48 / 226 = 0
    16'b00110000_11100011 : OUT <= 0;  //48 / 227 = 0
    16'b00110000_11100100 : OUT <= 0;  //48 / 228 = 0
    16'b00110000_11100101 : OUT <= 0;  //48 / 229 = 0
    16'b00110000_11100110 : OUT <= 0;  //48 / 230 = 0
    16'b00110000_11100111 : OUT <= 0;  //48 / 231 = 0
    16'b00110000_11101000 : OUT <= 0;  //48 / 232 = 0
    16'b00110000_11101001 : OUT <= 0;  //48 / 233 = 0
    16'b00110000_11101010 : OUT <= 0;  //48 / 234 = 0
    16'b00110000_11101011 : OUT <= 0;  //48 / 235 = 0
    16'b00110000_11101100 : OUT <= 0;  //48 / 236 = 0
    16'b00110000_11101101 : OUT <= 0;  //48 / 237 = 0
    16'b00110000_11101110 : OUT <= 0;  //48 / 238 = 0
    16'b00110000_11101111 : OUT <= 0;  //48 / 239 = 0
    16'b00110000_11110000 : OUT <= 0;  //48 / 240 = 0
    16'b00110000_11110001 : OUT <= 0;  //48 / 241 = 0
    16'b00110000_11110010 : OUT <= 0;  //48 / 242 = 0
    16'b00110000_11110011 : OUT <= 0;  //48 / 243 = 0
    16'b00110000_11110100 : OUT <= 0;  //48 / 244 = 0
    16'b00110000_11110101 : OUT <= 0;  //48 / 245 = 0
    16'b00110000_11110110 : OUT <= 0;  //48 / 246 = 0
    16'b00110000_11110111 : OUT <= 0;  //48 / 247 = 0
    16'b00110000_11111000 : OUT <= 0;  //48 / 248 = 0
    16'b00110000_11111001 : OUT <= 0;  //48 / 249 = 0
    16'b00110000_11111010 : OUT <= 0;  //48 / 250 = 0
    16'b00110000_11111011 : OUT <= 0;  //48 / 251 = 0
    16'b00110000_11111100 : OUT <= 0;  //48 / 252 = 0
    16'b00110000_11111101 : OUT <= 0;  //48 / 253 = 0
    16'b00110000_11111110 : OUT <= 0;  //48 / 254 = 0
    16'b00110000_11111111 : OUT <= 0;  //48 / 255 = 0
    16'b00110001_00000000 : OUT <= 0;  //49 / 0 = 0
    16'b00110001_00000001 : OUT <= 49;  //49 / 1 = 49
    16'b00110001_00000010 : OUT <= 24;  //49 / 2 = 24
    16'b00110001_00000011 : OUT <= 16;  //49 / 3 = 16
    16'b00110001_00000100 : OUT <= 12;  //49 / 4 = 12
    16'b00110001_00000101 : OUT <= 9;  //49 / 5 = 9
    16'b00110001_00000110 : OUT <= 8;  //49 / 6 = 8
    16'b00110001_00000111 : OUT <= 7;  //49 / 7 = 7
    16'b00110001_00001000 : OUT <= 6;  //49 / 8 = 6
    16'b00110001_00001001 : OUT <= 5;  //49 / 9 = 5
    16'b00110001_00001010 : OUT <= 4;  //49 / 10 = 4
    16'b00110001_00001011 : OUT <= 4;  //49 / 11 = 4
    16'b00110001_00001100 : OUT <= 4;  //49 / 12 = 4
    16'b00110001_00001101 : OUT <= 3;  //49 / 13 = 3
    16'b00110001_00001110 : OUT <= 3;  //49 / 14 = 3
    16'b00110001_00001111 : OUT <= 3;  //49 / 15 = 3
    16'b00110001_00010000 : OUT <= 3;  //49 / 16 = 3
    16'b00110001_00010001 : OUT <= 2;  //49 / 17 = 2
    16'b00110001_00010010 : OUT <= 2;  //49 / 18 = 2
    16'b00110001_00010011 : OUT <= 2;  //49 / 19 = 2
    16'b00110001_00010100 : OUT <= 2;  //49 / 20 = 2
    16'b00110001_00010101 : OUT <= 2;  //49 / 21 = 2
    16'b00110001_00010110 : OUT <= 2;  //49 / 22 = 2
    16'b00110001_00010111 : OUT <= 2;  //49 / 23 = 2
    16'b00110001_00011000 : OUT <= 2;  //49 / 24 = 2
    16'b00110001_00011001 : OUT <= 1;  //49 / 25 = 1
    16'b00110001_00011010 : OUT <= 1;  //49 / 26 = 1
    16'b00110001_00011011 : OUT <= 1;  //49 / 27 = 1
    16'b00110001_00011100 : OUT <= 1;  //49 / 28 = 1
    16'b00110001_00011101 : OUT <= 1;  //49 / 29 = 1
    16'b00110001_00011110 : OUT <= 1;  //49 / 30 = 1
    16'b00110001_00011111 : OUT <= 1;  //49 / 31 = 1
    16'b00110001_00100000 : OUT <= 1;  //49 / 32 = 1
    16'b00110001_00100001 : OUT <= 1;  //49 / 33 = 1
    16'b00110001_00100010 : OUT <= 1;  //49 / 34 = 1
    16'b00110001_00100011 : OUT <= 1;  //49 / 35 = 1
    16'b00110001_00100100 : OUT <= 1;  //49 / 36 = 1
    16'b00110001_00100101 : OUT <= 1;  //49 / 37 = 1
    16'b00110001_00100110 : OUT <= 1;  //49 / 38 = 1
    16'b00110001_00100111 : OUT <= 1;  //49 / 39 = 1
    16'b00110001_00101000 : OUT <= 1;  //49 / 40 = 1
    16'b00110001_00101001 : OUT <= 1;  //49 / 41 = 1
    16'b00110001_00101010 : OUT <= 1;  //49 / 42 = 1
    16'b00110001_00101011 : OUT <= 1;  //49 / 43 = 1
    16'b00110001_00101100 : OUT <= 1;  //49 / 44 = 1
    16'b00110001_00101101 : OUT <= 1;  //49 / 45 = 1
    16'b00110001_00101110 : OUT <= 1;  //49 / 46 = 1
    16'b00110001_00101111 : OUT <= 1;  //49 / 47 = 1
    16'b00110001_00110000 : OUT <= 1;  //49 / 48 = 1
    16'b00110001_00110001 : OUT <= 1;  //49 / 49 = 1
    16'b00110001_00110010 : OUT <= 0;  //49 / 50 = 0
    16'b00110001_00110011 : OUT <= 0;  //49 / 51 = 0
    16'b00110001_00110100 : OUT <= 0;  //49 / 52 = 0
    16'b00110001_00110101 : OUT <= 0;  //49 / 53 = 0
    16'b00110001_00110110 : OUT <= 0;  //49 / 54 = 0
    16'b00110001_00110111 : OUT <= 0;  //49 / 55 = 0
    16'b00110001_00111000 : OUT <= 0;  //49 / 56 = 0
    16'b00110001_00111001 : OUT <= 0;  //49 / 57 = 0
    16'b00110001_00111010 : OUT <= 0;  //49 / 58 = 0
    16'b00110001_00111011 : OUT <= 0;  //49 / 59 = 0
    16'b00110001_00111100 : OUT <= 0;  //49 / 60 = 0
    16'b00110001_00111101 : OUT <= 0;  //49 / 61 = 0
    16'b00110001_00111110 : OUT <= 0;  //49 / 62 = 0
    16'b00110001_00111111 : OUT <= 0;  //49 / 63 = 0
    16'b00110001_01000000 : OUT <= 0;  //49 / 64 = 0
    16'b00110001_01000001 : OUT <= 0;  //49 / 65 = 0
    16'b00110001_01000010 : OUT <= 0;  //49 / 66 = 0
    16'b00110001_01000011 : OUT <= 0;  //49 / 67 = 0
    16'b00110001_01000100 : OUT <= 0;  //49 / 68 = 0
    16'b00110001_01000101 : OUT <= 0;  //49 / 69 = 0
    16'b00110001_01000110 : OUT <= 0;  //49 / 70 = 0
    16'b00110001_01000111 : OUT <= 0;  //49 / 71 = 0
    16'b00110001_01001000 : OUT <= 0;  //49 / 72 = 0
    16'b00110001_01001001 : OUT <= 0;  //49 / 73 = 0
    16'b00110001_01001010 : OUT <= 0;  //49 / 74 = 0
    16'b00110001_01001011 : OUT <= 0;  //49 / 75 = 0
    16'b00110001_01001100 : OUT <= 0;  //49 / 76 = 0
    16'b00110001_01001101 : OUT <= 0;  //49 / 77 = 0
    16'b00110001_01001110 : OUT <= 0;  //49 / 78 = 0
    16'b00110001_01001111 : OUT <= 0;  //49 / 79 = 0
    16'b00110001_01010000 : OUT <= 0;  //49 / 80 = 0
    16'b00110001_01010001 : OUT <= 0;  //49 / 81 = 0
    16'b00110001_01010010 : OUT <= 0;  //49 / 82 = 0
    16'b00110001_01010011 : OUT <= 0;  //49 / 83 = 0
    16'b00110001_01010100 : OUT <= 0;  //49 / 84 = 0
    16'b00110001_01010101 : OUT <= 0;  //49 / 85 = 0
    16'b00110001_01010110 : OUT <= 0;  //49 / 86 = 0
    16'b00110001_01010111 : OUT <= 0;  //49 / 87 = 0
    16'b00110001_01011000 : OUT <= 0;  //49 / 88 = 0
    16'b00110001_01011001 : OUT <= 0;  //49 / 89 = 0
    16'b00110001_01011010 : OUT <= 0;  //49 / 90 = 0
    16'b00110001_01011011 : OUT <= 0;  //49 / 91 = 0
    16'b00110001_01011100 : OUT <= 0;  //49 / 92 = 0
    16'b00110001_01011101 : OUT <= 0;  //49 / 93 = 0
    16'b00110001_01011110 : OUT <= 0;  //49 / 94 = 0
    16'b00110001_01011111 : OUT <= 0;  //49 / 95 = 0
    16'b00110001_01100000 : OUT <= 0;  //49 / 96 = 0
    16'b00110001_01100001 : OUT <= 0;  //49 / 97 = 0
    16'b00110001_01100010 : OUT <= 0;  //49 / 98 = 0
    16'b00110001_01100011 : OUT <= 0;  //49 / 99 = 0
    16'b00110001_01100100 : OUT <= 0;  //49 / 100 = 0
    16'b00110001_01100101 : OUT <= 0;  //49 / 101 = 0
    16'b00110001_01100110 : OUT <= 0;  //49 / 102 = 0
    16'b00110001_01100111 : OUT <= 0;  //49 / 103 = 0
    16'b00110001_01101000 : OUT <= 0;  //49 / 104 = 0
    16'b00110001_01101001 : OUT <= 0;  //49 / 105 = 0
    16'b00110001_01101010 : OUT <= 0;  //49 / 106 = 0
    16'b00110001_01101011 : OUT <= 0;  //49 / 107 = 0
    16'b00110001_01101100 : OUT <= 0;  //49 / 108 = 0
    16'b00110001_01101101 : OUT <= 0;  //49 / 109 = 0
    16'b00110001_01101110 : OUT <= 0;  //49 / 110 = 0
    16'b00110001_01101111 : OUT <= 0;  //49 / 111 = 0
    16'b00110001_01110000 : OUT <= 0;  //49 / 112 = 0
    16'b00110001_01110001 : OUT <= 0;  //49 / 113 = 0
    16'b00110001_01110010 : OUT <= 0;  //49 / 114 = 0
    16'b00110001_01110011 : OUT <= 0;  //49 / 115 = 0
    16'b00110001_01110100 : OUT <= 0;  //49 / 116 = 0
    16'b00110001_01110101 : OUT <= 0;  //49 / 117 = 0
    16'b00110001_01110110 : OUT <= 0;  //49 / 118 = 0
    16'b00110001_01110111 : OUT <= 0;  //49 / 119 = 0
    16'b00110001_01111000 : OUT <= 0;  //49 / 120 = 0
    16'b00110001_01111001 : OUT <= 0;  //49 / 121 = 0
    16'b00110001_01111010 : OUT <= 0;  //49 / 122 = 0
    16'b00110001_01111011 : OUT <= 0;  //49 / 123 = 0
    16'b00110001_01111100 : OUT <= 0;  //49 / 124 = 0
    16'b00110001_01111101 : OUT <= 0;  //49 / 125 = 0
    16'b00110001_01111110 : OUT <= 0;  //49 / 126 = 0
    16'b00110001_01111111 : OUT <= 0;  //49 / 127 = 0
    16'b00110001_10000000 : OUT <= 0;  //49 / 128 = 0
    16'b00110001_10000001 : OUT <= 0;  //49 / 129 = 0
    16'b00110001_10000010 : OUT <= 0;  //49 / 130 = 0
    16'b00110001_10000011 : OUT <= 0;  //49 / 131 = 0
    16'b00110001_10000100 : OUT <= 0;  //49 / 132 = 0
    16'b00110001_10000101 : OUT <= 0;  //49 / 133 = 0
    16'b00110001_10000110 : OUT <= 0;  //49 / 134 = 0
    16'b00110001_10000111 : OUT <= 0;  //49 / 135 = 0
    16'b00110001_10001000 : OUT <= 0;  //49 / 136 = 0
    16'b00110001_10001001 : OUT <= 0;  //49 / 137 = 0
    16'b00110001_10001010 : OUT <= 0;  //49 / 138 = 0
    16'b00110001_10001011 : OUT <= 0;  //49 / 139 = 0
    16'b00110001_10001100 : OUT <= 0;  //49 / 140 = 0
    16'b00110001_10001101 : OUT <= 0;  //49 / 141 = 0
    16'b00110001_10001110 : OUT <= 0;  //49 / 142 = 0
    16'b00110001_10001111 : OUT <= 0;  //49 / 143 = 0
    16'b00110001_10010000 : OUT <= 0;  //49 / 144 = 0
    16'b00110001_10010001 : OUT <= 0;  //49 / 145 = 0
    16'b00110001_10010010 : OUT <= 0;  //49 / 146 = 0
    16'b00110001_10010011 : OUT <= 0;  //49 / 147 = 0
    16'b00110001_10010100 : OUT <= 0;  //49 / 148 = 0
    16'b00110001_10010101 : OUT <= 0;  //49 / 149 = 0
    16'b00110001_10010110 : OUT <= 0;  //49 / 150 = 0
    16'b00110001_10010111 : OUT <= 0;  //49 / 151 = 0
    16'b00110001_10011000 : OUT <= 0;  //49 / 152 = 0
    16'b00110001_10011001 : OUT <= 0;  //49 / 153 = 0
    16'b00110001_10011010 : OUT <= 0;  //49 / 154 = 0
    16'b00110001_10011011 : OUT <= 0;  //49 / 155 = 0
    16'b00110001_10011100 : OUT <= 0;  //49 / 156 = 0
    16'b00110001_10011101 : OUT <= 0;  //49 / 157 = 0
    16'b00110001_10011110 : OUT <= 0;  //49 / 158 = 0
    16'b00110001_10011111 : OUT <= 0;  //49 / 159 = 0
    16'b00110001_10100000 : OUT <= 0;  //49 / 160 = 0
    16'b00110001_10100001 : OUT <= 0;  //49 / 161 = 0
    16'b00110001_10100010 : OUT <= 0;  //49 / 162 = 0
    16'b00110001_10100011 : OUT <= 0;  //49 / 163 = 0
    16'b00110001_10100100 : OUT <= 0;  //49 / 164 = 0
    16'b00110001_10100101 : OUT <= 0;  //49 / 165 = 0
    16'b00110001_10100110 : OUT <= 0;  //49 / 166 = 0
    16'b00110001_10100111 : OUT <= 0;  //49 / 167 = 0
    16'b00110001_10101000 : OUT <= 0;  //49 / 168 = 0
    16'b00110001_10101001 : OUT <= 0;  //49 / 169 = 0
    16'b00110001_10101010 : OUT <= 0;  //49 / 170 = 0
    16'b00110001_10101011 : OUT <= 0;  //49 / 171 = 0
    16'b00110001_10101100 : OUT <= 0;  //49 / 172 = 0
    16'b00110001_10101101 : OUT <= 0;  //49 / 173 = 0
    16'b00110001_10101110 : OUT <= 0;  //49 / 174 = 0
    16'b00110001_10101111 : OUT <= 0;  //49 / 175 = 0
    16'b00110001_10110000 : OUT <= 0;  //49 / 176 = 0
    16'b00110001_10110001 : OUT <= 0;  //49 / 177 = 0
    16'b00110001_10110010 : OUT <= 0;  //49 / 178 = 0
    16'b00110001_10110011 : OUT <= 0;  //49 / 179 = 0
    16'b00110001_10110100 : OUT <= 0;  //49 / 180 = 0
    16'b00110001_10110101 : OUT <= 0;  //49 / 181 = 0
    16'b00110001_10110110 : OUT <= 0;  //49 / 182 = 0
    16'b00110001_10110111 : OUT <= 0;  //49 / 183 = 0
    16'b00110001_10111000 : OUT <= 0;  //49 / 184 = 0
    16'b00110001_10111001 : OUT <= 0;  //49 / 185 = 0
    16'b00110001_10111010 : OUT <= 0;  //49 / 186 = 0
    16'b00110001_10111011 : OUT <= 0;  //49 / 187 = 0
    16'b00110001_10111100 : OUT <= 0;  //49 / 188 = 0
    16'b00110001_10111101 : OUT <= 0;  //49 / 189 = 0
    16'b00110001_10111110 : OUT <= 0;  //49 / 190 = 0
    16'b00110001_10111111 : OUT <= 0;  //49 / 191 = 0
    16'b00110001_11000000 : OUT <= 0;  //49 / 192 = 0
    16'b00110001_11000001 : OUT <= 0;  //49 / 193 = 0
    16'b00110001_11000010 : OUT <= 0;  //49 / 194 = 0
    16'b00110001_11000011 : OUT <= 0;  //49 / 195 = 0
    16'b00110001_11000100 : OUT <= 0;  //49 / 196 = 0
    16'b00110001_11000101 : OUT <= 0;  //49 / 197 = 0
    16'b00110001_11000110 : OUT <= 0;  //49 / 198 = 0
    16'b00110001_11000111 : OUT <= 0;  //49 / 199 = 0
    16'b00110001_11001000 : OUT <= 0;  //49 / 200 = 0
    16'b00110001_11001001 : OUT <= 0;  //49 / 201 = 0
    16'b00110001_11001010 : OUT <= 0;  //49 / 202 = 0
    16'b00110001_11001011 : OUT <= 0;  //49 / 203 = 0
    16'b00110001_11001100 : OUT <= 0;  //49 / 204 = 0
    16'b00110001_11001101 : OUT <= 0;  //49 / 205 = 0
    16'b00110001_11001110 : OUT <= 0;  //49 / 206 = 0
    16'b00110001_11001111 : OUT <= 0;  //49 / 207 = 0
    16'b00110001_11010000 : OUT <= 0;  //49 / 208 = 0
    16'b00110001_11010001 : OUT <= 0;  //49 / 209 = 0
    16'b00110001_11010010 : OUT <= 0;  //49 / 210 = 0
    16'b00110001_11010011 : OUT <= 0;  //49 / 211 = 0
    16'b00110001_11010100 : OUT <= 0;  //49 / 212 = 0
    16'b00110001_11010101 : OUT <= 0;  //49 / 213 = 0
    16'b00110001_11010110 : OUT <= 0;  //49 / 214 = 0
    16'b00110001_11010111 : OUT <= 0;  //49 / 215 = 0
    16'b00110001_11011000 : OUT <= 0;  //49 / 216 = 0
    16'b00110001_11011001 : OUT <= 0;  //49 / 217 = 0
    16'b00110001_11011010 : OUT <= 0;  //49 / 218 = 0
    16'b00110001_11011011 : OUT <= 0;  //49 / 219 = 0
    16'b00110001_11011100 : OUT <= 0;  //49 / 220 = 0
    16'b00110001_11011101 : OUT <= 0;  //49 / 221 = 0
    16'b00110001_11011110 : OUT <= 0;  //49 / 222 = 0
    16'b00110001_11011111 : OUT <= 0;  //49 / 223 = 0
    16'b00110001_11100000 : OUT <= 0;  //49 / 224 = 0
    16'b00110001_11100001 : OUT <= 0;  //49 / 225 = 0
    16'b00110001_11100010 : OUT <= 0;  //49 / 226 = 0
    16'b00110001_11100011 : OUT <= 0;  //49 / 227 = 0
    16'b00110001_11100100 : OUT <= 0;  //49 / 228 = 0
    16'b00110001_11100101 : OUT <= 0;  //49 / 229 = 0
    16'b00110001_11100110 : OUT <= 0;  //49 / 230 = 0
    16'b00110001_11100111 : OUT <= 0;  //49 / 231 = 0
    16'b00110001_11101000 : OUT <= 0;  //49 / 232 = 0
    16'b00110001_11101001 : OUT <= 0;  //49 / 233 = 0
    16'b00110001_11101010 : OUT <= 0;  //49 / 234 = 0
    16'b00110001_11101011 : OUT <= 0;  //49 / 235 = 0
    16'b00110001_11101100 : OUT <= 0;  //49 / 236 = 0
    16'b00110001_11101101 : OUT <= 0;  //49 / 237 = 0
    16'b00110001_11101110 : OUT <= 0;  //49 / 238 = 0
    16'b00110001_11101111 : OUT <= 0;  //49 / 239 = 0
    16'b00110001_11110000 : OUT <= 0;  //49 / 240 = 0
    16'b00110001_11110001 : OUT <= 0;  //49 / 241 = 0
    16'b00110001_11110010 : OUT <= 0;  //49 / 242 = 0
    16'b00110001_11110011 : OUT <= 0;  //49 / 243 = 0
    16'b00110001_11110100 : OUT <= 0;  //49 / 244 = 0
    16'b00110001_11110101 : OUT <= 0;  //49 / 245 = 0
    16'b00110001_11110110 : OUT <= 0;  //49 / 246 = 0
    16'b00110001_11110111 : OUT <= 0;  //49 / 247 = 0
    16'b00110001_11111000 : OUT <= 0;  //49 / 248 = 0
    16'b00110001_11111001 : OUT <= 0;  //49 / 249 = 0
    16'b00110001_11111010 : OUT <= 0;  //49 / 250 = 0
    16'b00110001_11111011 : OUT <= 0;  //49 / 251 = 0
    16'b00110001_11111100 : OUT <= 0;  //49 / 252 = 0
    16'b00110001_11111101 : OUT <= 0;  //49 / 253 = 0
    16'b00110001_11111110 : OUT <= 0;  //49 / 254 = 0
    16'b00110001_11111111 : OUT <= 0;  //49 / 255 = 0
    16'b00110010_00000000 : OUT <= 0;  //50 / 0 = 0
    16'b00110010_00000001 : OUT <= 50;  //50 / 1 = 50
    16'b00110010_00000010 : OUT <= 25;  //50 / 2 = 25
    16'b00110010_00000011 : OUT <= 16;  //50 / 3 = 16
    16'b00110010_00000100 : OUT <= 12;  //50 / 4 = 12
    16'b00110010_00000101 : OUT <= 10;  //50 / 5 = 10
    16'b00110010_00000110 : OUT <= 8;  //50 / 6 = 8
    16'b00110010_00000111 : OUT <= 7;  //50 / 7 = 7
    16'b00110010_00001000 : OUT <= 6;  //50 / 8 = 6
    16'b00110010_00001001 : OUT <= 5;  //50 / 9 = 5
    16'b00110010_00001010 : OUT <= 5;  //50 / 10 = 5
    16'b00110010_00001011 : OUT <= 4;  //50 / 11 = 4
    16'b00110010_00001100 : OUT <= 4;  //50 / 12 = 4
    16'b00110010_00001101 : OUT <= 3;  //50 / 13 = 3
    16'b00110010_00001110 : OUT <= 3;  //50 / 14 = 3
    16'b00110010_00001111 : OUT <= 3;  //50 / 15 = 3
    16'b00110010_00010000 : OUT <= 3;  //50 / 16 = 3
    16'b00110010_00010001 : OUT <= 2;  //50 / 17 = 2
    16'b00110010_00010010 : OUT <= 2;  //50 / 18 = 2
    16'b00110010_00010011 : OUT <= 2;  //50 / 19 = 2
    16'b00110010_00010100 : OUT <= 2;  //50 / 20 = 2
    16'b00110010_00010101 : OUT <= 2;  //50 / 21 = 2
    16'b00110010_00010110 : OUT <= 2;  //50 / 22 = 2
    16'b00110010_00010111 : OUT <= 2;  //50 / 23 = 2
    16'b00110010_00011000 : OUT <= 2;  //50 / 24 = 2
    16'b00110010_00011001 : OUT <= 2;  //50 / 25 = 2
    16'b00110010_00011010 : OUT <= 1;  //50 / 26 = 1
    16'b00110010_00011011 : OUT <= 1;  //50 / 27 = 1
    16'b00110010_00011100 : OUT <= 1;  //50 / 28 = 1
    16'b00110010_00011101 : OUT <= 1;  //50 / 29 = 1
    16'b00110010_00011110 : OUT <= 1;  //50 / 30 = 1
    16'b00110010_00011111 : OUT <= 1;  //50 / 31 = 1
    16'b00110010_00100000 : OUT <= 1;  //50 / 32 = 1
    16'b00110010_00100001 : OUT <= 1;  //50 / 33 = 1
    16'b00110010_00100010 : OUT <= 1;  //50 / 34 = 1
    16'b00110010_00100011 : OUT <= 1;  //50 / 35 = 1
    16'b00110010_00100100 : OUT <= 1;  //50 / 36 = 1
    16'b00110010_00100101 : OUT <= 1;  //50 / 37 = 1
    16'b00110010_00100110 : OUT <= 1;  //50 / 38 = 1
    16'b00110010_00100111 : OUT <= 1;  //50 / 39 = 1
    16'b00110010_00101000 : OUT <= 1;  //50 / 40 = 1
    16'b00110010_00101001 : OUT <= 1;  //50 / 41 = 1
    16'b00110010_00101010 : OUT <= 1;  //50 / 42 = 1
    16'b00110010_00101011 : OUT <= 1;  //50 / 43 = 1
    16'b00110010_00101100 : OUT <= 1;  //50 / 44 = 1
    16'b00110010_00101101 : OUT <= 1;  //50 / 45 = 1
    16'b00110010_00101110 : OUT <= 1;  //50 / 46 = 1
    16'b00110010_00101111 : OUT <= 1;  //50 / 47 = 1
    16'b00110010_00110000 : OUT <= 1;  //50 / 48 = 1
    16'b00110010_00110001 : OUT <= 1;  //50 / 49 = 1
    16'b00110010_00110010 : OUT <= 1;  //50 / 50 = 1
    16'b00110010_00110011 : OUT <= 0;  //50 / 51 = 0
    16'b00110010_00110100 : OUT <= 0;  //50 / 52 = 0
    16'b00110010_00110101 : OUT <= 0;  //50 / 53 = 0
    16'b00110010_00110110 : OUT <= 0;  //50 / 54 = 0
    16'b00110010_00110111 : OUT <= 0;  //50 / 55 = 0
    16'b00110010_00111000 : OUT <= 0;  //50 / 56 = 0
    16'b00110010_00111001 : OUT <= 0;  //50 / 57 = 0
    16'b00110010_00111010 : OUT <= 0;  //50 / 58 = 0
    16'b00110010_00111011 : OUT <= 0;  //50 / 59 = 0
    16'b00110010_00111100 : OUT <= 0;  //50 / 60 = 0
    16'b00110010_00111101 : OUT <= 0;  //50 / 61 = 0
    16'b00110010_00111110 : OUT <= 0;  //50 / 62 = 0
    16'b00110010_00111111 : OUT <= 0;  //50 / 63 = 0
    16'b00110010_01000000 : OUT <= 0;  //50 / 64 = 0
    16'b00110010_01000001 : OUT <= 0;  //50 / 65 = 0
    16'b00110010_01000010 : OUT <= 0;  //50 / 66 = 0
    16'b00110010_01000011 : OUT <= 0;  //50 / 67 = 0
    16'b00110010_01000100 : OUT <= 0;  //50 / 68 = 0
    16'b00110010_01000101 : OUT <= 0;  //50 / 69 = 0
    16'b00110010_01000110 : OUT <= 0;  //50 / 70 = 0
    16'b00110010_01000111 : OUT <= 0;  //50 / 71 = 0
    16'b00110010_01001000 : OUT <= 0;  //50 / 72 = 0
    16'b00110010_01001001 : OUT <= 0;  //50 / 73 = 0
    16'b00110010_01001010 : OUT <= 0;  //50 / 74 = 0
    16'b00110010_01001011 : OUT <= 0;  //50 / 75 = 0
    16'b00110010_01001100 : OUT <= 0;  //50 / 76 = 0
    16'b00110010_01001101 : OUT <= 0;  //50 / 77 = 0
    16'b00110010_01001110 : OUT <= 0;  //50 / 78 = 0
    16'b00110010_01001111 : OUT <= 0;  //50 / 79 = 0
    16'b00110010_01010000 : OUT <= 0;  //50 / 80 = 0
    16'b00110010_01010001 : OUT <= 0;  //50 / 81 = 0
    16'b00110010_01010010 : OUT <= 0;  //50 / 82 = 0
    16'b00110010_01010011 : OUT <= 0;  //50 / 83 = 0
    16'b00110010_01010100 : OUT <= 0;  //50 / 84 = 0
    16'b00110010_01010101 : OUT <= 0;  //50 / 85 = 0
    16'b00110010_01010110 : OUT <= 0;  //50 / 86 = 0
    16'b00110010_01010111 : OUT <= 0;  //50 / 87 = 0
    16'b00110010_01011000 : OUT <= 0;  //50 / 88 = 0
    16'b00110010_01011001 : OUT <= 0;  //50 / 89 = 0
    16'b00110010_01011010 : OUT <= 0;  //50 / 90 = 0
    16'b00110010_01011011 : OUT <= 0;  //50 / 91 = 0
    16'b00110010_01011100 : OUT <= 0;  //50 / 92 = 0
    16'b00110010_01011101 : OUT <= 0;  //50 / 93 = 0
    16'b00110010_01011110 : OUT <= 0;  //50 / 94 = 0
    16'b00110010_01011111 : OUT <= 0;  //50 / 95 = 0
    16'b00110010_01100000 : OUT <= 0;  //50 / 96 = 0
    16'b00110010_01100001 : OUT <= 0;  //50 / 97 = 0
    16'b00110010_01100010 : OUT <= 0;  //50 / 98 = 0
    16'b00110010_01100011 : OUT <= 0;  //50 / 99 = 0
    16'b00110010_01100100 : OUT <= 0;  //50 / 100 = 0
    16'b00110010_01100101 : OUT <= 0;  //50 / 101 = 0
    16'b00110010_01100110 : OUT <= 0;  //50 / 102 = 0
    16'b00110010_01100111 : OUT <= 0;  //50 / 103 = 0
    16'b00110010_01101000 : OUT <= 0;  //50 / 104 = 0
    16'b00110010_01101001 : OUT <= 0;  //50 / 105 = 0
    16'b00110010_01101010 : OUT <= 0;  //50 / 106 = 0
    16'b00110010_01101011 : OUT <= 0;  //50 / 107 = 0
    16'b00110010_01101100 : OUT <= 0;  //50 / 108 = 0
    16'b00110010_01101101 : OUT <= 0;  //50 / 109 = 0
    16'b00110010_01101110 : OUT <= 0;  //50 / 110 = 0
    16'b00110010_01101111 : OUT <= 0;  //50 / 111 = 0
    16'b00110010_01110000 : OUT <= 0;  //50 / 112 = 0
    16'b00110010_01110001 : OUT <= 0;  //50 / 113 = 0
    16'b00110010_01110010 : OUT <= 0;  //50 / 114 = 0
    16'b00110010_01110011 : OUT <= 0;  //50 / 115 = 0
    16'b00110010_01110100 : OUT <= 0;  //50 / 116 = 0
    16'b00110010_01110101 : OUT <= 0;  //50 / 117 = 0
    16'b00110010_01110110 : OUT <= 0;  //50 / 118 = 0
    16'b00110010_01110111 : OUT <= 0;  //50 / 119 = 0
    16'b00110010_01111000 : OUT <= 0;  //50 / 120 = 0
    16'b00110010_01111001 : OUT <= 0;  //50 / 121 = 0
    16'b00110010_01111010 : OUT <= 0;  //50 / 122 = 0
    16'b00110010_01111011 : OUT <= 0;  //50 / 123 = 0
    16'b00110010_01111100 : OUT <= 0;  //50 / 124 = 0
    16'b00110010_01111101 : OUT <= 0;  //50 / 125 = 0
    16'b00110010_01111110 : OUT <= 0;  //50 / 126 = 0
    16'b00110010_01111111 : OUT <= 0;  //50 / 127 = 0
    16'b00110010_10000000 : OUT <= 0;  //50 / 128 = 0
    16'b00110010_10000001 : OUT <= 0;  //50 / 129 = 0
    16'b00110010_10000010 : OUT <= 0;  //50 / 130 = 0
    16'b00110010_10000011 : OUT <= 0;  //50 / 131 = 0
    16'b00110010_10000100 : OUT <= 0;  //50 / 132 = 0
    16'b00110010_10000101 : OUT <= 0;  //50 / 133 = 0
    16'b00110010_10000110 : OUT <= 0;  //50 / 134 = 0
    16'b00110010_10000111 : OUT <= 0;  //50 / 135 = 0
    16'b00110010_10001000 : OUT <= 0;  //50 / 136 = 0
    16'b00110010_10001001 : OUT <= 0;  //50 / 137 = 0
    16'b00110010_10001010 : OUT <= 0;  //50 / 138 = 0
    16'b00110010_10001011 : OUT <= 0;  //50 / 139 = 0
    16'b00110010_10001100 : OUT <= 0;  //50 / 140 = 0
    16'b00110010_10001101 : OUT <= 0;  //50 / 141 = 0
    16'b00110010_10001110 : OUT <= 0;  //50 / 142 = 0
    16'b00110010_10001111 : OUT <= 0;  //50 / 143 = 0
    16'b00110010_10010000 : OUT <= 0;  //50 / 144 = 0
    16'b00110010_10010001 : OUT <= 0;  //50 / 145 = 0
    16'b00110010_10010010 : OUT <= 0;  //50 / 146 = 0
    16'b00110010_10010011 : OUT <= 0;  //50 / 147 = 0
    16'b00110010_10010100 : OUT <= 0;  //50 / 148 = 0
    16'b00110010_10010101 : OUT <= 0;  //50 / 149 = 0
    16'b00110010_10010110 : OUT <= 0;  //50 / 150 = 0
    16'b00110010_10010111 : OUT <= 0;  //50 / 151 = 0
    16'b00110010_10011000 : OUT <= 0;  //50 / 152 = 0
    16'b00110010_10011001 : OUT <= 0;  //50 / 153 = 0
    16'b00110010_10011010 : OUT <= 0;  //50 / 154 = 0
    16'b00110010_10011011 : OUT <= 0;  //50 / 155 = 0
    16'b00110010_10011100 : OUT <= 0;  //50 / 156 = 0
    16'b00110010_10011101 : OUT <= 0;  //50 / 157 = 0
    16'b00110010_10011110 : OUT <= 0;  //50 / 158 = 0
    16'b00110010_10011111 : OUT <= 0;  //50 / 159 = 0
    16'b00110010_10100000 : OUT <= 0;  //50 / 160 = 0
    16'b00110010_10100001 : OUT <= 0;  //50 / 161 = 0
    16'b00110010_10100010 : OUT <= 0;  //50 / 162 = 0
    16'b00110010_10100011 : OUT <= 0;  //50 / 163 = 0
    16'b00110010_10100100 : OUT <= 0;  //50 / 164 = 0
    16'b00110010_10100101 : OUT <= 0;  //50 / 165 = 0
    16'b00110010_10100110 : OUT <= 0;  //50 / 166 = 0
    16'b00110010_10100111 : OUT <= 0;  //50 / 167 = 0
    16'b00110010_10101000 : OUT <= 0;  //50 / 168 = 0
    16'b00110010_10101001 : OUT <= 0;  //50 / 169 = 0
    16'b00110010_10101010 : OUT <= 0;  //50 / 170 = 0
    16'b00110010_10101011 : OUT <= 0;  //50 / 171 = 0
    16'b00110010_10101100 : OUT <= 0;  //50 / 172 = 0
    16'b00110010_10101101 : OUT <= 0;  //50 / 173 = 0
    16'b00110010_10101110 : OUT <= 0;  //50 / 174 = 0
    16'b00110010_10101111 : OUT <= 0;  //50 / 175 = 0
    16'b00110010_10110000 : OUT <= 0;  //50 / 176 = 0
    16'b00110010_10110001 : OUT <= 0;  //50 / 177 = 0
    16'b00110010_10110010 : OUT <= 0;  //50 / 178 = 0
    16'b00110010_10110011 : OUT <= 0;  //50 / 179 = 0
    16'b00110010_10110100 : OUT <= 0;  //50 / 180 = 0
    16'b00110010_10110101 : OUT <= 0;  //50 / 181 = 0
    16'b00110010_10110110 : OUT <= 0;  //50 / 182 = 0
    16'b00110010_10110111 : OUT <= 0;  //50 / 183 = 0
    16'b00110010_10111000 : OUT <= 0;  //50 / 184 = 0
    16'b00110010_10111001 : OUT <= 0;  //50 / 185 = 0
    16'b00110010_10111010 : OUT <= 0;  //50 / 186 = 0
    16'b00110010_10111011 : OUT <= 0;  //50 / 187 = 0
    16'b00110010_10111100 : OUT <= 0;  //50 / 188 = 0
    16'b00110010_10111101 : OUT <= 0;  //50 / 189 = 0
    16'b00110010_10111110 : OUT <= 0;  //50 / 190 = 0
    16'b00110010_10111111 : OUT <= 0;  //50 / 191 = 0
    16'b00110010_11000000 : OUT <= 0;  //50 / 192 = 0
    16'b00110010_11000001 : OUT <= 0;  //50 / 193 = 0
    16'b00110010_11000010 : OUT <= 0;  //50 / 194 = 0
    16'b00110010_11000011 : OUT <= 0;  //50 / 195 = 0
    16'b00110010_11000100 : OUT <= 0;  //50 / 196 = 0
    16'b00110010_11000101 : OUT <= 0;  //50 / 197 = 0
    16'b00110010_11000110 : OUT <= 0;  //50 / 198 = 0
    16'b00110010_11000111 : OUT <= 0;  //50 / 199 = 0
    16'b00110010_11001000 : OUT <= 0;  //50 / 200 = 0
    16'b00110010_11001001 : OUT <= 0;  //50 / 201 = 0
    16'b00110010_11001010 : OUT <= 0;  //50 / 202 = 0
    16'b00110010_11001011 : OUT <= 0;  //50 / 203 = 0
    16'b00110010_11001100 : OUT <= 0;  //50 / 204 = 0
    16'b00110010_11001101 : OUT <= 0;  //50 / 205 = 0
    16'b00110010_11001110 : OUT <= 0;  //50 / 206 = 0
    16'b00110010_11001111 : OUT <= 0;  //50 / 207 = 0
    16'b00110010_11010000 : OUT <= 0;  //50 / 208 = 0
    16'b00110010_11010001 : OUT <= 0;  //50 / 209 = 0
    16'b00110010_11010010 : OUT <= 0;  //50 / 210 = 0
    16'b00110010_11010011 : OUT <= 0;  //50 / 211 = 0
    16'b00110010_11010100 : OUT <= 0;  //50 / 212 = 0
    16'b00110010_11010101 : OUT <= 0;  //50 / 213 = 0
    16'b00110010_11010110 : OUT <= 0;  //50 / 214 = 0
    16'b00110010_11010111 : OUT <= 0;  //50 / 215 = 0
    16'b00110010_11011000 : OUT <= 0;  //50 / 216 = 0
    16'b00110010_11011001 : OUT <= 0;  //50 / 217 = 0
    16'b00110010_11011010 : OUT <= 0;  //50 / 218 = 0
    16'b00110010_11011011 : OUT <= 0;  //50 / 219 = 0
    16'b00110010_11011100 : OUT <= 0;  //50 / 220 = 0
    16'b00110010_11011101 : OUT <= 0;  //50 / 221 = 0
    16'b00110010_11011110 : OUT <= 0;  //50 / 222 = 0
    16'b00110010_11011111 : OUT <= 0;  //50 / 223 = 0
    16'b00110010_11100000 : OUT <= 0;  //50 / 224 = 0
    16'b00110010_11100001 : OUT <= 0;  //50 / 225 = 0
    16'b00110010_11100010 : OUT <= 0;  //50 / 226 = 0
    16'b00110010_11100011 : OUT <= 0;  //50 / 227 = 0
    16'b00110010_11100100 : OUT <= 0;  //50 / 228 = 0
    16'b00110010_11100101 : OUT <= 0;  //50 / 229 = 0
    16'b00110010_11100110 : OUT <= 0;  //50 / 230 = 0
    16'b00110010_11100111 : OUT <= 0;  //50 / 231 = 0
    16'b00110010_11101000 : OUT <= 0;  //50 / 232 = 0
    16'b00110010_11101001 : OUT <= 0;  //50 / 233 = 0
    16'b00110010_11101010 : OUT <= 0;  //50 / 234 = 0
    16'b00110010_11101011 : OUT <= 0;  //50 / 235 = 0
    16'b00110010_11101100 : OUT <= 0;  //50 / 236 = 0
    16'b00110010_11101101 : OUT <= 0;  //50 / 237 = 0
    16'b00110010_11101110 : OUT <= 0;  //50 / 238 = 0
    16'b00110010_11101111 : OUT <= 0;  //50 / 239 = 0
    16'b00110010_11110000 : OUT <= 0;  //50 / 240 = 0
    16'b00110010_11110001 : OUT <= 0;  //50 / 241 = 0
    16'b00110010_11110010 : OUT <= 0;  //50 / 242 = 0
    16'b00110010_11110011 : OUT <= 0;  //50 / 243 = 0
    16'b00110010_11110100 : OUT <= 0;  //50 / 244 = 0
    16'b00110010_11110101 : OUT <= 0;  //50 / 245 = 0
    16'b00110010_11110110 : OUT <= 0;  //50 / 246 = 0
    16'b00110010_11110111 : OUT <= 0;  //50 / 247 = 0
    16'b00110010_11111000 : OUT <= 0;  //50 / 248 = 0
    16'b00110010_11111001 : OUT <= 0;  //50 / 249 = 0
    16'b00110010_11111010 : OUT <= 0;  //50 / 250 = 0
    16'b00110010_11111011 : OUT <= 0;  //50 / 251 = 0
    16'b00110010_11111100 : OUT <= 0;  //50 / 252 = 0
    16'b00110010_11111101 : OUT <= 0;  //50 / 253 = 0
    16'b00110010_11111110 : OUT <= 0;  //50 / 254 = 0
    16'b00110010_11111111 : OUT <= 0;  //50 / 255 = 0
    16'b00110011_00000000 : OUT <= 0;  //51 / 0 = 0
    16'b00110011_00000001 : OUT <= 51;  //51 / 1 = 51
    16'b00110011_00000010 : OUT <= 25;  //51 / 2 = 25
    16'b00110011_00000011 : OUT <= 17;  //51 / 3 = 17
    16'b00110011_00000100 : OUT <= 12;  //51 / 4 = 12
    16'b00110011_00000101 : OUT <= 10;  //51 / 5 = 10
    16'b00110011_00000110 : OUT <= 8;  //51 / 6 = 8
    16'b00110011_00000111 : OUT <= 7;  //51 / 7 = 7
    16'b00110011_00001000 : OUT <= 6;  //51 / 8 = 6
    16'b00110011_00001001 : OUT <= 5;  //51 / 9 = 5
    16'b00110011_00001010 : OUT <= 5;  //51 / 10 = 5
    16'b00110011_00001011 : OUT <= 4;  //51 / 11 = 4
    16'b00110011_00001100 : OUT <= 4;  //51 / 12 = 4
    16'b00110011_00001101 : OUT <= 3;  //51 / 13 = 3
    16'b00110011_00001110 : OUT <= 3;  //51 / 14 = 3
    16'b00110011_00001111 : OUT <= 3;  //51 / 15 = 3
    16'b00110011_00010000 : OUT <= 3;  //51 / 16 = 3
    16'b00110011_00010001 : OUT <= 3;  //51 / 17 = 3
    16'b00110011_00010010 : OUT <= 2;  //51 / 18 = 2
    16'b00110011_00010011 : OUT <= 2;  //51 / 19 = 2
    16'b00110011_00010100 : OUT <= 2;  //51 / 20 = 2
    16'b00110011_00010101 : OUT <= 2;  //51 / 21 = 2
    16'b00110011_00010110 : OUT <= 2;  //51 / 22 = 2
    16'b00110011_00010111 : OUT <= 2;  //51 / 23 = 2
    16'b00110011_00011000 : OUT <= 2;  //51 / 24 = 2
    16'b00110011_00011001 : OUT <= 2;  //51 / 25 = 2
    16'b00110011_00011010 : OUT <= 1;  //51 / 26 = 1
    16'b00110011_00011011 : OUT <= 1;  //51 / 27 = 1
    16'b00110011_00011100 : OUT <= 1;  //51 / 28 = 1
    16'b00110011_00011101 : OUT <= 1;  //51 / 29 = 1
    16'b00110011_00011110 : OUT <= 1;  //51 / 30 = 1
    16'b00110011_00011111 : OUT <= 1;  //51 / 31 = 1
    16'b00110011_00100000 : OUT <= 1;  //51 / 32 = 1
    16'b00110011_00100001 : OUT <= 1;  //51 / 33 = 1
    16'b00110011_00100010 : OUT <= 1;  //51 / 34 = 1
    16'b00110011_00100011 : OUT <= 1;  //51 / 35 = 1
    16'b00110011_00100100 : OUT <= 1;  //51 / 36 = 1
    16'b00110011_00100101 : OUT <= 1;  //51 / 37 = 1
    16'b00110011_00100110 : OUT <= 1;  //51 / 38 = 1
    16'b00110011_00100111 : OUT <= 1;  //51 / 39 = 1
    16'b00110011_00101000 : OUT <= 1;  //51 / 40 = 1
    16'b00110011_00101001 : OUT <= 1;  //51 / 41 = 1
    16'b00110011_00101010 : OUT <= 1;  //51 / 42 = 1
    16'b00110011_00101011 : OUT <= 1;  //51 / 43 = 1
    16'b00110011_00101100 : OUT <= 1;  //51 / 44 = 1
    16'b00110011_00101101 : OUT <= 1;  //51 / 45 = 1
    16'b00110011_00101110 : OUT <= 1;  //51 / 46 = 1
    16'b00110011_00101111 : OUT <= 1;  //51 / 47 = 1
    16'b00110011_00110000 : OUT <= 1;  //51 / 48 = 1
    16'b00110011_00110001 : OUT <= 1;  //51 / 49 = 1
    16'b00110011_00110010 : OUT <= 1;  //51 / 50 = 1
    16'b00110011_00110011 : OUT <= 1;  //51 / 51 = 1
    16'b00110011_00110100 : OUT <= 0;  //51 / 52 = 0
    16'b00110011_00110101 : OUT <= 0;  //51 / 53 = 0
    16'b00110011_00110110 : OUT <= 0;  //51 / 54 = 0
    16'b00110011_00110111 : OUT <= 0;  //51 / 55 = 0
    16'b00110011_00111000 : OUT <= 0;  //51 / 56 = 0
    16'b00110011_00111001 : OUT <= 0;  //51 / 57 = 0
    16'b00110011_00111010 : OUT <= 0;  //51 / 58 = 0
    16'b00110011_00111011 : OUT <= 0;  //51 / 59 = 0
    16'b00110011_00111100 : OUT <= 0;  //51 / 60 = 0
    16'b00110011_00111101 : OUT <= 0;  //51 / 61 = 0
    16'b00110011_00111110 : OUT <= 0;  //51 / 62 = 0
    16'b00110011_00111111 : OUT <= 0;  //51 / 63 = 0
    16'b00110011_01000000 : OUT <= 0;  //51 / 64 = 0
    16'b00110011_01000001 : OUT <= 0;  //51 / 65 = 0
    16'b00110011_01000010 : OUT <= 0;  //51 / 66 = 0
    16'b00110011_01000011 : OUT <= 0;  //51 / 67 = 0
    16'b00110011_01000100 : OUT <= 0;  //51 / 68 = 0
    16'b00110011_01000101 : OUT <= 0;  //51 / 69 = 0
    16'b00110011_01000110 : OUT <= 0;  //51 / 70 = 0
    16'b00110011_01000111 : OUT <= 0;  //51 / 71 = 0
    16'b00110011_01001000 : OUT <= 0;  //51 / 72 = 0
    16'b00110011_01001001 : OUT <= 0;  //51 / 73 = 0
    16'b00110011_01001010 : OUT <= 0;  //51 / 74 = 0
    16'b00110011_01001011 : OUT <= 0;  //51 / 75 = 0
    16'b00110011_01001100 : OUT <= 0;  //51 / 76 = 0
    16'b00110011_01001101 : OUT <= 0;  //51 / 77 = 0
    16'b00110011_01001110 : OUT <= 0;  //51 / 78 = 0
    16'b00110011_01001111 : OUT <= 0;  //51 / 79 = 0
    16'b00110011_01010000 : OUT <= 0;  //51 / 80 = 0
    16'b00110011_01010001 : OUT <= 0;  //51 / 81 = 0
    16'b00110011_01010010 : OUT <= 0;  //51 / 82 = 0
    16'b00110011_01010011 : OUT <= 0;  //51 / 83 = 0
    16'b00110011_01010100 : OUT <= 0;  //51 / 84 = 0
    16'b00110011_01010101 : OUT <= 0;  //51 / 85 = 0
    16'b00110011_01010110 : OUT <= 0;  //51 / 86 = 0
    16'b00110011_01010111 : OUT <= 0;  //51 / 87 = 0
    16'b00110011_01011000 : OUT <= 0;  //51 / 88 = 0
    16'b00110011_01011001 : OUT <= 0;  //51 / 89 = 0
    16'b00110011_01011010 : OUT <= 0;  //51 / 90 = 0
    16'b00110011_01011011 : OUT <= 0;  //51 / 91 = 0
    16'b00110011_01011100 : OUT <= 0;  //51 / 92 = 0
    16'b00110011_01011101 : OUT <= 0;  //51 / 93 = 0
    16'b00110011_01011110 : OUT <= 0;  //51 / 94 = 0
    16'b00110011_01011111 : OUT <= 0;  //51 / 95 = 0
    16'b00110011_01100000 : OUT <= 0;  //51 / 96 = 0
    16'b00110011_01100001 : OUT <= 0;  //51 / 97 = 0
    16'b00110011_01100010 : OUT <= 0;  //51 / 98 = 0
    16'b00110011_01100011 : OUT <= 0;  //51 / 99 = 0
    16'b00110011_01100100 : OUT <= 0;  //51 / 100 = 0
    16'b00110011_01100101 : OUT <= 0;  //51 / 101 = 0
    16'b00110011_01100110 : OUT <= 0;  //51 / 102 = 0
    16'b00110011_01100111 : OUT <= 0;  //51 / 103 = 0
    16'b00110011_01101000 : OUT <= 0;  //51 / 104 = 0
    16'b00110011_01101001 : OUT <= 0;  //51 / 105 = 0
    16'b00110011_01101010 : OUT <= 0;  //51 / 106 = 0
    16'b00110011_01101011 : OUT <= 0;  //51 / 107 = 0
    16'b00110011_01101100 : OUT <= 0;  //51 / 108 = 0
    16'b00110011_01101101 : OUT <= 0;  //51 / 109 = 0
    16'b00110011_01101110 : OUT <= 0;  //51 / 110 = 0
    16'b00110011_01101111 : OUT <= 0;  //51 / 111 = 0
    16'b00110011_01110000 : OUT <= 0;  //51 / 112 = 0
    16'b00110011_01110001 : OUT <= 0;  //51 / 113 = 0
    16'b00110011_01110010 : OUT <= 0;  //51 / 114 = 0
    16'b00110011_01110011 : OUT <= 0;  //51 / 115 = 0
    16'b00110011_01110100 : OUT <= 0;  //51 / 116 = 0
    16'b00110011_01110101 : OUT <= 0;  //51 / 117 = 0
    16'b00110011_01110110 : OUT <= 0;  //51 / 118 = 0
    16'b00110011_01110111 : OUT <= 0;  //51 / 119 = 0
    16'b00110011_01111000 : OUT <= 0;  //51 / 120 = 0
    16'b00110011_01111001 : OUT <= 0;  //51 / 121 = 0
    16'b00110011_01111010 : OUT <= 0;  //51 / 122 = 0
    16'b00110011_01111011 : OUT <= 0;  //51 / 123 = 0
    16'b00110011_01111100 : OUT <= 0;  //51 / 124 = 0
    16'b00110011_01111101 : OUT <= 0;  //51 / 125 = 0
    16'b00110011_01111110 : OUT <= 0;  //51 / 126 = 0
    16'b00110011_01111111 : OUT <= 0;  //51 / 127 = 0
    16'b00110011_10000000 : OUT <= 0;  //51 / 128 = 0
    16'b00110011_10000001 : OUT <= 0;  //51 / 129 = 0
    16'b00110011_10000010 : OUT <= 0;  //51 / 130 = 0
    16'b00110011_10000011 : OUT <= 0;  //51 / 131 = 0
    16'b00110011_10000100 : OUT <= 0;  //51 / 132 = 0
    16'b00110011_10000101 : OUT <= 0;  //51 / 133 = 0
    16'b00110011_10000110 : OUT <= 0;  //51 / 134 = 0
    16'b00110011_10000111 : OUT <= 0;  //51 / 135 = 0
    16'b00110011_10001000 : OUT <= 0;  //51 / 136 = 0
    16'b00110011_10001001 : OUT <= 0;  //51 / 137 = 0
    16'b00110011_10001010 : OUT <= 0;  //51 / 138 = 0
    16'b00110011_10001011 : OUT <= 0;  //51 / 139 = 0
    16'b00110011_10001100 : OUT <= 0;  //51 / 140 = 0
    16'b00110011_10001101 : OUT <= 0;  //51 / 141 = 0
    16'b00110011_10001110 : OUT <= 0;  //51 / 142 = 0
    16'b00110011_10001111 : OUT <= 0;  //51 / 143 = 0
    16'b00110011_10010000 : OUT <= 0;  //51 / 144 = 0
    16'b00110011_10010001 : OUT <= 0;  //51 / 145 = 0
    16'b00110011_10010010 : OUT <= 0;  //51 / 146 = 0
    16'b00110011_10010011 : OUT <= 0;  //51 / 147 = 0
    16'b00110011_10010100 : OUT <= 0;  //51 / 148 = 0
    16'b00110011_10010101 : OUT <= 0;  //51 / 149 = 0
    16'b00110011_10010110 : OUT <= 0;  //51 / 150 = 0
    16'b00110011_10010111 : OUT <= 0;  //51 / 151 = 0
    16'b00110011_10011000 : OUT <= 0;  //51 / 152 = 0
    16'b00110011_10011001 : OUT <= 0;  //51 / 153 = 0
    16'b00110011_10011010 : OUT <= 0;  //51 / 154 = 0
    16'b00110011_10011011 : OUT <= 0;  //51 / 155 = 0
    16'b00110011_10011100 : OUT <= 0;  //51 / 156 = 0
    16'b00110011_10011101 : OUT <= 0;  //51 / 157 = 0
    16'b00110011_10011110 : OUT <= 0;  //51 / 158 = 0
    16'b00110011_10011111 : OUT <= 0;  //51 / 159 = 0
    16'b00110011_10100000 : OUT <= 0;  //51 / 160 = 0
    16'b00110011_10100001 : OUT <= 0;  //51 / 161 = 0
    16'b00110011_10100010 : OUT <= 0;  //51 / 162 = 0
    16'b00110011_10100011 : OUT <= 0;  //51 / 163 = 0
    16'b00110011_10100100 : OUT <= 0;  //51 / 164 = 0
    16'b00110011_10100101 : OUT <= 0;  //51 / 165 = 0
    16'b00110011_10100110 : OUT <= 0;  //51 / 166 = 0
    16'b00110011_10100111 : OUT <= 0;  //51 / 167 = 0
    16'b00110011_10101000 : OUT <= 0;  //51 / 168 = 0
    16'b00110011_10101001 : OUT <= 0;  //51 / 169 = 0
    16'b00110011_10101010 : OUT <= 0;  //51 / 170 = 0
    16'b00110011_10101011 : OUT <= 0;  //51 / 171 = 0
    16'b00110011_10101100 : OUT <= 0;  //51 / 172 = 0
    16'b00110011_10101101 : OUT <= 0;  //51 / 173 = 0
    16'b00110011_10101110 : OUT <= 0;  //51 / 174 = 0
    16'b00110011_10101111 : OUT <= 0;  //51 / 175 = 0
    16'b00110011_10110000 : OUT <= 0;  //51 / 176 = 0
    16'b00110011_10110001 : OUT <= 0;  //51 / 177 = 0
    16'b00110011_10110010 : OUT <= 0;  //51 / 178 = 0
    16'b00110011_10110011 : OUT <= 0;  //51 / 179 = 0
    16'b00110011_10110100 : OUT <= 0;  //51 / 180 = 0
    16'b00110011_10110101 : OUT <= 0;  //51 / 181 = 0
    16'b00110011_10110110 : OUT <= 0;  //51 / 182 = 0
    16'b00110011_10110111 : OUT <= 0;  //51 / 183 = 0
    16'b00110011_10111000 : OUT <= 0;  //51 / 184 = 0
    16'b00110011_10111001 : OUT <= 0;  //51 / 185 = 0
    16'b00110011_10111010 : OUT <= 0;  //51 / 186 = 0
    16'b00110011_10111011 : OUT <= 0;  //51 / 187 = 0
    16'b00110011_10111100 : OUT <= 0;  //51 / 188 = 0
    16'b00110011_10111101 : OUT <= 0;  //51 / 189 = 0
    16'b00110011_10111110 : OUT <= 0;  //51 / 190 = 0
    16'b00110011_10111111 : OUT <= 0;  //51 / 191 = 0
    16'b00110011_11000000 : OUT <= 0;  //51 / 192 = 0
    16'b00110011_11000001 : OUT <= 0;  //51 / 193 = 0
    16'b00110011_11000010 : OUT <= 0;  //51 / 194 = 0
    16'b00110011_11000011 : OUT <= 0;  //51 / 195 = 0
    16'b00110011_11000100 : OUT <= 0;  //51 / 196 = 0
    16'b00110011_11000101 : OUT <= 0;  //51 / 197 = 0
    16'b00110011_11000110 : OUT <= 0;  //51 / 198 = 0
    16'b00110011_11000111 : OUT <= 0;  //51 / 199 = 0
    16'b00110011_11001000 : OUT <= 0;  //51 / 200 = 0
    16'b00110011_11001001 : OUT <= 0;  //51 / 201 = 0
    16'b00110011_11001010 : OUT <= 0;  //51 / 202 = 0
    16'b00110011_11001011 : OUT <= 0;  //51 / 203 = 0
    16'b00110011_11001100 : OUT <= 0;  //51 / 204 = 0
    16'b00110011_11001101 : OUT <= 0;  //51 / 205 = 0
    16'b00110011_11001110 : OUT <= 0;  //51 / 206 = 0
    16'b00110011_11001111 : OUT <= 0;  //51 / 207 = 0
    16'b00110011_11010000 : OUT <= 0;  //51 / 208 = 0
    16'b00110011_11010001 : OUT <= 0;  //51 / 209 = 0
    16'b00110011_11010010 : OUT <= 0;  //51 / 210 = 0
    16'b00110011_11010011 : OUT <= 0;  //51 / 211 = 0
    16'b00110011_11010100 : OUT <= 0;  //51 / 212 = 0
    16'b00110011_11010101 : OUT <= 0;  //51 / 213 = 0
    16'b00110011_11010110 : OUT <= 0;  //51 / 214 = 0
    16'b00110011_11010111 : OUT <= 0;  //51 / 215 = 0
    16'b00110011_11011000 : OUT <= 0;  //51 / 216 = 0
    16'b00110011_11011001 : OUT <= 0;  //51 / 217 = 0
    16'b00110011_11011010 : OUT <= 0;  //51 / 218 = 0
    16'b00110011_11011011 : OUT <= 0;  //51 / 219 = 0
    16'b00110011_11011100 : OUT <= 0;  //51 / 220 = 0
    16'b00110011_11011101 : OUT <= 0;  //51 / 221 = 0
    16'b00110011_11011110 : OUT <= 0;  //51 / 222 = 0
    16'b00110011_11011111 : OUT <= 0;  //51 / 223 = 0
    16'b00110011_11100000 : OUT <= 0;  //51 / 224 = 0
    16'b00110011_11100001 : OUT <= 0;  //51 / 225 = 0
    16'b00110011_11100010 : OUT <= 0;  //51 / 226 = 0
    16'b00110011_11100011 : OUT <= 0;  //51 / 227 = 0
    16'b00110011_11100100 : OUT <= 0;  //51 / 228 = 0
    16'b00110011_11100101 : OUT <= 0;  //51 / 229 = 0
    16'b00110011_11100110 : OUT <= 0;  //51 / 230 = 0
    16'b00110011_11100111 : OUT <= 0;  //51 / 231 = 0
    16'b00110011_11101000 : OUT <= 0;  //51 / 232 = 0
    16'b00110011_11101001 : OUT <= 0;  //51 / 233 = 0
    16'b00110011_11101010 : OUT <= 0;  //51 / 234 = 0
    16'b00110011_11101011 : OUT <= 0;  //51 / 235 = 0
    16'b00110011_11101100 : OUT <= 0;  //51 / 236 = 0
    16'b00110011_11101101 : OUT <= 0;  //51 / 237 = 0
    16'b00110011_11101110 : OUT <= 0;  //51 / 238 = 0
    16'b00110011_11101111 : OUT <= 0;  //51 / 239 = 0
    16'b00110011_11110000 : OUT <= 0;  //51 / 240 = 0
    16'b00110011_11110001 : OUT <= 0;  //51 / 241 = 0
    16'b00110011_11110010 : OUT <= 0;  //51 / 242 = 0
    16'b00110011_11110011 : OUT <= 0;  //51 / 243 = 0
    16'b00110011_11110100 : OUT <= 0;  //51 / 244 = 0
    16'b00110011_11110101 : OUT <= 0;  //51 / 245 = 0
    16'b00110011_11110110 : OUT <= 0;  //51 / 246 = 0
    16'b00110011_11110111 : OUT <= 0;  //51 / 247 = 0
    16'b00110011_11111000 : OUT <= 0;  //51 / 248 = 0
    16'b00110011_11111001 : OUT <= 0;  //51 / 249 = 0
    16'b00110011_11111010 : OUT <= 0;  //51 / 250 = 0
    16'b00110011_11111011 : OUT <= 0;  //51 / 251 = 0
    16'b00110011_11111100 : OUT <= 0;  //51 / 252 = 0
    16'b00110011_11111101 : OUT <= 0;  //51 / 253 = 0
    16'b00110011_11111110 : OUT <= 0;  //51 / 254 = 0
    16'b00110011_11111111 : OUT <= 0;  //51 / 255 = 0
    16'b00110100_00000000 : OUT <= 0;  //52 / 0 = 0
    16'b00110100_00000001 : OUT <= 52;  //52 / 1 = 52
    16'b00110100_00000010 : OUT <= 26;  //52 / 2 = 26
    16'b00110100_00000011 : OUT <= 17;  //52 / 3 = 17
    16'b00110100_00000100 : OUT <= 13;  //52 / 4 = 13
    16'b00110100_00000101 : OUT <= 10;  //52 / 5 = 10
    16'b00110100_00000110 : OUT <= 8;  //52 / 6 = 8
    16'b00110100_00000111 : OUT <= 7;  //52 / 7 = 7
    16'b00110100_00001000 : OUT <= 6;  //52 / 8 = 6
    16'b00110100_00001001 : OUT <= 5;  //52 / 9 = 5
    16'b00110100_00001010 : OUT <= 5;  //52 / 10 = 5
    16'b00110100_00001011 : OUT <= 4;  //52 / 11 = 4
    16'b00110100_00001100 : OUT <= 4;  //52 / 12 = 4
    16'b00110100_00001101 : OUT <= 4;  //52 / 13 = 4
    16'b00110100_00001110 : OUT <= 3;  //52 / 14 = 3
    16'b00110100_00001111 : OUT <= 3;  //52 / 15 = 3
    16'b00110100_00010000 : OUT <= 3;  //52 / 16 = 3
    16'b00110100_00010001 : OUT <= 3;  //52 / 17 = 3
    16'b00110100_00010010 : OUT <= 2;  //52 / 18 = 2
    16'b00110100_00010011 : OUT <= 2;  //52 / 19 = 2
    16'b00110100_00010100 : OUT <= 2;  //52 / 20 = 2
    16'b00110100_00010101 : OUT <= 2;  //52 / 21 = 2
    16'b00110100_00010110 : OUT <= 2;  //52 / 22 = 2
    16'b00110100_00010111 : OUT <= 2;  //52 / 23 = 2
    16'b00110100_00011000 : OUT <= 2;  //52 / 24 = 2
    16'b00110100_00011001 : OUT <= 2;  //52 / 25 = 2
    16'b00110100_00011010 : OUT <= 2;  //52 / 26 = 2
    16'b00110100_00011011 : OUT <= 1;  //52 / 27 = 1
    16'b00110100_00011100 : OUT <= 1;  //52 / 28 = 1
    16'b00110100_00011101 : OUT <= 1;  //52 / 29 = 1
    16'b00110100_00011110 : OUT <= 1;  //52 / 30 = 1
    16'b00110100_00011111 : OUT <= 1;  //52 / 31 = 1
    16'b00110100_00100000 : OUT <= 1;  //52 / 32 = 1
    16'b00110100_00100001 : OUT <= 1;  //52 / 33 = 1
    16'b00110100_00100010 : OUT <= 1;  //52 / 34 = 1
    16'b00110100_00100011 : OUT <= 1;  //52 / 35 = 1
    16'b00110100_00100100 : OUT <= 1;  //52 / 36 = 1
    16'b00110100_00100101 : OUT <= 1;  //52 / 37 = 1
    16'b00110100_00100110 : OUT <= 1;  //52 / 38 = 1
    16'b00110100_00100111 : OUT <= 1;  //52 / 39 = 1
    16'b00110100_00101000 : OUT <= 1;  //52 / 40 = 1
    16'b00110100_00101001 : OUT <= 1;  //52 / 41 = 1
    16'b00110100_00101010 : OUT <= 1;  //52 / 42 = 1
    16'b00110100_00101011 : OUT <= 1;  //52 / 43 = 1
    16'b00110100_00101100 : OUT <= 1;  //52 / 44 = 1
    16'b00110100_00101101 : OUT <= 1;  //52 / 45 = 1
    16'b00110100_00101110 : OUT <= 1;  //52 / 46 = 1
    16'b00110100_00101111 : OUT <= 1;  //52 / 47 = 1
    16'b00110100_00110000 : OUT <= 1;  //52 / 48 = 1
    16'b00110100_00110001 : OUT <= 1;  //52 / 49 = 1
    16'b00110100_00110010 : OUT <= 1;  //52 / 50 = 1
    16'b00110100_00110011 : OUT <= 1;  //52 / 51 = 1
    16'b00110100_00110100 : OUT <= 1;  //52 / 52 = 1
    16'b00110100_00110101 : OUT <= 0;  //52 / 53 = 0
    16'b00110100_00110110 : OUT <= 0;  //52 / 54 = 0
    16'b00110100_00110111 : OUT <= 0;  //52 / 55 = 0
    16'b00110100_00111000 : OUT <= 0;  //52 / 56 = 0
    16'b00110100_00111001 : OUT <= 0;  //52 / 57 = 0
    16'b00110100_00111010 : OUT <= 0;  //52 / 58 = 0
    16'b00110100_00111011 : OUT <= 0;  //52 / 59 = 0
    16'b00110100_00111100 : OUT <= 0;  //52 / 60 = 0
    16'b00110100_00111101 : OUT <= 0;  //52 / 61 = 0
    16'b00110100_00111110 : OUT <= 0;  //52 / 62 = 0
    16'b00110100_00111111 : OUT <= 0;  //52 / 63 = 0
    16'b00110100_01000000 : OUT <= 0;  //52 / 64 = 0
    16'b00110100_01000001 : OUT <= 0;  //52 / 65 = 0
    16'b00110100_01000010 : OUT <= 0;  //52 / 66 = 0
    16'b00110100_01000011 : OUT <= 0;  //52 / 67 = 0
    16'b00110100_01000100 : OUT <= 0;  //52 / 68 = 0
    16'b00110100_01000101 : OUT <= 0;  //52 / 69 = 0
    16'b00110100_01000110 : OUT <= 0;  //52 / 70 = 0
    16'b00110100_01000111 : OUT <= 0;  //52 / 71 = 0
    16'b00110100_01001000 : OUT <= 0;  //52 / 72 = 0
    16'b00110100_01001001 : OUT <= 0;  //52 / 73 = 0
    16'b00110100_01001010 : OUT <= 0;  //52 / 74 = 0
    16'b00110100_01001011 : OUT <= 0;  //52 / 75 = 0
    16'b00110100_01001100 : OUT <= 0;  //52 / 76 = 0
    16'b00110100_01001101 : OUT <= 0;  //52 / 77 = 0
    16'b00110100_01001110 : OUT <= 0;  //52 / 78 = 0
    16'b00110100_01001111 : OUT <= 0;  //52 / 79 = 0
    16'b00110100_01010000 : OUT <= 0;  //52 / 80 = 0
    16'b00110100_01010001 : OUT <= 0;  //52 / 81 = 0
    16'b00110100_01010010 : OUT <= 0;  //52 / 82 = 0
    16'b00110100_01010011 : OUT <= 0;  //52 / 83 = 0
    16'b00110100_01010100 : OUT <= 0;  //52 / 84 = 0
    16'b00110100_01010101 : OUT <= 0;  //52 / 85 = 0
    16'b00110100_01010110 : OUT <= 0;  //52 / 86 = 0
    16'b00110100_01010111 : OUT <= 0;  //52 / 87 = 0
    16'b00110100_01011000 : OUT <= 0;  //52 / 88 = 0
    16'b00110100_01011001 : OUT <= 0;  //52 / 89 = 0
    16'b00110100_01011010 : OUT <= 0;  //52 / 90 = 0
    16'b00110100_01011011 : OUT <= 0;  //52 / 91 = 0
    16'b00110100_01011100 : OUT <= 0;  //52 / 92 = 0
    16'b00110100_01011101 : OUT <= 0;  //52 / 93 = 0
    16'b00110100_01011110 : OUT <= 0;  //52 / 94 = 0
    16'b00110100_01011111 : OUT <= 0;  //52 / 95 = 0
    16'b00110100_01100000 : OUT <= 0;  //52 / 96 = 0
    16'b00110100_01100001 : OUT <= 0;  //52 / 97 = 0
    16'b00110100_01100010 : OUT <= 0;  //52 / 98 = 0
    16'b00110100_01100011 : OUT <= 0;  //52 / 99 = 0
    16'b00110100_01100100 : OUT <= 0;  //52 / 100 = 0
    16'b00110100_01100101 : OUT <= 0;  //52 / 101 = 0
    16'b00110100_01100110 : OUT <= 0;  //52 / 102 = 0
    16'b00110100_01100111 : OUT <= 0;  //52 / 103 = 0
    16'b00110100_01101000 : OUT <= 0;  //52 / 104 = 0
    16'b00110100_01101001 : OUT <= 0;  //52 / 105 = 0
    16'b00110100_01101010 : OUT <= 0;  //52 / 106 = 0
    16'b00110100_01101011 : OUT <= 0;  //52 / 107 = 0
    16'b00110100_01101100 : OUT <= 0;  //52 / 108 = 0
    16'b00110100_01101101 : OUT <= 0;  //52 / 109 = 0
    16'b00110100_01101110 : OUT <= 0;  //52 / 110 = 0
    16'b00110100_01101111 : OUT <= 0;  //52 / 111 = 0
    16'b00110100_01110000 : OUT <= 0;  //52 / 112 = 0
    16'b00110100_01110001 : OUT <= 0;  //52 / 113 = 0
    16'b00110100_01110010 : OUT <= 0;  //52 / 114 = 0
    16'b00110100_01110011 : OUT <= 0;  //52 / 115 = 0
    16'b00110100_01110100 : OUT <= 0;  //52 / 116 = 0
    16'b00110100_01110101 : OUT <= 0;  //52 / 117 = 0
    16'b00110100_01110110 : OUT <= 0;  //52 / 118 = 0
    16'b00110100_01110111 : OUT <= 0;  //52 / 119 = 0
    16'b00110100_01111000 : OUT <= 0;  //52 / 120 = 0
    16'b00110100_01111001 : OUT <= 0;  //52 / 121 = 0
    16'b00110100_01111010 : OUT <= 0;  //52 / 122 = 0
    16'b00110100_01111011 : OUT <= 0;  //52 / 123 = 0
    16'b00110100_01111100 : OUT <= 0;  //52 / 124 = 0
    16'b00110100_01111101 : OUT <= 0;  //52 / 125 = 0
    16'b00110100_01111110 : OUT <= 0;  //52 / 126 = 0
    16'b00110100_01111111 : OUT <= 0;  //52 / 127 = 0
    16'b00110100_10000000 : OUT <= 0;  //52 / 128 = 0
    16'b00110100_10000001 : OUT <= 0;  //52 / 129 = 0
    16'b00110100_10000010 : OUT <= 0;  //52 / 130 = 0
    16'b00110100_10000011 : OUT <= 0;  //52 / 131 = 0
    16'b00110100_10000100 : OUT <= 0;  //52 / 132 = 0
    16'b00110100_10000101 : OUT <= 0;  //52 / 133 = 0
    16'b00110100_10000110 : OUT <= 0;  //52 / 134 = 0
    16'b00110100_10000111 : OUT <= 0;  //52 / 135 = 0
    16'b00110100_10001000 : OUT <= 0;  //52 / 136 = 0
    16'b00110100_10001001 : OUT <= 0;  //52 / 137 = 0
    16'b00110100_10001010 : OUT <= 0;  //52 / 138 = 0
    16'b00110100_10001011 : OUT <= 0;  //52 / 139 = 0
    16'b00110100_10001100 : OUT <= 0;  //52 / 140 = 0
    16'b00110100_10001101 : OUT <= 0;  //52 / 141 = 0
    16'b00110100_10001110 : OUT <= 0;  //52 / 142 = 0
    16'b00110100_10001111 : OUT <= 0;  //52 / 143 = 0
    16'b00110100_10010000 : OUT <= 0;  //52 / 144 = 0
    16'b00110100_10010001 : OUT <= 0;  //52 / 145 = 0
    16'b00110100_10010010 : OUT <= 0;  //52 / 146 = 0
    16'b00110100_10010011 : OUT <= 0;  //52 / 147 = 0
    16'b00110100_10010100 : OUT <= 0;  //52 / 148 = 0
    16'b00110100_10010101 : OUT <= 0;  //52 / 149 = 0
    16'b00110100_10010110 : OUT <= 0;  //52 / 150 = 0
    16'b00110100_10010111 : OUT <= 0;  //52 / 151 = 0
    16'b00110100_10011000 : OUT <= 0;  //52 / 152 = 0
    16'b00110100_10011001 : OUT <= 0;  //52 / 153 = 0
    16'b00110100_10011010 : OUT <= 0;  //52 / 154 = 0
    16'b00110100_10011011 : OUT <= 0;  //52 / 155 = 0
    16'b00110100_10011100 : OUT <= 0;  //52 / 156 = 0
    16'b00110100_10011101 : OUT <= 0;  //52 / 157 = 0
    16'b00110100_10011110 : OUT <= 0;  //52 / 158 = 0
    16'b00110100_10011111 : OUT <= 0;  //52 / 159 = 0
    16'b00110100_10100000 : OUT <= 0;  //52 / 160 = 0
    16'b00110100_10100001 : OUT <= 0;  //52 / 161 = 0
    16'b00110100_10100010 : OUT <= 0;  //52 / 162 = 0
    16'b00110100_10100011 : OUT <= 0;  //52 / 163 = 0
    16'b00110100_10100100 : OUT <= 0;  //52 / 164 = 0
    16'b00110100_10100101 : OUT <= 0;  //52 / 165 = 0
    16'b00110100_10100110 : OUT <= 0;  //52 / 166 = 0
    16'b00110100_10100111 : OUT <= 0;  //52 / 167 = 0
    16'b00110100_10101000 : OUT <= 0;  //52 / 168 = 0
    16'b00110100_10101001 : OUT <= 0;  //52 / 169 = 0
    16'b00110100_10101010 : OUT <= 0;  //52 / 170 = 0
    16'b00110100_10101011 : OUT <= 0;  //52 / 171 = 0
    16'b00110100_10101100 : OUT <= 0;  //52 / 172 = 0
    16'b00110100_10101101 : OUT <= 0;  //52 / 173 = 0
    16'b00110100_10101110 : OUT <= 0;  //52 / 174 = 0
    16'b00110100_10101111 : OUT <= 0;  //52 / 175 = 0
    16'b00110100_10110000 : OUT <= 0;  //52 / 176 = 0
    16'b00110100_10110001 : OUT <= 0;  //52 / 177 = 0
    16'b00110100_10110010 : OUT <= 0;  //52 / 178 = 0
    16'b00110100_10110011 : OUT <= 0;  //52 / 179 = 0
    16'b00110100_10110100 : OUT <= 0;  //52 / 180 = 0
    16'b00110100_10110101 : OUT <= 0;  //52 / 181 = 0
    16'b00110100_10110110 : OUT <= 0;  //52 / 182 = 0
    16'b00110100_10110111 : OUT <= 0;  //52 / 183 = 0
    16'b00110100_10111000 : OUT <= 0;  //52 / 184 = 0
    16'b00110100_10111001 : OUT <= 0;  //52 / 185 = 0
    16'b00110100_10111010 : OUT <= 0;  //52 / 186 = 0
    16'b00110100_10111011 : OUT <= 0;  //52 / 187 = 0
    16'b00110100_10111100 : OUT <= 0;  //52 / 188 = 0
    16'b00110100_10111101 : OUT <= 0;  //52 / 189 = 0
    16'b00110100_10111110 : OUT <= 0;  //52 / 190 = 0
    16'b00110100_10111111 : OUT <= 0;  //52 / 191 = 0
    16'b00110100_11000000 : OUT <= 0;  //52 / 192 = 0
    16'b00110100_11000001 : OUT <= 0;  //52 / 193 = 0
    16'b00110100_11000010 : OUT <= 0;  //52 / 194 = 0
    16'b00110100_11000011 : OUT <= 0;  //52 / 195 = 0
    16'b00110100_11000100 : OUT <= 0;  //52 / 196 = 0
    16'b00110100_11000101 : OUT <= 0;  //52 / 197 = 0
    16'b00110100_11000110 : OUT <= 0;  //52 / 198 = 0
    16'b00110100_11000111 : OUT <= 0;  //52 / 199 = 0
    16'b00110100_11001000 : OUT <= 0;  //52 / 200 = 0
    16'b00110100_11001001 : OUT <= 0;  //52 / 201 = 0
    16'b00110100_11001010 : OUT <= 0;  //52 / 202 = 0
    16'b00110100_11001011 : OUT <= 0;  //52 / 203 = 0
    16'b00110100_11001100 : OUT <= 0;  //52 / 204 = 0
    16'b00110100_11001101 : OUT <= 0;  //52 / 205 = 0
    16'b00110100_11001110 : OUT <= 0;  //52 / 206 = 0
    16'b00110100_11001111 : OUT <= 0;  //52 / 207 = 0
    16'b00110100_11010000 : OUT <= 0;  //52 / 208 = 0
    16'b00110100_11010001 : OUT <= 0;  //52 / 209 = 0
    16'b00110100_11010010 : OUT <= 0;  //52 / 210 = 0
    16'b00110100_11010011 : OUT <= 0;  //52 / 211 = 0
    16'b00110100_11010100 : OUT <= 0;  //52 / 212 = 0
    16'b00110100_11010101 : OUT <= 0;  //52 / 213 = 0
    16'b00110100_11010110 : OUT <= 0;  //52 / 214 = 0
    16'b00110100_11010111 : OUT <= 0;  //52 / 215 = 0
    16'b00110100_11011000 : OUT <= 0;  //52 / 216 = 0
    16'b00110100_11011001 : OUT <= 0;  //52 / 217 = 0
    16'b00110100_11011010 : OUT <= 0;  //52 / 218 = 0
    16'b00110100_11011011 : OUT <= 0;  //52 / 219 = 0
    16'b00110100_11011100 : OUT <= 0;  //52 / 220 = 0
    16'b00110100_11011101 : OUT <= 0;  //52 / 221 = 0
    16'b00110100_11011110 : OUT <= 0;  //52 / 222 = 0
    16'b00110100_11011111 : OUT <= 0;  //52 / 223 = 0
    16'b00110100_11100000 : OUT <= 0;  //52 / 224 = 0
    16'b00110100_11100001 : OUT <= 0;  //52 / 225 = 0
    16'b00110100_11100010 : OUT <= 0;  //52 / 226 = 0
    16'b00110100_11100011 : OUT <= 0;  //52 / 227 = 0
    16'b00110100_11100100 : OUT <= 0;  //52 / 228 = 0
    16'b00110100_11100101 : OUT <= 0;  //52 / 229 = 0
    16'b00110100_11100110 : OUT <= 0;  //52 / 230 = 0
    16'b00110100_11100111 : OUT <= 0;  //52 / 231 = 0
    16'b00110100_11101000 : OUT <= 0;  //52 / 232 = 0
    16'b00110100_11101001 : OUT <= 0;  //52 / 233 = 0
    16'b00110100_11101010 : OUT <= 0;  //52 / 234 = 0
    16'b00110100_11101011 : OUT <= 0;  //52 / 235 = 0
    16'b00110100_11101100 : OUT <= 0;  //52 / 236 = 0
    16'b00110100_11101101 : OUT <= 0;  //52 / 237 = 0
    16'b00110100_11101110 : OUT <= 0;  //52 / 238 = 0
    16'b00110100_11101111 : OUT <= 0;  //52 / 239 = 0
    16'b00110100_11110000 : OUT <= 0;  //52 / 240 = 0
    16'b00110100_11110001 : OUT <= 0;  //52 / 241 = 0
    16'b00110100_11110010 : OUT <= 0;  //52 / 242 = 0
    16'b00110100_11110011 : OUT <= 0;  //52 / 243 = 0
    16'b00110100_11110100 : OUT <= 0;  //52 / 244 = 0
    16'b00110100_11110101 : OUT <= 0;  //52 / 245 = 0
    16'b00110100_11110110 : OUT <= 0;  //52 / 246 = 0
    16'b00110100_11110111 : OUT <= 0;  //52 / 247 = 0
    16'b00110100_11111000 : OUT <= 0;  //52 / 248 = 0
    16'b00110100_11111001 : OUT <= 0;  //52 / 249 = 0
    16'b00110100_11111010 : OUT <= 0;  //52 / 250 = 0
    16'b00110100_11111011 : OUT <= 0;  //52 / 251 = 0
    16'b00110100_11111100 : OUT <= 0;  //52 / 252 = 0
    16'b00110100_11111101 : OUT <= 0;  //52 / 253 = 0
    16'b00110100_11111110 : OUT <= 0;  //52 / 254 = 0
    16'b00110100_11111111 : OUT <= 0;  //52 / 255 = 0
    16'b00110101_00000000 : OUT <= 0;  //53 / 0 = 0
    16'b00110101_00000001 : OUT <= 53;  //53 / 1 = 53
    16'b00110101_00000010 : OUT <= 26;  //53 / 2 = 26
    16'b00110101_00000011 : OUT <= 17;  //53 / 3 = 17
    16'b00110101_00000100 : OUT <= 13;  //53 / 4 = 13
    16'b00110101_00000101 : OUT <= 10;  //53 / 5 = 10
    16'b00110101_00000110 : OUT <= 8;  //53 / 6 = 8
    16'b00110101_00000111 : OUT <= 7;  //53 / 7 = 7
    16'b00110101_00001000 : OUT <= 6;  //53 / 8 = 6
    16'b00110101_00001001 : OUT <= 5;  //53 / 9 = 5
    16'b00110101_00001010 : OUT <= 5;  //53 / 10 = 5
    16'b00110101_00001011 : OUT <= 4;  //53 / 11 = 4
    16'b00110101_00001100 : OUT <= 4;  //53 / 12 = 4
    16'b00110101_00001101 : OUT <= 4;  //53 / 13 = 4
    16'b00110101_00001110 : OUT <= 3;  //53 / 14 = 3
    16'b00110101_00001111 : OUT <= 3;  //53 / 15 = 3
    16'b00110101_00010000 : OUT <= 3;  //53 / 16 = 3
    16'b00110101_00010001 : OUT <= 3;  //53 / 17 = 3
    16'b00110101_00010010 : OUT <= 2;  //53 / 18 = 2
    16'b00110101_00010011 : OUT <= 2;  //53 / 19 = 2
    16'b00110101_00010100 : OUT <= 2;  //53 / 20 = 2
    16'b00110101_00010101 : OUT <= 2;  //53 / 21 = 2
    16'b00110101_00010110 : OUT <= 2;  //53 / 22 = 2
    16'b00110101_00010111 : OUT <= 2;  //53 / 23 = 2
    16'b00110101_00011000 : OUT <= 2;  //53 / 24 = 2
    16'b00110101_00011001 : OUT <= 2;  //53 / 25 = 2
    16'b00110101_00011010 : OUT <= 2;  //53 / 26 = 2
    16'b00110101_00011011 : OUT <= 1;  //53 / 27 = 1
    16'b00110101_00011100 : OUT <= 1;  //53 / 28 = 1
    16'b00110101_00011101 : OUT <= 1;  //53 / 29 = 1
    16'b00110101_00011110 : OUT <= 1;  //53 / 30 = 1
    16'b00110101_00011111 : OUT <= 1;  //53 / 31 = 1
    16'b00110101_00100000 : OUT <= 1;  //53 / 32 = 1
    16'b00110101_00100001 : OUT <= 1;  //53 / 33 = 1
    16'b00110101_00100010 : OUT <= 1;  //53 / 34 = 1
    16'b00110101_00100011 : OUT <= 1;  //53 / 35 = 1
    16'b00110101_00100100 : OUT <= 1;  //53 / 36 = 1
    16'b00110101_00100101 : OUT <= 1;  //53 / 37 = 1
    16'b00110101_00100110 : OUT <= 1;  //53 / 38 = 1
    16'b00110101_00100111 : OUT <= 1;  //53 / 39 = 1
    16'b00110101_00101000 : OUT <= 1;  //53 / 40 = 1
    16'b00110101_00101001 : OUT <= 1;  //53 / 41 = 1
    16'b00110101_00101010 : OUT <= 1;  //53 / 42 = 1
    16'b00110101_00101011 : OUT <= 1;  //53 / 43 = 1
    16'b00110101_00101100 : OUT <= 1;  //53 / 44 = 1
    16'b00110101_00101101 : OUT <= 1;  //53 / 45 = 1
    16'b00110101_00101110 : OUT <= 1;  //53 / 46 = 1
    16'b00110101_00101111 : OUT <= 1;  //53 / 47 = 1
    16'b00110101_00110000 : OUT <= 1;  //53 / 48 = 1
    16'b00110101_00110001 : OUT <= 1;  //53 / 49 = 1
    16'b00110101_00110010 : OUT <= 1;  //53 / 50 = 1
    16'b00110101_00110011 : OUT <= 1;  //53 / 51 = 1
    16'b00110101_00110100 : OUT <= 1;  //53 / 52 = 1
    16'b00110101_00110101 : OUT <= 1;  //53 / 53 = 1
    16'b00110101_00110110 : OUT <= 0;  //53 / 54 = 0
    16'b00110101_00110111 : OUT <= 0;  //53 / 55 = 0
    16'b00110101_00111000 : OUT <= 0;  //53 / 56 = 0
    16'b00110101_00111001 : OUT <= 0;  //53 / 57 = 0
    16'b00110101_00111010 : OUT <= 0;  //53 / 58 = 0
    16'b00110101_00111011 : OUT <= 0;  //53 / 59 = 0
    16'b00110101_00111100 : OUT <= 0;  //53 / 60 = 0
    16'b00110101_00111101 : OUT <= 0;  //53 / 61 = 0
    16'b00110101_00111110 : OUT <= 0;  //53 / 62 = 0
    16'b00110101_00111111 : OUT <= 0;  //53 / 63 = 0
    16'b00110101_01000000 : OUT <= 0;  //53 / 64 = 0
    16'b00110101_01000001 : OUT <= 0;  //53 / 65 = 0
    16'b00110101_01000010 : OUT <= 0;  //53 / 66 = 0
    16'b00110101_01000011 : OUT <= 0;  //53 / 67 = 0
    16'b00110101_01000100 : OUT <= 0;  //53 / 68 = 0
    16'b00110101_01000101 : OUT <= 0;  //53 / 69 = 0
    16'b00110101_01000110 : OUT <= 0;  //53 / 70 = 0
    16'b00110101_01000111 : OUT <= 0;  //53 / 71 = 0
    16'b00110101_01001000 : OUT <= 0;  //53 / 72 = 0
    16'b00110101_01001001 : OUT <= 0;  //53 / 73 = 0
    16'b00110101_01001010 : OUT <= 0;  //53 / 74 = 0
    16'b00110101_01001011 : OUT <= 0;  //53 / 75 = 0
    16'b00110101_01001100 : OUT <= 0;  //53 / 76 = 0
    16'b00110101_01001101 : OUT <= 0;  //53 / 77 = 0
    16'b00110101_01001110 : OUT <= 0;  //53 / 78 = 0
    16'b00110101_01001111 : OUT <= 0;  //53 / 79 = 0
    16'b00110101_01010000 : OUT <= 0;  //53 / 80 = 0
    16'b00110101_01010001 : OUT <= 0;  //53 / 81 = 0
    16'b00110101_01010010 : OUT <= 0;  //53 / 82 = 0
    16'b00110101_01010011 : OUT <= 0;  //53 / 83 = 0
    16'b00110101_01010100 : OUT <= 0;  //53 / 84 = 0
    16'b00110101_01010101 : OUT <= 0;  //53 / 85 = 0
    16'b00110101_01010110 : OUT <= 0;  //53 / 86 = 0
    16'b00110101_01010111 : OUT <= 0;  //53 / 87 = 0
    16'b00110101_01011000 : OUT <= 0;  //53 / 88 = 0
    16'b00110101_01011001 : OUT <= 0;  //53 / 89 = 0
    16'b00110101_01011010 : OUT <= 0;  //53 / 90 = 0
    16'b00110101_01011011 : OUT <= 0;  //53 / 91 = 0
    16'b00110101_01011100 : OUT <= 0;  //53 / 92 = 0
    16'b00110101_01011101 : OUT <= 0;  //53 / 93 = 0
    16'b00110101_01011110 : OUT <= 0;  //53 / 94 = 0
    16'b00110101_01011111 : OUT <= 0;  //53 / 95 = 0
    16'b00110101_01100000 : OUT <= 0;  //53 / 96 = 0
    16'b00110101_01100001 : OUT <= 0;  //53 / 97 = 0
    16'b00110101_01100010 : OUT <= 0;  //53 / 98 = 0
    16'b00110101_01100011 : OUT <= 0;  //53 / 99 = 0
    16'b00110101_01100100 : OUT <= 0;  //53 / 100 = 0
    16'b00110101_01100101 : OUT <= 0;  //53 / 101 = 0
    16'b00110101_01100110 : OUT <= 0;  //53 / 102 = 0
    16'b00110101_01100111 : OUT <= 0;  //53 / 103 = 0
    16'b00110101_01101000 : OUT <= 0;  //53 / 104 = 0
    16'b00110101_01101001 : OUT <= 0;  //53 / 105 = 0
    16'b00110101_01101010 : OUT <= 0;  //53 / 106 = 0
    16'b00110101_01101011 : OUT <= 0;  //53 / 107 = 0
    16'b00110101_01101100 : OUT <= 0;  //53 / 108 = 0
    16'b00110101_01101101 : OUT <= 0;  //53 / 109 = 0
    16'b00110101_01101110 : OUT <= 0;  //53 / 110 = 0
    16'b00110101_01101111 : OUT <= 0;  //53 / 111 = 0
    16'b00110101_01110000 : OUT <= 0;  //53 / 112 = 0
    16'b00110101_01110001 : OUT <= 0;  //53 / 113 = 0
    16'b00110101_01110010 : OUT <= 0;  //53 / 114 = 0
    16'b00110101_01110011 : OUT <= 0;  //53 / 115 = 0
    16'b00110101_01110100 : OUT <= 0;  //53 / 116 = 0
    16'b00110101_01110101 : OUT <= 0;  //53 / 117 = 0
    16'b00110101_01110110 : OUT <= 0;  //53 / 118 = 0
    16'b00110101_01110111 : OUT <= 0;  //53 / 119 = 0
    16'b00110101_01111000 : OUT <= 0;  //53 / 120 = 0
    16'b00110101_01111001 : OUT <= 0;  //53 / 121 = 0
    16'b00110101_01111010 : OUT <= 0;  //53 / 122 = 0
    16'b00110101_01111011 : OUT <= 0;  //53 / 123 = 0
    16'b00110101_01111100 : OUT <= 0;  //53 / 124 = 0
    16'b00110101_01111101 : OUT <= 0;  //53 / 125 = 0
    16'b00110101_01111110 : OUT <= 0;  //53 / 126 = 0
    16'b00110101_01111111 : OUT <= 0;  //53 / 127 = 0
    16'b00110101_10000000 : OUT <= 0;  //53 / 128 = 0
    16'b00110101_10000001 : OUT <= 0;  //53 / 129 = 0
    16'b00110101_10000010 : OUT <= 0;  //53 / 130 = 0
    16'b00110101_10000011 : OUT <= 0;  //53 / 131 = 0
    16'b00110101_10000100 : OUT <= 0;  //53 / 132 = 0
    16'b00110101_10000101 : OUT <= 0;  //53 / 133 = 0
    16'b00110101_10000110 : OUT <= 0;  //53 / 134 = 0
    16'b00110101_10000111 : OUT <= 0;  //53 / 135 = 0
    16'b00110101_10001000 : OUT <= 0;  //53 / 136 = 0
    16'b00110101_10001001 : OUT <= 0;  //53 / 137 = 0
    16'b00110101_10001010 : OUT <= 0;  //53 / 138 = 0
    16'b00110101_10001011 : OUT <= 0;  //53 / 139 = 0
    16'b00110101_10001100 : OUT <= 0;  //53 / 140 = 0
    16'b00110101_10001101 : OUT <= 0;  //53 / 141 = 0
    16'b00110101_10001110 : OUT <= 0;  //53 / 142 = 0
    16'b00110101_10001111 : OUT <= 0;  //53 / 143 = 0
    16'b00110101_10010000 : OUT <= 0;  //53 / 144 = 0
    16'b00110101_10010001 : OUT <= 0;  //53 / 145 = 0
    16'b00110101_10010010 : OUT <= 0;  //53 / 146 = 0
    16'b00110101_10010011 : OUT <= 0;  //53 / 147 = 0
    16'b00110101_10010100 : OUT <= 0;  //53 / 148 = 0
    16'b00110101_10010101 : OUT <= 0;  //53 / 149 = 0
    16'b00110101_10010110 : OUT <= 0;  //53 / 150 = 0
    16'b00110101_10010111 : OUT <= 0;  //53 / 151 = 0
    16'b00110101_10011000 : OUT <= 0;  //53 / 152 = 0
    16'b00110101_10011001 : OUT <= 0;  //53 / 153 = 0
    16'b00110101_10011010 : OUT <= 0;  //53 / 154 = 0
    16'b00110101_10011011 : OUT <= 0;  //53 / 155 = 0
    16'b00110101_10011100 : OUT <= 0;  //53 / 156 = 0
    16'b00110101_10011101 : OUT <= 0;  //53 / 157 = 0
    16'b00110101_10011110 : OUT <= 0;  //53 / 158 = 0
    16'b00110101_10011111 : OUT <= 0;  //53 / 159 = 0
    16'b00110101_10100000 : OUT <= 0;  //53 / 160 = 0
    16'b00110101_10100001 : OUT <= 0;  //53 / 161 = 0
    16'b00110101_10100010 : OUT <= 0;  //53 / 162 = 0
    16'b00110101_10100011 : OUT <= 0;  //53 / 163 = 0
    16'b00110101_10100100 : OUT <= 0;  //53 / 164 = 0
    16'b00110101_10100101 : OUT <= 0;  //53 / 165 = 0
    16'b00110101_10100110 : OUT <= 0;  //53 / 166 = 0
    16'b00110101_10100111 : OUT <= 0;  //53 / 167 = 0
    16'b00110101_10101000 : OUT <= 0;  //53 / 168 = 0
    16'b00110101_10101001 : OUT <= 0;  //53 / 169 = 0
    16'b00110101_10101010 : OUT <= 0;  //53 / 170 = 0
    16'b00110101_10101011 : OUT <= 0;  //53 / 171 = 0
    16'b00110101_10101100 : OUT <= 0;  //53 / 172 = 0
    16'b00110101_10101101 : OUT <= 0;  //53 / 173 = 0
    16'b00110101_10101110 : OUT <= 0;  //53 / 174 = 0
    16'b00110101_10101111 : OUT <= 0;  //53 / 175 = 0
    16'b00110101_10110000 : OUT <= 0;  //53 / 176 = 0
    16'b00110101_10110001 : OUT <= 0;  //53 / 177 = 0
    16'b00110101_10110010 : OUT <= 0;  //53 / 178 = 0
    16'b00110101_10110011 : OUT <= 0;  //53 / 179 = 0
    16'b00110101_10110100 : OUT <= 0;  //53 / 180 = 0
    16'b00110101_10110101 : OUT <= 0;  //53 / 181 = 0
    16'b00110101_10110110 : OUT <= 0;  //53 / 182 = 0
    16'b00110101_10110111 : OUT <= 0;  //53 / 183 = 0
    16'b00110101_10111000 : OUT <= 0;  //53 / 184 = 0
    16'b00110101_10111001 : OUT <= 0;  //53 / 185 = 0
    16'b00110101_10111010 : OUT <= 0;  //53 / 186 = 0
    16'b00110101_10111011 : OUT <= 0;  //53 / 187 = 0
    16'b00110101_10111100 : OUT <= 0;  //53 / 188 = 0
    16'b00110101_10111101 : OUT <= 0;  //53 / 189 = 0
    16'b00110101_10111110 : OUT <= 0;  //53 / 190 = 0
    16'b00110101_10111111 : OUT <= 0;  //53 / 191 = 0
    16'b00110101_11000000 : OUT <= 0;  //53 / 192 = 0
    16'b00110101_11000001 : OUT <= 0;  //53 / 193 = 0
    16'b00110101_11000010 : OUT <= 0;  //53 / 194 = 0
    16'b00110101_11000011 : OUT <= 0;  //53 / 195 = 0
    16'b00110101_11000100 : OUT <= 0;  //53 / 196 = 0
    16'b00110101_11000101 : OUT <= 0;  //53 / 197 = 0
    16'b00110101_11000110 : OUT <= 0;  //53 / 198 = 0
    16'b00110101_11000111 : OUT <= 0;  //53 / 199 = 0
    16'b00110101_11001000 : OUT <= 0;  //53 / 200 = 0
    16'b00110101_11001001 : OUT <= 0;  //53 / 201 = 0
    16'b00110101_11001010 : OUT <= 0;  //53 / 202 = 0
    16'b00110101_11001011 : OUT <= 0;  //53 / 203 = 0
    16'b00110101_11001100 : OUT <= 0;  //53 / 204 = 0
    16'b00110101_11001101 : OUT <= 0;  //53 / 205 = 0
    16'b00110101_11001110 : OUT <= 0;  //53 / 206 = 0
    16'b00110101_11001111 : OUT <= 0;  //53 / 207 = 0
    16'b00110101_11010000 : OUT <= 0;  //53 / 208 = 0
    16'b00110101_11010001 : OUT <= 0;  //53 / 209 = 0
    16'b00110101_11010010 : OUT <= 0;  //53 / 210 = 0
    16'b00110101_11010011 : OUT <= 0;  //53 / 211 = 0
    16'b00110101_11010100 : OUT <= 0;  //53 / 212 = 0
    16'b00110101_11010101 : OUT <= 0;  //53 / 213 = 0
    16'b00110101_11010110 : OUT <= 0;  //53 / 214 = 0
    16'b00110101_11010111 : OUT <= 0;  //53 / 215 = 0
    16'b00110101_11011000 : OUT <= 0;  //53 / 216 = 0
    16'b00110101_11011001 : OUT <= 0;  //53 / 217 = 0
    16'b00110101_11011010 : OUT <= 0;  //53 / 218 = 0
    16'b00110101_11011011 : OUT <= 0;  //53 / 219 = 0
    16'b00110101_11011100 : OUT <= 0;  //53 / 220 = 0
    16'b00110101_11011101 : OUT <= 0;  //53 / 221 = 0
    16'b00110101_11011110 : OUT <= 0;  //53 / 222 = 0
    16'b00110101_11011111 : OUT <= 0;  //53 / 223 = 0
    16'b00110101_11100000 : OUT <= 0;  //53 / 224 = 0
    16'b00110101_11100001 : OUT <= 0;  //53 / 225 = 0
    16'b00110101_11100010 : OUT <= 0;  //53 / 226 = 0
    16'b00110101_11100011 : OUT <= 0;  //53 / 227 = 0
    16'b00110101_11100100 : OUT <= 0;  //53 / 228 = 0
    16'b00110101_11100101 : OUT <= 0;  //53 / 229 = 0
    16'b00110101_11100110 : OUT <= 0;  //53 / 230 = 0
    16'b00110101_11100111 : OUT <= 0;  //53 / 231 = 0
    16'b00110101_11101000 : OUT <= 0;  //53 / 232 = 0
    16'b00110101_11101001 : OUT <= 0;  //53 / 233 = 0
    16'b00110101_11101010 : OUT <= 0;  //53 / 234 = 0
    16'b00110101_11101011 : OUT <= 0;  //53 / 235 = 0
    16'b00110101_11101100 : OUT <= 0;  //53 / 236 = 0
    16'b00110101_11101101 : OUT <= 0;  //53 / 237 = 0
    16'b00110101_11101110 : OUT <= 0;  //53 / 238 = 0
    16'b00110101_11101111 : OUT <= 0;  //53 / 239 = 0
    16'b00110101_11110000 : OUT <= 0;  //53 / 240 = 0
    16'b00110101_11110001 : OUT <= 0;  //53 / 241 = 0
    16'b00110101_11110010 : OUT <= 0;  //53 / 242 = 0
    16'b00110101_11110011 : OUT <= 0;  //53 / 243 = 0
    16'b00110101_11110100 : OUT <= 0;  //53 / 244 = 0
    16'b00110101_11110101 : OUT <= 0;  //53 / 245 = 0
    16'b00110101_11110110 : OUT <= 0;  //53 / 246 = 0
    16'b00110101_11110111 : OUT <= 0;  //53 / 247 = 0
    16'b00110101_11111000 : OUT <= 0;  //53 / 248 = 0
    16'b00110101_11111001 : OUT <= 0;  //53 / 249 = 0
    16'b00110101_11111010 : OUT <= 0;  //53 / 250 = 0
    16'b00110101_11111011 : OUT <= 0;  //53 / 251 = 0
    16'b00110101_11111100 : OUT <= 0;  //53 / 252 = 0
    16'b00110101_11111101 : OUT <= 0;  //53 / 253 = 0
    16'b00110101_11111110 : OUT <= 0;  //53 / 254 = 0
    16'b00110101_11111111 : OUT <= 0;  //53 / 255 = 0
    16'b00110110_00000000 : OUT <= 0;  //54 / 0 = 0
    16'b00110110_00000001 : OUT <= 54;  //54 / 1 = 54
    16'b00110110_00000010 : OUT <= 27;  //54 / 2 = 27
    16'b00110110_00000011 : OUT <= 18;  //54 / 3 = 18
    16'b00110110_00000100 : OUT <= 13;  //54 / 4 = 13
    16'b00110110_00000101 : OUT <= 10;  //54 / 5 = 10
    16'b00110110_00000110 : OUT <= 9;  //54 / 6 = 9
    16'b00110110_00000111 : OUT <= 7;  //54 / 7 = 7
    16'b00110110_00001000 : OUT <= 6;  //54 / 8 = 6
    16'b00110110_00001001 : OUT <= 6;  //54 / 9 = 6
    16'b00110110_00001010 : OUT <= 5;  //54 / 10 = 5
    16'b00110110_00001011 : OUT <= 4;  //54 / 11 = 4
    16'b00110110_00001100 : OUT <= 4;  //54 / 12 = 4
    16'b00110110_00001101 : OUT <= 4;  //54 / 13 = 4
    16'b00110110_00001110 : OUT <= 3;  //54 / 14 = 3
    16'b00110110_00001111 : OUT <= 3;  //54 / 15 = 3
    16'b00110110_00010000 : OUT <= 3;  //54 / 16 = 3
    16'b00110110_00010001 : OUT <= 3;  //54 / 17 = 3
    16'b00110110_00010010 : OUT <= 3;  //54 / 18 = 3
    16'b00110110_00010011 : OUT <= 2;  //54 / 19 = 2
    16'b00110110_00010100 : OUT <= 2;  //54 / 20 = 2
    16'b00110110_00010101 : OUT <= 2;  //54 / 21 = 2
    16'b00110110_00010110 : OUT <= 2;  //54 / 22 = 2
    16'b00110110_00010111 : OUT <= 2;  //54 / 23 = 2
    16'b00110110_00011000 : OUT <= 2;  //54 / 24 = 2
    16'b00110110_00011001 : OUT <= 2;  //54 / 25 = 2
    16'b00110110_00011010 : OUT <= 2;  //54 / 26 = 2
    16'b00110110_00011011 : OUT <= 2;  //54 / 27 = 2
    16'b00110110_00011100 : OUT <= 1;  //54 / 28 = 1
    16'b00110110_00011101 : OUT <= 1;  //54 / 29 = 1
    16'b00110110_00011110 : OUT <= 1;  //54 / 30 = 1
    16'b00110110_00011111 : OUT <= 1;  //54 / 31 = 1
    16'b00110110_00100000 : OUT <= 1;  //54 / 32 = 1
    16'b00110110_00100001 : OUT <= 1;  //54 / 33 = 1
    16'b00110110_00100010 : OUT <= 1;  //54 / 34 = 1
    16'b00110110_00100011 : OUT <= 1;  //54 / 35 = 1
    16'b00110110_00100100 : OUT <= 1;  //54 / 36 = 1
    16'b00110110_00100101 : OUT <= 1;  //54 / 37 = 1
    16'b00110110_00100110 : OUT <= 1;  //54 / 38 = 1
    16'b00110110_00100111 : OUT <= 1;  //54 / 39 = 1
    16'b00110110_00101000 : OUT <= 1;  //54 / 40 = 1
    16'b00110110_00101001 : OUT <= 1;  //54 / 41 = 1
    16'b00110110_00101010 : OUT <= 1;  //54 / 42 = 1
    16'b00110110_00101011 : OUT <= 1;  //54 / 43 = 1
    16'b00110110_00101100 : OUT <= 1;  //54 / 44 = 1
    16'b00110110_00101101 : OUT <= 1;  //54 / 45 = 1
    16'b00110110_00101110 : OUT <= 1;  //54 / 46 = 1
    16'b00110110_00101111 : OUT <= 1;  //54 / 47 = 1
    16'b00110110_00110000 : OUT <= 1;  //54 / 48 = 1
    16'b00110110_00110001 : OUT <= 1;  //54 / 49 = 1
    16'b00110110_00110010 : OUT <= 1;  //54 / 50 = 1
    16'b00110110_00110011 : OUT <= 1;  //54 / 51 = 1
    16'b00110110_00110100 : OUT <= 1;  //54 / 52 = 1
    16'b00110110_00110101 : OUT <= 1;  //54 / 53 = 1
    16'b00110110_00110110 : OUT <= 1;  //54 / 54 = 1
    16'b00110110_00110111 : OUT <= 0;  //54 / 55 = 0
    16'b00110110_00111000 : OUT <= 0;  //54 / 56 = 0
    16'b00110110_00111001 : OUT <= 0;  //54 / 57 = 0
    16'b00110110_00111010 : OUT <= 0;  //54 / 58 = 0
    16'b00110110_00111011 : OUT <= 0;  //54 / 59 = 0
    16'b00110110_00111100 : OUT <= 0;  //54 / 60 = 0
    16'b00110110_00111101 : OUT <= 0;  //54 / 61 = 0
    16'b00110110_00111110 : OUT <= 0;  //54 / 62 = 0
    16'b00110110_00111111 : OUT <= 0;  //54 / 63 = 0
    16'b00110110_01000000 : OUT <= 0;  //54 / 64 = 0
    16'b00110110_01000001 : OUT <= 0;  //54 / 65 = 0
    16'b00110110_01000010 : OUT <= 0;  //54 / 66 = 0
    16'b00110110_01000011 : OUT <= 0;  //54 / 67 = 0
    16'b00110110_01000100 : OUT <= 0;  //54 / 68 = 0
    16'b00110110_01000101 : OUT <= 0;  //54 / 69 = 0
    16'b00110110_01000110 : OUT <= 0;  //54 / 70 = 0
    16'b00110110_01000111 : OUT <= 0;  //54 / 71 = 0
    16'b00110110_01001000 : OUT <= 0;  //54 / 72 = 0
    16'b00110110_01001001 : OUT <= 0;  //54 / 73 = 0
    16'b00110110_01001010 : OUT <= 0;  //54 / 74 = 0
    16'b00110110_01001011 : OUT <= 0;  //54 / 75 = 0
    16'b00110110_01001100 : OUT <= 0;  //54 / 76 = 0
    16'b00110110_01001101 : OUT <= 0;  //54 / 77 = 0
    16'b00110110_01001110 : OUT <= 0;  //54 / 78 = 0
    16'b00110110_01001111 : OUT <= 0;  //54 / 79 = 0
    16'b00110110_01010000 : OUT <= 0;  //54 / 80 = 0
    16'b00110110_01010001 : OUT <= 0;  //54 / 81 = 0
    16'b00110110_01010010 : OUT <= 0;  //54 / 82 = 0
    16'b00110110_01010011 : OUT <= 0;  //54 / 83 = 0
    16'b00110110_01010100 : OUT <= 0;  //54 / 84 = 0
    16'b00110110_01010101 : OUT <= 0;  //54 / 85 = 0
    16'b00110110_01010110 : OUT <= 0;  //54 / 86 = 0
    16'b00110110_01010111 : OUT <= 0;  //54 / 87 = 0
    16'b00110110_01011000 : OUT <= 0;  //54 / 88 = 0
    16'b00110110_01011001 : OUT <= 0;  //54 / 89 = 0
    16'b00110110_01011010 : OUT <= 0;  //54 / 90 = 0
    16'b00110110_01011011 : OUT <= 0;  //54 / 91 = 0
    16'b00110110_01011100 : OUT <= 0;  //54 / 92 = 0
    16'b00110110_01011101 : OUT <= 0;  //54 / 93 = 0
    16'b00110110_01011110 : OUT <= 0;  //54 / 94 = 0
    16'b00110110_01011111 : OUT <= 0;  //54 / 95 = 0
    16'b00110110_01100000 : OUT <= 0;  //54 / 96 = 0
    16'b00110110_01100001 : OUT <= 0;  //54 / 97 = 0
    16'b00110110_01100010 : OUT <= 0;  //54 / 98 = 0
    16'b00110110_01100011 : OUT <= 0;  //54 / 99 = 0
    16'b00110110_01100100 : OUT <= 0;  //54 / 100 = 0
    16'b00110110_01100101 : OUT <= 0;  //54 / 101 = 0
    16'b00110110_01100110 : OUT <= 0;  //54 / 102 = 0
    16'b00110110_01100111 : OUT <= 0;  //54 / 103 = 0
    16'b00110110_01101000 : OUT <= 0;  //54 / 104 = 0
    16'b00110110_01101001 : OUT <= 0;  //54 / 105 = 0
    16'b00110110_01101010 : OUT <= 0;  //54 / 106 = 0
    16'b00110110_01101011 : OUT <= 0;  //54 / 107 = 0
    16'b00110110_01101100 : OUT <= 0;  //54 / 108 = 0
    16'b00110110_01101101 : OUT <= 0;  //54 / 109 = 0
    16'b00110110_01101110 : OUT <= 0;  //54 / 110 = 0
    16'b00110110_01101111 : OUT <= 0;  //54 / 111 = 0
    16'b00110110_01110000 : OUT <= 0;  //54 / 112 = 0
    16'b00110110_01110001 : OUT <= 0;  //54 / 113 = 0
    16'b00110110_01110010 : OUT <= 0;  //54 / 114 = 0
    16'b00110110_01110011 : OUT <= 0;  //54 / 115 = 0
    16'b00110110_01110100 : OUT <= 0;  //54 / 116 = 0
    16'b00110110_01110101 : OUT <= 0;  //54 / 117 = 0
    16'b00110110_01110110 : OUT <= 0;  //54 / 118 = 0
    16'b00110110_01110111 : OUT <= 0;  //54 / 119 = 0
    16'b00110110_01111000 : OUT <= 0;  //54 / 120 = 0
    16'b00110110_01111001 : OUT <= 0;  //54 / 121 = 0
    16'b00110110_01111010 : OUT <= 0;  //54 / 122 = 0
    16'b00110110_01111011 : OUT <= 0;  //54 / 123 = 0
    16'b00110110_01111100 : OUT <= 0;  //54 / 124 = 0
    16'b00110110_01111101 : OUT <= 0;  //54 / 125 = 0
    16'b00110110_01111110 : OUT <= 0;  //54 / 126 = 0
    16'b00110110_01111111 : OUT <= 0;  //54 / 127 = 0
    16'b00110110_10000000 : OUT <= 0;  //54 / 128 = 0
    16'b00110110_10000001 : OUT <= 0;  //54 / 129 = 0
    16'b00110110_10000010 : OUT <= 0;  //54 / 130 = 0
    16'b00110110_10000011 : OUT <= 0;  //54 / 131 = 0
    16'b00110110_10000100 : OUT <= 0;  //54 / 132 = 0
    16'b00110110_10000101 : OUT <= 0;  //54 / 133 = 0
    16'b00110110_10000110 : OUT <= 0;  //54 / 134 = 0
    16'b00110110_10000111 : OUT <= 0;  //54 / 135 = 0
    16'b00110110_10001000 : OUT <= 0;  //54 / 136 = 0
    16'b00110110_10001001 : OUT <= 0;  //54 / 137 = 0
    16'b00110110_10001010 : OUT <= 0;  //54 / 138 = 0
    16'b00110110_10001011 : OUT <= 0;  //54 / 139 = 0
    16'b00110110_10001100 : OUT <= 0;  //54 / 140 = 0
    16'b00110110_10001101 : OUT <= 0;  //54 / 141 = 0
    16'b00110110_10001110 : OUT <= 0;  //54 / 142 = 0
    16'b00110110_10001111 : OUT <= 0;  //54 / 143 = 0
    16'b00110110_10010000 : OUT <= 0;  //54 / 144 = 0
    16'b00110110_10010001 : OUT <= 0;  //54 / 145 = 0
    16'b00110110_10010010 : OUT <= 0;  //54 / 146 = 0
    16'b00110110_10010011 : OUT <= 0;  //54 / 147 = 0
    16'b00110110_10010100 : OUT <= 0;  //54 / 148 = 0
    16'b00110110_10010101 : OUT <= 0;  //54 / 149 = 0
    16'b00110110_10010110 : OUT <= 0;  //54 / 150 = 0
    16'b00110110_10010111 : OUT <= 0;  //54 / 151 = 0
    16'b00110110_10011000 : OUT <= 0;  //54 / 152 = 0
    16'b00110110_10011001 : OUT <= 0;  //54 / 153 = 0
    16'b00110110_10011010 : OUT <= 0;  //54 / 154 = 0
    16'b00110110_10011011 : OUT <= 0;  //54 / 155 = 0
    16'b00110110_10011100 : OUT <= 0;  //54 / 156 = 0
    16'b00110110_10011101 : OUT <= 0;  //54 / 157 = 0
    16'b00110110_10011110 : OUT <= 0;  //54 / 158 = 0
    16'b00110110_10011111 : OUT <= 0;  //54 / 159 = 0
    16'b00110110_10100000 : OUT <= 0;  //54 / 160 = 0
    16'b00110110_10100001 : OUT <= 0;  //54 / 161 = 0
    16'b00110110_10100010 : OUT <= 0;  //54 / 162 = 0
    16'b00110110_10100011 : OUT <= 0;  //54 / 163 = 0
    16'b00110110_10100100 : OUT <= 0;  //54 / 164 = 0
    16'b00110110_10100101 : OUT <= 0;  //54 / 165 = 0
    16'b00110110_10100110 : OUT <= 0;  //54 / 166 = 0
    16'b00110110_10100111 : OUT <= 0;  //54 / 167 = 0
    16'b00110110_10101000 : OUT <= 0;  //54 / 168 = 0
    16'b00110110_10101001 : OUT <= 0;  //54 / 169 = 0
    16'b00110110_10101010 : OUT <= 0;  //54 / 170 = 0
    16'b00110110_10101011 : OUT <= 0;  //54 / 171 = 0
    16'b00110110_10101100 : OUT <= 0;  //54 / 172 = 0
    16'b00110110_10101101 : OUT <= 0;  //54 / 173 = 0
    16'b00110110_10101110 : OUT <= 0;  //54 / 174 = 0
    16'b00110110_10101111 : OUT <= 0;  //54 / 175 = 0
    16'b00110110_10110000 : OUT <= 0;  //54 / 176 = 0
    16'b00110110_10110001 : OUT <= 0;  //54 / 177 = 0
    16'b00110110_10110010 : OUT <= 0;  //54 / 178 = 0
    16'b00110110_10110011 : OUT <= 0;  //54 / 179 = 0
    16'b00110110_10110100 : OUT <= 0;  //54 / 180 = 0
    16'b00110110_10110101 : OUT <= 0;  //54 / 181 = 0
    16'b00110110_10110110 : OUT <= 0;  //54 / 182 = 0
    16'b00110110_10110111 : OUT <= 0;  //54 / 183 = 0
    16'b00110110_10111000 : OUT <= 0;  //54 / 184 = 0
    16'b00110110_10111001 : OUT <= 0;  //54 / 185 = 0
    16'b00110110_10111010 : OUT <= 0;  //54 / 186 = 0
    16'b00110110_10111011 : OUT <= 0;  //54 / 187 = 0
    16'b00110110_10111100 : OUT <= 0;  //54 / 188 = 0
    16'b00110110_10111101 : OUT <= 0;  //54 / 189 = 0
    16'b00110110_10111110 : OUT <= 0;  //54 / 190 = 0
    16'b00110110_10111111 : OUT <= 0;  //54 / 191 = 0
    16'b00110110_11000000 : OUT <= 0;  //54 / 192 = 0
    16'b00110110_11000001 : OUT <= 0;  //54 / 193 = 0
    16'b00110110_11000010 : OUT <= 0;  //54 / 194 = 0
    16'b00110110_11000011 : OUT <= 0;  //54 / 195 = 0
    16'b00110110_11000100 : OUT <= 0;  //54 / 196 = 0
    16'b00110110_11000101 : OUT <= 0;  //54 / 197 = 0
    16'b00110110_11000110 : OUT <= 0;  //54 / 198 = 0
    16'b00110110_11000111 : OUT <= 0;  //54 / 199 = 0
    16'b00110110_11001000 : OUT <= 0;  //54 / 200 = 0
    16'b00110110_11001001 : OUT <= 0;  //54 / 201 = 0
    16'b00110110_11001010 : OUT <= 0;  //54 / 202 = 0
    16'b00110110_11001011 : OUT <= 0;  //54 / 203 = 0
    16'b00110110_11001100 : OUT <= 0;  //54 / 204 = 0
    16'b00110110_11001101 : OUT <= 0;  //54 / 205 = 0
    16'b00110110_11001110 : OUT <= 0;  //54 / 206 = 0
    16'b00110110_11001111 : OUT <= 0;  //54 / 207 = 0
    16'b00110110_11010000 : OUT <= 0;  //54 / 208 = 0
    16'b00110110_11010001 : OUT <= 0;  //54 / 209 = 0
    16'b00110110_11010010 : OUT <= 0;  //54 / 210 = 0
    16'b00110110_11010011 : OUT <= 0;  //54 / 211 = 0
    16'b00110110_11010100 : OUT <= 0;  //54 / 212 = 0
    16'b00110110_11010101 : OUT <= 0;  //54 / 213 = 0
    16'b00110110_11010110 : OUT <= 0;  //54 / 214 = 0
    16'b00110110_11010111 : OUT <= 0;  //54 / 215 = 0
    16'b00110110_11011000 : OUT <= 0;  //54 / 216 = 0
    16'b00110110_11011001 : OUT <= 0;  //54 / 217 = 0
    16'b00110110_11011010 : OUT <= 0;  //54 / 218 = 0
    16'b00110110_11011011 : OUT <= 0;  //54 / 219 = 0
    16'b00110110_11011100 : OUT <= 0;  //54 / 220 = 0
    16'b00110110_11011101 : OUT <= 0;  //54 / 221 = 0
    16'b00110110_11011110 : OUT <= 0;  //54 / 222 = 0
    16'b00110110_11011111 : OUT <= 0;  //54 / 223 = 0
    16'b00110110_11100000 : OUT <= 0;  //54 / 224 = 0
    16'b00110110_11100001 : OUT <= 0;  //54 / 225 = 0
    16'b00110110_11100010 : OUT <= 0;  //54 / 226 = 0
    16'b00110110_11100011 : OUT <= 0;  //54 / 227 = 0
    16'b00110110_11100100 : OUT <= 0;  //54 / 228 = 0
    16'b00110110_11100101 : OUT <= 0;  //54 / 229 = 0
    16'b00110110_11100110 : OUT <= 0;  //54 / 230 = 0
    16'b00110110_11100111 : OUT <= 0;  //54 / 231 = 0
    16'b00110110_11101000 : OUT <= 0;  //54 / 232 = 0
    16'b00110110_11101001 : OUT <= 0;  //54 / 233 = 0
    16'b00110110_11101010 : OUT <= 0;  //54 / 234 = 0
    16'b00110110_11101011 : OUT <= 0;  //54 / 235 = 0
    16'b00110110_11101100 : OUT <= 0;  //54 / 236 = 0
    16'b00110110_11101101 : OUT <= 0;  //54 / 237 = 0
    16'b00110110_11101110 : OUT <= 0;  //54 / 238 = 0
    16'b00110110_11101111 : OUT <= 0;  //54 / 239 = 0
    16'b00110110_11110000 : OUT <= 0;  //54 / 240 = 0
    16'b00110110_11110001 : OUT <= 0;  //54 / 241 = 0
    16'b00110110_11110010 : OUT <= 0;  //54 / 242 = 0
    16'b00110110_11110011 : OUT <= 0;  //54 / 243 = 0
    16'b00110110_11110100 : OUT <= 0;  //54 / 244 = 0
    16'b00110110_11110101 : OUT <= 0;  //54 / 245 = 0
    16'b00110110_11110110 : OUT <= 0;  //54 / 246 = 0
    16'b00110110_11110111 : OUT <= 0;  //54 / 247 = 0
    16'b00110110_11111000 : OUT <= 0;  //54 / 248 = 0
    16'b00110110_11111001 : OUT <= 0;  //54 / 249 = 0
    16'b00110110_11111010 : OUT <= 0;  //54 / 250 = 0
    16'b00110110_11111011 : OUT <= 0;  //54 / 251 = 0
    16'b00110110_11111100 : OUT <= 0;  //54 / 252 = 0
    16'b00110110_11111101 : OUT <= 0;  //54 / 253 = 0
    16'b00110110_11111110 : OUT <= 0;  //54 / 254 = 0
    16'b00110110_11111111 : OUT <= 0;  //54 / 255 = 0
    16'b00110111_00000000 : OUT <= 0;  //55 / 0 = 0
    16'b00110111_00000001 : OUT <= 55;  //55 / 1 = 55
    16'b00110111_00000010 : OUT <= 27;  //55 / 2 = 27
    16'b00110111_00000011 : OUT <= 18;  //55 / 3 = 18
    16'b00110111_00000100 : OUT <= 13;  //55 / 4 = 13
    16'b00110111_00000101 : OUT <= 11;  //55 / 5 = 11
    16'b00110111_00000110 : OUT <= 9;  //55 / 6 = 9
    16'b00110111_00000111 : OUT <= 7;  //55 / 7 = 7
    16'b00110111_00001000 : OUT <= 6;  //55 / 8 = 6
    16'b00110111_00001001 : OUT <= 6;  //55 / 9 = 6
    16'b00110111_00001010 : OUT <= 5;  //55 / 10 = 5
    16'b00110111_00001011 : OUT <= 5;  //55 / 11 = 5
    16'b00110111_00001100 : OUT <= 4;  //55 / 12 = 4
    16'b00110111_00001101 : OUT <= 4;  //55 / 13 = 4
    16'b00110111_00001110 : OUT <= 3;  //55 / 14 = 3
    16'b00110111_00001111 : OUT <= 3;  //55 / 15 = 3
    16'b00110111_00010000 : OUT <= 3;  //55 / 16 = 3
    16'b00110111_00010001 : OUT <= 3;  //55 / 17 = 3
    16'b00110111_00010010 : OUT <= 3;  //55 / 18 = 3
    16'b00110111_00010011 : OUT <= 2;  //55 / 19 = 2
    16'b00110111_00010100 : OUT <= 2;  //55 / 20 = 2
    16'b00110111_00010101 : OUT <= 2;  //55 / 21 = 2
    16'b00110111_00010110 : OUT <= 2;  //55 / 22 = 2
    16'b00110111_00010111 : OUT <= 2;  //55 / 23 = 2
    16'b00110111_00011000 : OUT <= 2;  //55 / 24 = 2
    16'b00110111_00011001 : OUT <= 2;  //55 / 25 = 2
    16'b00110111_00011010 : OUT <= 2;  //55 / 26 = 2
    16'b00110111_00011011 : OUT <= 2;  //55 / 27 = 2
    16'b00110111_00011100 : OUT <= 1;  //55 / 28 = 1
    16'b00110111_00011101 : OUT <= 1;  //55 / 29 = 1
    16'b00110111_00011110 : OUT <= 1;  //55 / 30 = 1
    16'b00110111_00011111 : OUT <= 1;  //55 / 31 = 1
    16'b00110111_00100000 : OUT <= 1;  //55 / 32 = 1
    16'b00110111_00100001 : OUT <= 1;  //55 / 33 = 1
    16'b00110111_00100010 : OUT <= 1;  //55 / 34 = 1
    16'b00110111_00100011 : OUT <= 1;  //55 / 35 = 1
    16'b00110111_00100100 : OUT <= 1;  //55 / 36 = 1
    16'b00110111_00100101 : OUT <= 1;  //55 / 37 = 1
    16'b00110111_00100110 : OUT <= 1;  //55 / 38 = 1
    16'b00110111_00100111 : OUT <= 1;  //55 / 39 = 1
    16'b00110111_00101000 : OUT <= 1;  //55 / 40 = 1
    16'b00110111_00101001 : OUT <= 1;  //55 / 41 = 1
    16'b00110111_00101010 : OUT <= 1;  //55 / 42 = 1
    16'b00110111_00101011 : OUT <= 1;  //55 / 43 = 1
    16'b00110111_00101100 : OUT <= 1;  //55 / 44 = 1
    16'b00110111_00101101 : OUT <= 1;  //55 / 45 = 1
    16'b00110111_00101110 : OUT <= 1;  //55 / 46 = 1
    16'b00110111_00101111 : OUT <= 1;  //55 / 47 = 1
    16'b00110111_00110000 : OUT <= 1;  //55 / 48 = 1
    16'b00110111_00110001 : OUT <= 1;  //55 / 49 = 1
    16'b00110111_00110010 : OUT <= 1;  //55 / 50 = 1
    16'b00110111_00110011 : OUT <= 1;  //55 / 51 = 1
    16'b00110111_00110100 : OUT <= 1;  //55 / 52 = 1
    16'b00110111_00110101 : OUT <= 1;  //55 / 53 = 1
    16'b00110111_00110110 : OUT <= 1;  //55 / 54 = 1
    16'b00110111_00110111 : OUT <= 1;  //55 / 55 = 1
    16'b00110111_00111000 : OUT <= 0;  //55 / 56 = 0
    16'b00110111_00111001 : OUT <= 0;  //55 / 57 = 0
    16'b00110111_00111010 : OUT <= 0;  //55 / 58 = 0
    16'b00110111_00111011 : OUT <= 0;  //55 / 59 = 0
    16'b00110111_00111100 : OUT <= 0;  //55 / 60 = 0
    16'b00110111_00111101 : OUT <= 0;  //55 / 61 = 0
    16'b00110111_00111110 : OUT <= 0;  //55 / 62 = 0
    16'b00110111_00111111 : OUT <= 0;  //55 / 63 = 0
    16'b00110111_01000000 : OUT <= 0;  //55 / 64 = 0
    16'b00110111_01000001 : OUT <= 0;  //55 / 65 = 0
    16'b00110111_01000010 : OUT <= 0;  //55 / 66 = 0
    16'b00110111_01000011 : OUT <= 0;  //55 / 67 = 0
    16'b00110111_01000100 : OUT <= 0;  //55 / 68 = 0
    16'b00110111_01000101 : OUT <= 0;  //55 / 69 = 0
    16'b00110111_01000110 : OUT <= 0;  //55 / 70 = 0
    16'b00110111_01000111 : OUT <= 0;  //55 / 71 = 0
    16'b00110111_01001000 : OUT <= 0;  //55 / 72 = 0
    16'b00110111_01001001 : OUT <= 0;  //55 / 73 = 0
    16'b00110111_01001010 : OUT <= 0;  //55 / 74 = 0
    16'b00110111_01001011 : OUT <= 0;  //55 / 75 = 0
    16'b00110111_01001100 : OUT <= 0;  //55 / 76 = 0
    16'b00110111_01001101 : OUT <= 0;  //55 / 77 = 0
    16'b00110111_01001110 : OUT <= 0;  //55 / 78 = 0
    16'b00110111_01001111 : OUT <= 0;  //55 / 79 = 0
    16'b00110111_01010000 : OUT <= 0;  //55 / 80 = 0
    16'b00110111_01010001 : OUT <= 0;  //55 / 81 = 0
    16'b00110111_01010010 : OUT <= 0;  //55 / 82 = 0
    16'b00110111_01010011 : OUT <= 0;  //55 / 83 = 0
    16'b00110111_01010100 : OUT <= 0;  //55 / 84 = 0
    16'b00110111_01010101 : OUT <= 0;  //55 / 85 = 0
    16'b00110111_01010110 : OUT <= 0;  //55 / 86 = 0
    16'b00110111_01010111 : OUT <= 0;  //55 / 87 = 0
    16'b00110111_01011000 : OUT <= 0;  //55 / 88 = 0
    16'b00110111_01011001 : OUT <= 0;  //55 / 89 = 0
    16'b00110111_01011010 : OUT <= 0;  //55 / 90 = 0
    16'b00110111_01011011 : OUT <= 0;  //55 / 91 = 0
    16'b00110111_01011100 : OUT <= 0;  //55 / 92 = 0
    16'b00110111_01011101 : OUT <= 0;  //55 / 93 = 0
    16'b00110111_01011110 : OUT <= 0;  //55 / 94 = 0
    16'b00110111_01011111 : OUT <= 0;  //55 / 95 = 0
    16'b00110111_01100000 : OUT <= 0;  //55 / 96 = 0
    16'b00110111_01100001 : OUT <= 0;  //55 / 97 = 0
    16'b00110111_01100010 : OUT <= 0;  //55 / 98 = 0
    16'b00110111_01100011 : OUT <= 0;  //55 / 99 = 0
    16'b00110111_01100100 : OUT <= 0;  //55 / 100 = 0
    16'b00110111_01100101 : OUT <= 0;  //55 / 101 = 0
    16'b00110111_01100110 : OUT <= 0;  //55 / 102 = 0
    16'b00110111_01100111 : OUT <= 0;  //55 / 103 = 0
    16'b00110111_01101000 : OUT <= 0;  //55 / 104 = 0
    16'b00110111_01101001 : OUT <= 0;  //55 / 105 = 0
    16'b00110111_01101010 : OUT <= 0;  //55 / 106 = 0
    16'b00110111_01101011 : OUT <= 0;  //55 / 107 = 0
    16'b00110111_01101100 : OUT <= 0;  //55 / 108 = 0
    16'b00110111_01101101 : OUT <= 0;  //55 / 109 = 0
    16'b00110111_01101110 : OUT <= 0;  //55 / 110 = 0
    16'b00110111_01101111 : OUT <= 0;  //55 / 111 = 0
    16'b00110111_01110000 : OUT <= 0;  //55 / 112 = 0
    16'b00110111_01110001 : OUT <= 0;  //55 / 113 = 0
    16'b00110111_01110010 : OUT <= 0;  //55 / 114 = 0
    16'b00110111_01110011 : OUT <= 0;  //55 / 115 = 0
    16'b00110111_01110100 : OUT <= 0;  //55 / 116 = 0
    16'b00110111_01110101 : OUT <= 0;  //55 / 117 = 0
    16'b00110111_01110110 : OUT <= 0;  //55 / 118 = 0
    16'b00110111_01110111 : OUT <= 0;  //55 / 119 = 0
    16'b00110111_01111000 : OUT <= 0;  //55 / 120 = 0
    16'b00110111_01111001 : OUT <= 0;  //55 / 121 = 0
    16'b00110111_01111010 : OUT <= 0;  //55 / 122 = 0
    16'b00110111_01111011 : OUT <= 0;  //55 / 123 = 0
    16'b00110111_01111100 : OUT <= 0;  //55 / 124 = 0
    16'b00110111_01111101 : OUT <= 0;  //55 / 125 = 0
    16'b00110111_01111110 : OUT <= 0;  //55 / 126 = 0
    16'b00110111_01111111 : OUT <= 0;  //55 / 127 = 0
    16'b00110111_10000000 : OUT <= 0;  //55 / 128 = 0
    16'b00110111_10000001 : OUT <= 0;  //55 / 129 = 0
    16'b00110111_10000010 : OUT <= 0;  //55 / 130 = 0
    16'b00110111_10000011 : OUT <= 0;  //55 / 131 = 0
    16'b00110111_10000100 : OUT <= 0;  //55 / 132 = 0
    16'b00110111_10000101 : OUT <= 0;  //55 / 133 = 0
    16'b00110111_10000110 : OUT <= 0;  //55 / 134 = 0
    16'b00110111_10000111 : OUT <= 0;  //55 / 135 = 0
    16'b00110111_10001000 : OUT <= 0;  //55 / 136 = 0
    16'b00110111_10001001 : OUT <= 0;  //55 / 137 = 0
    16'b00110111_10001010 : OUT <= 0;  //55 / 138 = 0
    16'b00110111_10001011 : OUT <= 0;  //55 / 139 = 0
    16'b00110111_10001100 : OUT <= 0;  //55 / 140 = 0
    16'b00110111_10001101 : OUT <= 0;  //55 / 141 = 0
    16'b00110111_10001110 : OUT <= 0;  //55 / 142 = 0
    16'b00110111_10001111 : OUT <= 0;  //55 / 143 = 0
    16'b00110111_10010000 : OUT <= 0;  //55 / 144 = 0
    16'b00110111_10010001 : OUT <= 0;  //55 / 145 = 0
    16'b00110111_10010010 : OUT <= 0;  //55 / 146 = 0
    16'b00110111_10010011 : OUT <= 0;  //55 / 147 = 0
    16'b00110111_10010100 : OUT <= 0;  //55 / 148 = 0
    16'b00110111_10010101 : OUT <= 0;  //55 / 149 = 0
    16'b00110111_10010110 : OUT <= 0;  //55 / 150 = 0
    16'b00110111_10010111 : OUT <= 0;  //55 / 151 = 0
    16'b00110111_10011000 : OUT <= 0;  //55 / 152 = 0
    16'b00110111_10011001 : OUT <= 0;  //55 / 153 = 0
    16'b00110111_10011010 : OUT <= 0;  //55 / 154 = 0
    16'b00110111_10011011 : OUT <= 0;  //55 / 155 = 0
    16'b00110111_10011100 : OUT <= 0;  //55 / 156 = 0
    16'b00110111_10011101 : OUT <= 0;  //55 / 157 = 0
    16'b00110111_10011110 : OUT <= 0;  //55 / 158 = 0
    16'b00110111_10011111 : OUT <= 0;  //55 / 159 = 0
    16'b00110111_10100000 : OUT <= 0;  //55 / 160 = 0
    16'b00110111_10100001 : OUT <= 0;  //55 / 161 = 0
    16'b00110111_10100010 : OUT <= 0;  //55 / 162 = 0
    16'b00110111_10100011 : OUT <= 0;  //55 / 163 = 0
    16'b00110111_10100100 : OUT <= 0;  //55 / 164 = 0
    16'b00110111_10100101 : OUT <= 0;  //55 / 165 = 0
    16'b00110111_10100110 : OUT <= 0;  //55 / 166 = 0
    16'b00110111_10100111 : OUT <= 0;  //55 / 167 = 0
    16'b00110111_10101000 : OUT <= 0;  //55 / 168 = 0
    16'b00110111_10101001 : OUT <= 0;  //55 / 169 = 0
    16'b00110111_10101010 : OUT <= 0;  //55 / 170 = 0
    16'b00110111_10101011 : OUT <= 0;  //55 / 171 = 0
    16'b00110111_10101100 : OUT <= 0;  //55 / 172 = 0
    16'b00110111_10101101 : OUT <= 0;  //55 / 173 = 0
    16'b00110111_10101110 : OUT <= 0;  //55 / 174 = 0
    16'b00110111_10101111 : OUT <= 0;  //55 / 175 = 0
    16'b00110111_10110000 : OUT <= 0;  //55 / 176 = 0
    16'b00110111_10110001 : OUT <= 0;  //55 / 177 = 0
    16'b00110111_10110010 : OUT <= 0;  //55 / 178 = 0
    16'b00110111_10110011 : OUT <= 0;  //55 / 179 = 0
    16'b00110111_10110100 : OUT <= 0;  //55 / 180 = 0
    16'b00110111_10110101 : OUT <= 0;  //55 / 181 = 0
    16'b00110111_10110110 : OUT <= 0;  //55 / 182 = 0
    16'b00110111_10110111 : OUT <= 0;  //55 / 183 = 0
    16'b00110111_10111000 : OUT <= 0;  //55 / 184 = 0
    16'b00110111_10111001 : OUT <= 0;  //55 / 185 = 0
    16'b00110111_10111010 : OUT <= 0;  //55 / 186 = 0
    16'b00110111_10111011 : OUT <= 0;  //55 / 187 = 0
    16'b00110111_10111100 : OUT <= 0;  //55 / 188 = 0
    16'b00110111_10111101 : OUT <= 0;  //55 / 189 = 0
    16'b00110111_10111110 : OUT <= 0;  //55 / 190 = 0
    16'b00110111_10111111 : OUT <= 0;  //55 / 191 = 0
    16'b00110111_11000000 : OUT <= 0;  //55 / 192 = 0
    16'b00110111_11000001 : OUT <= 0;  //55 / 193 = 0
    16'b00110111_11000010 : OUT <= 0;  //55 / 194 = 0
    16'b00110111_11000011 : OUT <= 0;  //55 / 195 = 0
    16'b00110111_11000100 : OUT <= 0;  //55 / 196 = 0
    16'b00110111_11000101 : OUT <= 0;  //55 / 197 = 0
    16'b00110111_11000110 : OUT <= 0;  //55 / 198 = 0
    16'b00110111_11000111 : OUT <= 0;  //55 / 199 = 0
    16'b00110111_11001000 : OUT <= 0;  //55 / 200 = 0
    16'b00110111_11001001 : OUT <= 0;  //55 / 201 = 0
    16'b00110111_11001010 : OUT <= 0;  //55 / 202 = 0
    16'b00110111_11001011 : OUT <= 0;  //55 / 203 = 0
    16'b00110111_11001100 : OUT <= 0;  //55 / 204 = 0
    16'b00110111_11001101 : OUT <= 0;  //55 / 205 = 0
    16'b00110111_11001110 : OUT <= 0;  //55 / 206 = 0
    16'b00110111_11001111 : OUT <= 0;  //55 / 207 = 0
    16'b00110111_11010000 : OUT <= 0;  //55 / 208 = 0
    16'b00110111_11010001 : OUT <= 0;  //55 / 209 = 0
    16'b00110111_11010010 : OUT <= 0;  //55 / 210 = 0
    16'b00110111_11010011 : OUT <= 0;  //55 / 211 = 0
    16'b00110111_11010100 : OUT <= 0;  //55 / 212 = 0
    16'b00110111_11010101 : OUT <= 0;  //55 / 213 = 0
    16'b00110111_11010110 : OUT <= 0;  //55 / 214 = 0
    16'b00110111_11010111 : OUT <= 0;  //55 / 215 = 0
    16'b00110111_11011000 : OUT <= 0;  //55 / 216 = 0
    16'b00110111_11011001 : OUT <= 0;  //55 / 217 = 0
    16'b00110111_11011010 : OUT <= 0;  //55 / 218 = 0
    16'b00110111_11011011 : OUT <= 0;  //55 / 219 = 0
    16'b00110111_11011100 : OUT <= 0;  //55 / 220 = 0
    16'b00110111_11011101 : OUT <= 0;  //55 / 221 = 0
    16'b00110111_11011110 : OUT <= 0;  //55 / 222 = 0
    16'b00110111_11011111 : OUT <= 0;  //55 / 223 = 0
    16'b00110111_11100000 : OUT <= 0;  //55 / 224 = 0
    16'b00110111_11100001 : OUT <= 0;  //55 / 225 = 0
    16'b00110111_11100010 : OUT <= 0;  //55 / 226 = 0
    16'b00110111_11100011 : OUT <= 0;  //55 / 227 = 0
    16'b00110111_11100100 : OUT <= 0;  //55 / 228 = 0
    16'b00110111_11100101 : OUT <= 0;  //55 / 229 = 0
    16'b00110111_11100110 : OUT <= 0;  //55 / 230 = 0
    16'b00110111_11100111 : OUT <= 0;  //55 / 231 = 0
    16'b00110111_11101000 : OUT <= 0;  //55 / 232 = 0
    16'b00110111_11101001 : OUT <= 0;  //55 / 233 = 0
    16'b00110111_11101010 : OUT <= 0;  //55 / 234 = 0
    16'b00110111_11101011 : OUT <= 0;  //55 / 235 = 0
    16'b00110111_11101100 : OUT <= 0;  //55 / 236 = 0
    16'b00110111_11101101 : OUT <= 0;  //55 / 237 = 0
    16'b00110111_11101110 : OUT <= 0;  //55 / 238 = 0
    16'b00110111_11101111 : OUT <= 0;  //55 / 239 = 0
    16'b00110111_11110000 : OUT <= 0;  //55 / 240 = 0
    16'b00110111_11110001 : OUT <= 0;  //55 / 241 = 0
    16'b00110111_11110010 : OUT <= 0;  //55 / 242 = 0
    16'b00110111_11110011 : OUT <= 0;  //55 / 243 = 0
    16'b00110111_11110100 : OUT <= 0;  //55 / 244 = 0
    16'b00110111_11110101 : OUT <= 0;  //55 / 245 = 0
    16'b00110111_11110110 : OUT <= 0;  //55 / 246 = 0
    16'b00110111_11110111 : OUT <= 0;  //55 / 247 = 0
    16'b00110111_11111000 : OUT <= 0;  //55 / 248 = 0
    16'b00110111_11111001 : OUT <= 0;  //55 / 249 = 0
    16'b00110111_11111010 : OUT <= 0;  //55 / 250 = 0
    16'b00110111_11111011 : OUT <= 0;  //55 / 251 = 0
    16'b00110111_11111100 : OUT <= 0;  //55 / 252 = 0
    16'b00110111_11111101 : OUT <= 0;  //55 / 253 = 0
    16'b00110111_11111110 : OUT <= 0;  //55 / 254 = 0
    16'b00110111_11111111 : OUT <= 0;  //55 / 255 = 0
    16'b00111000_00000000 : OUT <= 0;  //56 / 0 = 0
    16'b00111000_00000001 : OUT <= 56;  //56 / 1 = 56
    16'b00111000_00000010 : OUT <= 28;  //56 / 2 = 28
    16'b00111000_00000011 : OUT <= 18;  //56 / 3 = 18
    16'b00111000_00000100 : OUT <= 14;  //56 / 4 = 14
    16'b00111000_00000101 : OUT <= 11;  //56 / 5 = 11
    16'b00111000_00000110 : OUT <= 9;  //56 / 6 = 9
    16'b00111000_00000111 : OUT <= 8;  //56 / 7 = 8
    16'b00111000_00001000 : OUT <= 7;  //56 / 8 = 7
    16'b00111000_00001001 : OUT <= 6;  //56 / 9 = 6
    16'b00111000_00001010 : OUT <= 5;  //56 / 10 = 5
    16'b00111000_00001011 : OUT <= 5;  //56 / 11 = 5
    16'b00111000_00001100 : OUT <= 4;  //56 / 12 = 4
    16'b00111000_00001101 : OUT <= 4;  //56 / 13 = 4
    16'b00111000_00001110 : OUT <= 4;  //56 / 14 = 4
    16'b00111000_00001111 : OUT <= 3;  //56 / 15 = 3
    16'b00111000_00010000 : OUT <= 3;  //56 / 16 = 3
    16'b00111000_00010001 : OUT <= 3;  //56 / 17 = 3
    16'b00111000_00010010 : OUT <= 3;  //56 / 18 = 3
    16'b00111000_00010011 : OUT <= 2;  //56 / 19 = 2
    16'b00111000_00010100 : OUT <= 2;  //56 / 20 = 2
    16'b00111000_00010101 : OUT <= 2;  //56 / 21 = 2
    16'b00111000_00010110 : OUT <= 2;  //56 / 22 = 2
    16'b00111000_00010111 : OUT <= 2;  //56 / 23 = 2
    16'b00111000_00011000 : OUT <= 2;  //56 / 24 = 2
    16'b00111000_00011001 : OUT <= 2;  //56 / 25 = 2
    16'b00111000_00011010 : OUT <= 2;  //56 / 26 = 2
    16'b00111000_00011011 : OUT <= 2;  //56 / 27 = 2
    16'b00111000_00011100 : OUT <= 2;  //56 / 28 = 2
    16'b00111000_00011101 : OUT <= 1;  //56 / 29 = 1
    16'b00111000_00011110 : OUT <= 1;  //56 / 30 = 1
    16'b00111000_00011111 : OUT <= 1;  //56 / 31 = 1
    16'b00111000_00100000 : OUT <= 1;  //56 / 32 = 1
    16'b00111000_00100001 : OUT <= 1;  //56 / 33 = 1
    16'b00111000_00100010 : OUT <= 1;  //56 / 34 = 1
    16'b00111000_00100011 : OUT <= 1;  //56 / 35 = 1
    16'b00111000_00100100 : OUT <= 1;  //56 / 36 = 1
    16'b00111000_00100101 : OUT <= 1;  //56 / 37 = 1
    16'b00111000_00100110 : OUT <= 1;  //56 / 38 = 1
    16'b00111000_00100111 : OUT <= 1;  //56 / 39 = 1
    16'b00111000_00101000 : OUT <= 1;  //56 / 40 = 1
    16'b00111000_00101001 : OUT <= 1;  //56 / 41 = 1
    16'b00111000_00101010 : OUT <= 1;  //56 / 42 = 1
    16'b00111000_00101011 : OUT <= 1;  //56 / 43 = 1
    16'b00111000_00101100 : OUT <= 1;  //56 / 44 = 1
    16'b00111000_00101101 : OUT <= 1;  //56 / 45 = 1
    16'b00111000_00101110 : OUT <= 1;  //56 / 46 = 1
    16'b00111000_00101111 : OUT <= 1;  //56 / 47 = 1
    16'b00111000_00110000 : OUT <= 1;  //56 / 48 = 1
    16'b00111000_00110001 : OUT <= 1;  //56 / 49 = 1
    16'b00111000_00110010 : OUT <= 1;  //56 / 50 = 1
    16'b00111000_00110011 : OUT <= 1;  //56 / 51 = 1
    16'b00111000_00110100 : OUT <= 1;  //56 / 52 = 1
    16'b00111000_00110101 : OUT <= 1;  //56 / 53 = 1
    16'b00111000_00110110 : OUT <= 1;  //56 / 54 = 1
    16'b00111000_00110111 : OUT <= 1;  //56 / 55 = 1
    16'b00111000_00111000 : OUT <= 1;  //56 / 56 = 1
    16'b00111000_00111001 : OUT <= 0;  //56 / 57 = 0
    16'b00111000_00111010 : OUT <= 0;  //56 / 58 = 0
    16'b00111000_00111011 : OUT <= 0;  //56 / 59 = 0
    16'b00111000_00111100 : OUT <= 0;  //56 / 60 = 0
    16'b00111000_00111101 : OUT <= 0;  //56 / 61 = 0
    16'b00111000_00111110 : OUT <= 0;  //56 / 62 = 0
    16'b00111000_00111111 : OUT <= 0;  //56 / 63 = 0
    16'b00111000_01000000 : OUT <= 0;  //56 / 64 = 0
    16'b00111000_01000001 : OUT <= 0;  //56 / 65 = 0
    16'b00111000_01000010 : OUT <= 0;  //56 / 66 = 0
    16'b00111000_01000011 : OUT <= 0;  //56 / 67 = 0
    16'b00111000_01000100 : OUT <= 0;  //56 / 68 = 0
    16'b00111000_01000101 : OUT <= 0;  //56 / 69 = 0
    16'b00111000_01000110 : OUT <= 0;  //56 / 70 = 0
    16'b00111000_01000111 : OUT <= 0;  //56 / 71 = 0
    16'b00111000_01001000 : OUT <= 0;  //56 / 72 = 0
    16'b00111000_01001001 : OUT <= 0;  //56 / 73 = 0
    16'b00111000_01001010 : OUT <= 0;  //56 / 74 = 0
    16'b00111000_01001011 : OUT <= 0;  //56 / 75 = 0
    16'b00111000_01001100 : OUT <= 0;  //56 / 76 = 0
    16'b00111000_01001101 : OUT <= 0;  //56 / 77 = 0
    16'b00111000_01001110 : OUT <= 0;  //56 / 78 = 0
    16'b00111000_01001111 : OUT <= 0;  //56 / 79 = 0
    16'b00111000_01010000 : OUT <= 0;  //56 / 80 = 0
    16'b00111000_01010001 : OUT <= 0;  //56 / 81 = 0
    16'b00111000_01010010 : OUT <= 0;  //56 / 82 = 0
    16'b00111000_01010011 : OUT <= 0;  //56 / 83 = 0
    16'b00111000_01010100 : OUT <= 0;  //56 / 84 = 0
    16'b00111000_01010101 : OUT <= 0;  //56 / 85 = 0
    16'b00111000_01010110 : OUT <= 0;  //56 / 86 = 0
    16'b00111000_01010111 : OUT <= 0;  //56 / 87 = 0
    16'b00111000_01011000 : OUT <= 0;  //56 / 88 = 0
    16'b00111000_01011001 : OUT <= 0;  //56 / 89 = 0
    16'b00111000_01011010 : OUT <= 0;  //56 / 90 = 0
    16'b00111000_01011011 : OUT <= 0;  //56 / 91 = 0
    16'b00111000_01011100 : OUT <= 0;  //56 / 92 = 0
    16'b00111000_01011101 : OUT <= 0;  //56 / 93 = 0
    16'b00111000_01011110 : OUT <= 0;  //56 / 94 = 0
    16'b00111000_01011111 : OUT <= 0;  //56 / 95 = 0
    16'b00111000_01100000 : OUT <= 0;  //56 / 96 = 0
    16'b00111000_01100001 : OUT <= 0;  //56 / 97 = 0
    16'b00111000_01100010 : OUT <= 0;  //56 / 98 = 0
    16'b00111000_01100011 : OUT <= 0;  //56 / 99 = 0
    16'b00111000_01100100 : OUT <= 0;  //56 / 100 = 0
    16'b00111000_01100101 : OUT <= 0;  //56 / 101 = 0
    16'b00111000_01100110 : OUT <= 0;  //56 / 102 = 0
    16'b00111000_01100111 : OUT <= 0;  //56 / 103 = 0
    16'b00111000_01101000 : OUT <= 0;  //56 / 104 = 0
    16'b00111000_01101001 : OUT <= 0;  //56 / 105 = 0
    16'b00111000_01101010 : OUT <= 0;  //56 / 106 = 0
    16'b00111000_01101011 : OUT <= 0;  //56 / 107 = 0
    16'b00111000_01101100 : OUT <= 0;  //56 / 108 = 0
    16'b00111000_01101101 : OUT <= 0;  //56 / 109 = 0
    16'b00111000_01101110 : OUT <= 0;  //56 / 110 = 0
    16'b00111000_01101111 : OUT <= 0;  //56 / 111 = 0
    16'b00111000_01110000 : OUT <= 0;  //56 / 112 = 0
    16'b00111000_01110001 : OUT <= 0;  //56 / 113 = 0
    16'b00111000_01110010 : OUT <= 0;  //56 / 114 = 0
    16'b00111000_01110011 : OUT <= 0;  //56 / 115 = 0
    16'b00111000_01110100 : OUT <= 0;  //56 / 116 = 0
    16'b00111000_01110101 : OUT <= 0;  //56 / 117 = 0
    16'b00111000_01110110 : OUT <= 0;  //56 / 118 = 0
    16'b00111000_01110111 : OUT <= 0;  //56 / 119 = 0
    16'b00111000_01111000 : OUT <= 0;  //56 / 120 = 0
    16'b00111000_01111001 : OUT <= 0;  //56 / 121 = 0
    16'b00111000_01111010 : OUT <= 0;  //56 / 122 = 0
    16'b00111000_01111011 : OUT <= 0;  //56 / 123 = 0
    16'b00111000_01111100 : OUT <= 0;  //56 / 124 = 0
    16'b00111000_01111101 : OUT <= 0;  //56 / 125 = 0
    16'b00111000_01111110 : OUT <= 0;  //56 / 126 = 0
    16'b00111000_01111111 : OUT <= 0;  //56 / 127 = 0
    16'b00111000_10000000 : OUT <= 0;  //56 / 128 = 0
    16'b00111000_10000001 : OUT <= 0;  //56 / 129 = 0
    16'b00111000_10000010 : OUT <= 0;  //56 / 130 = 0
    16'b00111000_10000011 : OUT <= 0;  //56 / 131 = 0
    16'b00111000_10000100 : OUT <= 0;  //56 / 132 = 0
    16'b00111000_10000101 : OUT <= 0;  //56 / 133 = 0
    16'b00111000_10000110 : OUT <= 0;  //56 / 134 = 0
    16'b00111000_10000111 : OUT <= 0;  //56 / 135 = 0
    16'b00111000_10001000 : OUT <= 0;  //56 / 136 = 0
    16'b00111000_10001001 : OUT <= 0;  //56 / 137 = 0
    16'b00111000_10001010 : OUT <= 0;  //56 / 138 = 0
    16'b00111000_10001011 : OUT <= 0;  //56 / 139 = 0
    16'b00111000_10001100 : OUT <= 0;  //56 / 140 = 0
    16'b00111000_10001101 : OUT <= 0;  //56 / 141 = 0
    16'b00111000_10001110 : OUT <= 0;  //56 / 142 = 0
    16'b00111000_10001111 : OUT <= 0;  //56 / 143 = 0
    16'b00111000_10010000 : OUT <= 0;  //56 / 144 = 0
    16'b00111000_10010001 : OUT <= 0;  //56 / 145 = 0
    16'b00111000_10010010 : OUT <= 0;  //56 / 146 = 0
    16'b00111000_10010011 : OUT <= 0;  //56 / 147 = 0
    16'b00111000_10010100 : OUT <= 0;  //56 / 148 = 0
    16'b00111000_10010101 : OUT <= 0;  //56 / 149 = 0
    16'b00111000_10010110 : OUT <= 0;  //56 / 150 = 0
    16'b00111000_10010111 : OUT <= 0;  //56 / 151 = 0
    16'b00111000_10011000 : OUT <= 0;  //56 / 152 = 0
    16'b00111000_10011001 : OUT <= 0;  //56 / 153 = 0
    16'b00111000_10011010 : OUT <= 0;  //56 / 154 = 0
    16'b00111000_10011011 : OUT <= 0;  //56 / 155 = 0
    16'b00111000_10011100 : OUT <= 0;  //56 / 156 = 0
    16'b00111000_10011101 : OUT <= 0;  //56 / 157 = 0
    16'b00111000_10011110 : OUT <= 0;  //56 / 158 = 0
    16'b00111000_10011111 : OUT <= 0;  //56 / 159 = 0
    16'b00111000_10100000 : OUT <= 0;  //56 / 160 = 0
    16'b00111000_10100001 : OUT <= 0;  //56 / 161 = 0
    16'b00111000_10100010 : OUT <= 0;  //56 / 162 = 0
    16'b00111000_10100011 : OUT <= 0;  //56 / 163 = 0
    16'b00111000_10100100 : OUT <= 0;  //56 / 164 = 0
    16'b00111000_10100101 : OUT <= 0;  //56 / 165 = 0
    16'b00111000_10100110 : OUT <= 0;  //56 / 166 = 0
    16'b00111000_10100111 : OUT <= 0;  //56 / 167 = 0
    16'b00111000_10101000 : OUT <= 0;  //56 / 168 = 0
    16'b00111000_10101001 : OUT <= 0;  //56 / 169 = 0
    16'b00111000_10101010 : OUT <= 0;  //56 / 170 = 0
    16'b00111000_10101011 : OUT <= 0;  //56 / 171 = 0
    16'b00111000_10101100 : OUT <= 0;  //56 / 172 = 0
    16'b00111000_10101101 : OUT <= 0;  //56 / 173 = 0
    16'b00111000_10101110 : OUT <= 0;  //56 / 174 = 0
    16'b00111000_10101111 : OUT <= 0;  //56 / 175 = 0
    16'b00111000_10110000 : OUT <= 0;  //56 / 176 = 0
    16'b00111000_10110001 : OUT <= 0;  //56 / 177 = 0
    16'b00111000_10110010 : OUT <= 0;  //56 / 178 = 0
    16'b00111000_10110011 : OUT <= 0;  //56 / 179 = 0
    16'b00111000_10110100 : OUT <= 0;  //56 / 180 = 0
    16'b00111000_10110101 : OUT <= 0;  //56 / 181 = 0
    16'b00111000_10110110 : OUT <= 0;  //56 / 182 = 0
    16'b00111000_10110111 : OUT <= 0;  //56 / 183 = 0
    16'b00111000_10111000 : OUT <= 0;  //56 / 184 = 0
    16'b00111000_10111001 : OUT <= 0;  //56 / 185 = 0
    16'b00111000_10111010 : OUT <= 0;  //56 / 186 = 0
    16'b00111000_10111011 : OUT <= 0;  //56 / 187 = 0
    16'b00111000_10111100 : OUT <= 0;  //56 / 188 = 0
    16'b00111000_10111101 : OUT <= 0;  //56 / 189 = 0
    16'b00111000_10111110 : OUT <= 0;  //56 / 190 = 0
    16'b00111000_10111111 : OUT <= 0;  //56 / 191 = 0
    16'b00111000_11000000 : OUT <= 0;  //56 / 192 = 0
    16'b00111000_11000001 : OUT <= 0;  //56 / 193 = 0
    16'b00111000_11000010 : OUT <= 0;  //56 / 194 = 0
    16'b00111000_11000011 : OUT <= 0;  //56 / 195 = 0
    16'b00111000_11000100 : OUT <= 0;  //56 / 196 = 0
    16'b00111000_11000101 : OUT <= 0;  //56 / 197 = 0
    16'b00111000_11000110 : OUT <= 0;  //56 / 198 = 0
    16'b00111000_11000111 : OUT <= 0;  //56 / 199 = 0
    16'b00111000_11001000 : OUT <= 0;  //56 / 200 = 0
    16'b00111000_11001001 : OUT <= 0;  //56 / 201 = 0
    16'b00111000_11001010 : OUT <= 0;  //56 / 202 = 0
    16'b00111000_11001011 : OUT <= 0;  //56 / 203 = 0
    16'b00111000_11001100 : OUT <= 0;  //56 / 204 = 0
    16'b00111000_11001101 : OUT <= 0;  //56 / 205 = 0
    16'b00111000_11001110 : OUT <= 0;  //56 / 206 = 0
    16'b00111000_11001111 : OUT <= 0;  //56 / 207 = 0
    16'b00111000_11010000 : OUT <= 0;  //56 / 208 = 0
    16'b00111000_11010001 : OUT <= 0;  //56 / 209 = 0
    16'b00111000_11010010 : OUT <= 0;  //56 / 210 = 0
    16'b00111000_11010011 : OUT <= 0;  //56 / 211 = 0
    16'b00111000_11010100 : OUT <= 0;  //56 / 212 = 0
    16'b00111000_11010101 : OUT <= 0;  //56 / 213 = 0
    16'b00111000_11010110 : OUT <= 0;  //56 / 214 = 0
    16'b00111000_11010111 : OUT <= 0;  //56 / 215 = 0
    16'b00111000_11011000 : OUT <= 0;  //56 / 216 = 0
    16'b00111000_11011001 : OUT <= 0;  //56 / 217 = 0
    16'b00111000_11011010 : OUT <= 0;  //56 / 218 = 0
    16'b00111000_11011011 : OUT <= 0;  //56 / 219 = 0
    16'b00111000_11011100 : OUT <= 0;  //56 / 220 = 0
    16'b00111000_11011101 : OUT <= 0;  //56 / 221 = 0
    16'b00111000_11011110 : OUT <= 0;  //56 / 222 = 0
    16'b00111000_11011111 : OUT <= 0;  //56 / 223 = 0
    16'b00111000_11100000 : OUT <= 0;  //56 / 224 = 0
    16'b00111000_11100001 : OUT <= 0;  //56 / 225 = 0
    16'b00111000_11100010 : OUT <= 0;  //56 / 226 = 0
    16'b00111000_11100011 : OUT <= 0;  //56 / 227 = 0
    16'b00111000_11100100 : OUT <= 0;  //56 / 228 = 0
    16'b00111000_11100101 : OUT <= 0;  //56 / 229 = 0
    16'b00111000_11100110 : OUT <= 0;  //56 / 230 = 0
    16'b00111000_11100111 : OUT <= 0;  //56 / 231 = 0
    16'b00111000_11101000 : OUT <= 0;  //56 / 232 = 0
    16'b00111000_11101001 : OUT <= 0;  //56 / 233 = 0
    16'b00111000_11101010 : OUT <= 0;  //56 / 234 = 0
    16'b00111000_11101011 : OUT <= 0;  //56 / 235 = 0
    16'b00111000_11101100 : OUT <= 0;  //56 / 236 = 0
    16'b00111000_11101101 : OUT <= 0;  //56 / 237 = 0
    16'b00111000_11101110 : OUT <= 0;  //56 / 238 = 0
    16'b00111000_11101111 : OUT <= 0;  //56 / 239 = 0
    16'b00111000_11110000 : OUT <= 0;  //56 / 240 = 0
    16'b00111000_11110001 : OUT <= 0;  //56 / 241 = 0
    16'b00111000_11110010 : OUT <= 0;  //56 / 242 = 0
    16'b00111000_11110011 : OUT <= 0;  //56 / 243 = 0
    16'b00111000_11110100 : OUT <= 0;  //56 / 244 = 0
    16'b00111000_11110101 : OUT <= 0;  //56 / 245 = 0
    16'b00111000_11110110 : OUT <= 0;  //56 / 246 = 0
    16'b00111000_11110111 : OUT <= 0;  //56 / 247 = 0
    16'b00111000_11111000 : OUT <= 0;  //56 / 248 = 0
    16'b00111000_11111001 : OUT <= 0;  //56 / 249 = 0
    16'b00111000_11111010 : OUT <= 0;  //56 / 250 = 0
    16'b00111000_11111011 : OUT <= 0;  //56 / 251 = 0
    16'b00111000_11111100 : OUT <= 0;  //56 / 252 = 0
    16'b00111000_11111101 : OUT <= 0;  //56 / 253 = 0
    16'b00111000_11111110 : OUT <= 0;  //56 / 254 = 0
    16'b00111000_11111111 : OUT <= 0;  //56 / 255 = 0
    16'b00111001_00000000 : OUT <= 0;  //57 / 0 = 0
    16'b00111001_00000001 : OUT <= 57;  //57 / 1 = 57
    16'b00111001_00000010 : OUT <= 28;  //57 / 2 = 28
    16'b00111001_00000011 : OUT <= 19;  //57 / 3 = 19
    16'b00111001_00000100 : OUT <= 14;  //57 / 4 = 14
    16'b00111001_00000101 : OUT <= 11;  //57 / 5 = 11
    16'b00111001_00000110 : OUT <= 9;  //57 / 6 = 9
    16'b00111001_00000111 : OUT <= 8;  //57 / 7 = 8
    16'b00111001_00001000 : OUT <= 7;  //57 / 8 = 7
    16'b00111001_00001001 : OUT <= 6;  //57 / 9 = 6
    16'b00111001_00001010 : OUT <= 5;  //57 / 10 = 5
    16'b00111001_00001011 : OUT <= 5;  //57 / 11 = 5
    16'b00111001_00001100 : OUT <= 4;  //57 / 12 = 4
    16'b00111001_00001101 : OUT <= 4;  //57 / 13 = 4
    16'b00111001_00001110 : OUT <= 4;  //57 / 14 = 4
    16'b00111001_00001111 : OUT <= 3;  //57 / 15 = 3
    16'b00111001_00010000 : OUT <= 3;  //57 / 16 = 3
    16'b00111001_00010001 : OUT <= 3;  //57 / 17 = 3
    16'b00111001_00010010 : OUT <= 3;  //57 / 18 = 3
    16'b00111001_00010011 : OUT <= 3;  //57 / 19 = 3
    16'b00111001_00010100 : OUT <= 2;  //57 / 20 = 2
    16'b00111001_00010101 : OUT <= 2;  //57 / 21 = 2
    16'b00111001_00010110 : OUT <= 2;  //57 / 22 = 2
    16'b00111001_00010111 : OUT <= 2;  //57 / 23 = 2
    16'b00111001_00011000 : OUT <= 2;  //57 / 24 = 2
    16'b00111001_00011001 : OUT <= 2;  //57 / 25 = 2
    16'b00111001_00011010 : OUT <= 2;  //57 / 26 = 2
    16'b00111001_00011011 : OUT <= 2;  //57 / 27 = 2
    16'b00111001_00011100 : OUT <= 2;  //57 / 28 = 2
    16'b00111001_00011101 : OUT <= 1;  //57 / 29 = 1
    16'b00111001_00011110 : OUT <= 1;  //57 / 30 = 1
    16'b00111001_00011111 : OUT <= 1;  //57 / 31 = 1
    16'b00111001_00100000 : OUT <= 1;  //57 / 32 = 1
    16'b00111001_00100001 : OUT <= 1;  //57 / 33 = 1
    16'b00111001_00100010 : OUT <= 1;  //57 / 34 = 1
    16'b00111001_00100011 : OUT <= 1;  //57 / 35 = 1
    16'b00111001_00100100 : OUT <= 1;  //57 / 36 = 1
    16'b00111001_00100101 : OUT <= 1;  //57 / 37 = 1
    16'b00111001_00100110 : OUT <= 1;  //57 / 38 = 1
    16'b00111001_00100111 : OUT <= 1;  //57 / 39 = 1
    16'b00111001_00101000 : OUT <= 1;  //57 / 40 = 1
    16'b00111001_00101001 : OUT <= 1;  //57 / 41 = 1
    16'b00111001_00101010 : OUT <= 1;  //57 / 42 = 1
    16'b00111001_00101011 : OUT <= 1;  //57 / 43 = 1
    16'b00111001_00101100 : OUT <= 1;  //57 / 44 = 1
    16'b00111001_00101101 : OUT <= 1;  //57 / 45 = 1
    16'b00111001_00101110 : OUT <= 1;  //57 / 46 = 1
    16'b00111001_00101111 : OUT <= 1;  //57 / 47 = 1
    16'b00111001_00110000 : OUT <= 1;  //57 / 48 = 1
    16'b00111001_00110001 : OUT <= 1;  //57 / 49 = 1
    16'b00111001_00110010 : OUT <= 1;  //57 / 50 = 1
    16'b00111001_00110011 : OUT <= 1;  //57 / 51 = 1
    16'b00111001_00110100 : OUT <= 1;  //57 / 52 = 1
    16'b00111001_00110101 : OUT <= 1;  //57 / 53 = 1
    16'b00111001_00110110 : OUT <= 1;  //57 / 54 = 1
    16'b00111001_00110111 : OUT <= 1;  //57 / 55 = 1
    16'b00111001_00111000 : OUT <= 1;  //57 / 56 = 1
    16'b00111001_00111001 : OUT <= 1;  //57 / 57 = 1
    16'b00111001_00111010 : OUT <= 0;  //57 / 58 = 0
    16'b00111001_00111011 : OUT <= 0;  //57 / 59 = 0
    16'b00111001_00111100 : OUT <= 0;  //57 / 60 = 0
    16'b00111001_00111101 : OUT <= 0;  //57 / 61 = 0
    16'b00111001_00111110 : OUT <= 0;  //57 / 62 = 0
    16'b00111001_00111111 : OUT <= 0;  //57 / 63 = 0
    16'b00111001_01000000 : OUT <= 0;  //57 / 64 = 0
    16'b00111001_01000001 : OUT <= 0;  //57 / 65 = 0
    16'b00111001_01000010 : OUT <= 0;  //57 / 66 = 0
    16'b00111001_01000011 : OUT <= 0;  //57 / 67 = 0
    16'b00111001_01000100 : OUT <= 0;  //57 / 68 = 0
    16'b00111001_01000101 : OUT <= 0;  //57 / 69 = 0
    16'b00111001_01000110 : OUT <= 0;  //57 / 70 = 0
    16'b00111001_01000111 : OUT <= 0;  //57 / 71 = 0
    16'b00111001_01001000 : OUT <= 0;  //57 / 72 = 0
    16'b00111001_01001001 : OUT <= 0;  //57 / 73 = 0
    16'b00111001_01001010 : OUT <= 0;  //57 / 74 = 0
    16'b00111001_01001011 : OUT <= 0;  //57 / 75 = 0
    16'b00111001_01001100 : OUT <= 0;  //57 / 76 = 0
    16'b00111001_01001101 : OUT <= 0;  //57 / 77 = 0
    16'b00111001_01001110 : OUT <= 0;  //57 / 78 = 0
    16'b00111001_01001111 : OUT <= 0;  //57 / 79 = 0
    16'b00111001_01010000 : OUT <= 0;  //57 / 80 = 0
    16'b00111001_01010001 : OUT <= 0;  //57 / 81 = 0
    16'b00111001_01010010 : OUT <= 0;  //57 / 82 = 0
    16'b00111001_01010011 : OUT <= 0;  //57 / 83 = 0
    16'b00111001_01010100 : OUT <= 0;  //57 / 84 = 0
    16'b00111001_01010101 : OUT <= 0;  //57 / 85 = 0
    16'b00111001_01010110 : OUT <= 0;  //57 / 86 = 0
    16'b00111001_01010111 : OUT <= 0;  //57 / 87 = 0
    16'b00111001_01011000 : OUT <= 0;  //57 / 88 = 0
    16'b00111001_01011001 : OUT <= 0;  //57 / 89 = 0
    16'b00111001_01011010 : OUT <= 0;  //57 / 90 = 0
    16'b00111001_01011011 : OUT <= 0;  //57 / 91 = 0
    16'b00111001_01011100 : OUT <= 0;  //57 / 92 = 0
    16'b00111001_01011101 : OUT <= 0;  //57 / 93 = 0
    16'b00111001_01011110 : OUT <= 0;  //57 / 94 = 0
    16'b00111001_01011111 : OUT <= 0;  //57 / 95 = 0
    16'b00111001_01100000 : OUT <= 0;  //57 / 96 = 0
    16'b00111001_01100001 : OUT <= 0;  //57 / 97 = 0
    16'b00111001_01100010 : OUT <= 0;  //57 / 98 = 0
    16'b00111001_01100011 : OUT <= 0;  //57 / 99 = 0
    16'b00111001_01100100 : OUT <= 0;  //57 / 100 = 0
    16'b00111001_01100101 : OUT <= 0;  //57 / 101 = 0
    16'b00111001_01100110 : OUT <= 0;  //57 / 102 = 0
    16'b00111001_01100111 : OUT <= 0;  //57 / 103 = 0
    16'b00111001_01101000 : OUT <= 0;  //57 / 104 = 0
    16'b00111001_01101001 : OUT <= 0;  //57 / 105 = 0
    16'b00111001_01101010 : OUT <= 0;  //57 / 106 = 0
    16'b00111001_01101011 : OUT <= 0;  //57 / 107 = 0
    16'b00111001_01101100 : OUT <= 0;  //57 / 108 = 0
    16'b00111001_01101101 : OUT <= 0;  //57 / 109 = 0
    16'b00111001_01101110 : OUT <= 0;  //57 / 110 = 0
    16'b00111001_01101111 : OUT <= 0;  //57 / 111 = 0
    16'b00111001_01110000 : OUT <= 0;  //57 / 112 = 0
    16'b00111001_01110001 : OUT <= 0;  //57 / 113 = 0
    16'b00111001_01110010 : OUT <= 0;  //57 / 114 = 0
    16'b00111001_01110011 : OUT <= 0;  //57 / 115 = 0
    16'b00111001_01110100 : OUT <= 0;  //57 / 116 = 0
    16'b00111001_01110101 : OUT <= 0;  //57 / 117 = 0
    16'b00111001_01110110 : OUT <= 0;  //57 / 118 = 0
    16'b00111001_01110111 : OUT <= 0;  //57 / 119 = 0
    16'b00111001_01111000 : OUT <= 0;  //57 / 120 = 0
    16'b00111001_01111001 : OUT <= 0;  //57 / 121 = 0
    16'b00111001_01111010 : OUT <= 0;  //57 / 122 = 0
    16'b00111001_01111011 : OUT <= 0;  //57 / 123 = 0
    16'b00111001_01111100 : OUT <= 0;  //57 / 124 = 0
    16'b00111001_01111101 : OUT <= 0;  //57 / 125 = 0
    16'b00111001_01111110 : OUT <= 0;  //57 / 126 = 0
    16'b00111001_01111111 : OUT <= 0;  //57 / 127 = 0
    16'b00111001_10000000 : OUT <= 0;  //57 / 128 = 0
    16'b00111001_10000001 : OUT <= 0;  //57 / 129 = 0
    16'b00111001_10000010 : OUT <= 0;  //57 / 130 = 0
    16'b00111001_10000011 : OUT <= 0;  //57 / 131 = 0
    16'b00111001_10000100 : OUT <= 0;  //57 / 132 = 0
    16'b00111001_10000101 : OUT <= 0;  //57 / 133 = 0
    16'b00111001_10000110 : OUT <= 0;  //57 / 134 = 0
    16'b00111001_10000111 : OUT <= 0;  //57 / 135 = 0
    16'b00111001_10001000 : OUT <= 0;  //57 / 136 = 0
    16'b00111001_10001001 : OUT <= 0;  //57 / 137 = 0
    16'b00111001_10001010 : OUT <= 0;  //57 / 138 = 0
    16'b00111001_10001011 : OUT <= 0;  //57 / 139 = 0
    16'b00111001_10001100 : OUT <= 0;  //57 / 140 = 0
    16'b00111001_10001101 : OUT <= 0;  //57 / 141 = 0
    16'b00111001_10001110 : OUT <= 0;  //57 / 142 = 0
    16'b00111001_10001111 : OUT <= 0;  //57 / 143 = 0
    16'b00111001_10010000 : OUT <= 0;  //57 / 144 = 0
    16'b00111001_10010001 : OUT <= 0;  //57 / 145 = 0
    16'b00111001_10010010 : OUT <= 0;  //57 / 146 = 0
    16'b00111001_10010011 : OUT <= 0;  //57 / 147 = 0
    16'b00111001_10010100 : OUT <= 0;  //57 / 148 = 0
    16'b00111001_10010101 : OUT <= 0;  //57 / 149 = 0
    16'b00111001_10010110 : OUT <= 0;  //57 / 150 = 0
    16'b00111001_10010111 : OUT <= 0;  //57 / 151 = 0
    16'b00111001_10011000 : OUT <= 0;  //57 / 152 = 0
    16'b00111001_10011001 : OUT <= 0;  //57 / 153 = 0
    16'b00111001_10011010 : OUT <= 0;  //57 / 154 = 0
    16'b00111001_10011011 : OUT <= 0;  //57 / 155 = 0
    16'b00111001_10011100 : OUT <= 0;  //57 / 156 = 0
    16'b00111001_10011101 : OUT <= 0;  //57 / 157 = 0
    16'b00111001_10011110 : OUT <= 0;  //57 / 158 = 0
    16'b00111001_10011111 : OUT <= 0;  //57 / 159 = 0
    16'b00111001_10100000 : OUT <= 0;  //57 / 160 = 0
    16'b00111001_10100001 : OUT <= 0;  //57 / 161 = 0
    16'b00111001_10100010 : OUT <= 0;  //57 / 162 = 0
    16'b00111001_10100011 : OUT <= 0;  //57 / 163 = 0
    16'b00111001_10100100 : OUT <= 0;  //57 / 164 = 0
    16'b00111001_10100101 : OUT <= 0;  //57 / 165 = 0
    16'b00111001_10100110 : OUT <= 0;  //57 / 166 = 0
    16'b00111001_10100111 : OUT <= 0;  //57 / 167 = 0
    16'b00111001_10101000 : OUT <= 0;  //57 / 168 = 0
    16'b00111001_10101001 : OUT <= 0;  //57 / 169 = 0
    16'b00111001_10101010 : OUT <= 0;  //57 / 170 = 0
    16'b00111001_10101011 : OUT <= 0;  //57 / 171 = 0
    16'b00111001_10101100 : OUT <= 0;  //57 / 172 = 0
    16'b00111001_10101101 : OUT <= 0;  //57 / 173 = 0
    16'b00111001_10101110 : OUT <= 0;  //57 / 174 = 0
    16'b00111001_10101111 : OUT <= 0;  //57 / 175 = 0
    16'b00111001_10110000 : OUT <= 0;  //57 / 176 = 0
    16'b00111001_10110001 : OUT <= 0;  //57 / 177 = 0
    16'b00111001_10110010 : OUT <= 0;  //57 / 178 = 0
    16'b00111001_10110011 : OUT <= 0;  //57 / 179 = 0
    16'b00111001_10110100 : OUT <= 0;  //57 / 180 = 0
    16'b00111001_10110101 : OUT <= 0;  //57 / 181 = 0
    16'b00111001_10110110 : OUT <= 0;  //57 / 182 = 0
    16'b00111001_10110111 : OUT <= 0;  //57 / 183 = 0
    16'b00111001_10111000 : OUT <= 0;  //57 / 184 = 0
    16'b00111001_10111001 : OUT <= 0;  //57 / 185 = 0
    16'b00111001_10111010 : OUT <= 0;  //57 / 186 = 0
    16'b00111001_10111011 : OUT <= 0;  //57 / 187 = 0
    16'b00111001_10111100 : OUT <= 0;  //57 / 188 = 0
    16'b00111001_10111101 : OUT <= 0;  //57 / 189 = 0
    16'b00111001_10111110 : OUT <= 0;  //57 / 190 = 0
    16'b00111001_10111111 : OUT <= 0;  //57 / 191 = 0
    16'b00111001_11000000 : OUT <= 0;  //57 / 192 = 0
    16'b00111001_11000001 : OUT <= 0;  //57 / 193 = 0
    16'b00111001_11000010 : OUT <= 0;  //57 / 194 = 0
    16'b00111001_11000011 : OUT <= 0;  //57 / 195 = 0
    16'b00111001_11000100 : OUT <= 0;  //57 / 196 = 0
    16'b00111001_11000101 : OUT <= 0;  //57 / 197 = 0
    16'b00111001_11000110 : OUT <= 0;  //57 / 198 = 0
    16'b00111001_11000111 : OUT <= 0;  //57 / 199 = 0
    16'b00111001_11001000 : OUT <= 0;  //57 / 200 = 0
    16'b00111001_11001001 : OUT <= 0;  //57 / 201 = 0
    16'b00111001_11001010 : OUT <= 0;  //57 / 202 = 0
    16'b00111001_11001011 : OUT <= 0;  //57 / 203 = 0
    16'b00111001_11001100 : OUT <= 0;  //57 / 204 = 0
    16'b00111001_11001101 : OUT <= 0;  //57 / 205 = 0
    16'b00111001_11001110 : OUT <= 0;  //57 / 206 = 0
    16'b00111001_11001111 : OUT <= 0;  //57 / 207 = 0
    16'b00111001_11010000 : OUT <= 0;  //57 / 208 = 0
    16'b00111001_11010001 : OUT <= 0;  //57 / 209 = 0
    16'b00111001_11010010 : OUT <= 0;  //57 / 210 = 0
    16'b00111001_11010011 : OUT <= 0;  //57 / 211 = 0
    16'b00111001_11010100 : OUT <= 0;  //57 / 212 = 0
    16'b00111001_11010101 : OUT <= 0;  //57 / 213 = 0
    16'b00111001_11010110 : OUT <= 0;  //57 / 214 = 0
    16'b00111001_11010111 : OUT <= 0;  //57 / 215 = 0
    16'b00111001_11011000 : OUT <= 0;  //57 / 216 = 0
    16'b00111001_11011001 : OUT <= 0;  //57 / 217 = 0
    16'b00111001_11011010 : OUT <= 0;  //57 / 218 = 0
    16'b00111001_11011011 : OUT <= 0;  //57 / 219 = 0
    16'b00111001_11011100 : OUT <= 0;  //57 / 220 = 0
    16'b00111001_11011101 : OUT <= 0;  //57 / 221 = 0
    16'b00111001_11011110 : OUT <= 0;  //57 / 222 = 0
    16'b00111001_11011111 : OUT <= 0;  //57 / 223 = 0
    16'b00111001_11100000 : OUT <= 0;  //57 / 224 = 0
    16'b00111001_11100001 : OUT <= 0;  //57 / 225 = 0
    16'b00111001_11100010 : OUT <= 0;  //57 / 226 = 0
    16'b00111001_11100011 : OUT <= 0;  //57 / 227 = 0
    16'b00111001_11100100 : OUT <= 0;  //57 / 228 = 0
    16'b00111001_11100101 : OUT <= 0;  //57 / 229 = 0
    16'b00111001_11100110 : OUT <= 0;  //57 / 230 = 0
    16'b00111001_11100111 : OUT <= 0;  //57 / 231 = 0
    16'b00111001_11101000 : OUT <= 0;  //57 / 232 = 0
    16'b00111001_11101001 : OUT <= 0;  //57 / 233 = 0
    16'b00111001_11101010 : OUT <= 0;  //57 / 234 = 0
    16'b00111001_11101011 : OUT <= 0;  //57 / 235 = 0
    16'b00111001_11101100 : OUT <= 0;  //57 / 236 = 0
    16'b00111001_11101101 : OUT <= 0;  //57 / 237 = 0
    16'b00111001_11101110 : OUT <= 0;  //57 / 238 = 0
    16'b00111001_11101111 : OUT <= 0;  //57 / 239 = 0
    16'b00111001_11110000 : OUT <= 0;  //57 / 240 = 0
    16'b00111001_11110001 : OUT <= 0;  //57 / 241 = 0
    16'b00111001_11110010 : OUT <= 0;  //57 / 242 = 0
    16'b00111001_11110011 : OUT <= 0;  //57 / 243 = 0
    16'b00111001_11110100 : OUT <= 0;  //57 / 244 = 0
    16'b00111001_11110101 : OUT <= 0;  //57 / 245 = 0
    16'b00111001_11110110 : OUT <= 0;  //57 / 246 = 0
    16'b00111001_11110111 : OUT <= 0;  //57 / 247 = 0
    16'b00111001_11111000 : OUT <= 0;  //57 / 248 = 0
    16'b00111001_11111001 : OUT <= 0;  //57 / 249 = 0
    16'b00111001_11111010 : OUT <= 0;  //57 / 250 = 0
    16'b00111001_11111011 : OUT <= 0;  //57 / 251 = 0
    16'b00111001_11111100 : OUT <= 0;  //57 / 252 = 0
    16'b00111001_11111101 : OUT <= 0;  //57 / 253 = 0
    16'b00111001_11111110 : OUT <= 0;  //57 / 254 = 0
    16'b00111001_11111111 : OUT <= 0;  //57 / 255 = 0
    16'b00111010_00000000 : OUT <= 0;  //58 / 0 = 0
    16'b00111010_00000001 : OUT <= 58;  //58 / 1 = 58
    16'b00111010_00000010 : OUT <= 29;  //58 / 2 = 29
    16'b00111010_00000011 : OUT <= 19;  //58 / 3 = 19
    16'b00111010_00000100 : OUT <= 14;  //58 / 4 = 14
    16'b00111010_00000101 : OUT <= 11;  //58 / 5 = 11
    16'b00111010_00000110 : OUT <= 9;  //58 / 6 = 9
    16'b00111010_00000111 : OUT <= 8;  //58 / 7 = 8
    16'b00111010_00001000 : OUT <= 7;  //58 / 8 = 7
    16'b00111010_00001001 : OUT <= 6;  //58 / 9 = 6
    16'b00111010_00001010 : OUT <= 5;  //58 / 10 = 5
    16'b00111010_00001011 : OUT <= 5;  //58 / 11 = 5
    16'b00111010_00001100 : OUT <= 4;  //58 / 12 = 4
    16'b00111010_00001101 : OUT <= 4;  //58 / 13 = 4
    16'b00111010_00001110 : OUT <= 4;  //58 / 14 = 4
    16'b00111010_00001111 : OUT <= 3;  //58 / 15 = 3
    16'b00111010_00010000 : OUT <= 3;  //58 / 16 = 3
    16'b00111010_00010001 : OUT <= 3;  //58 / 17 = 3
    16'b00111010_00010010 : OUT <= 3;  //58 / 18 = 3
    16'b00111010_00010011 : OUT <= 3;  //58 / 19 = 3
    16'b00111010_00010100 : OUT <= 2;  //58 / 20 = 2
    16'b00111010_00010101 : OUT <= 2;  //58 / 21 = 2
    16'b00111010_00010110 : OUT <= 2;  //58 / 22 = 2
    16'b00111010_00010111 : OUT <= 2;  //58 / 23 = 2
    16'b00111010_00011000 : OUT <= 2;  //58 / 24 = 2
    16'b00111010_00011001 : OUT <= 2;  //58 / 25 = 2
    16'b00111010_00011010 : OUT <= 2;  //58 / 26 = 2
    16'b00111010_00011011 : OUT <= 2;  //58 / 27 = 2
    16'b00111010_00011100 : OUT <= 2;  //58 / 28 = 2
    16'b00111010_00011101 : OUT <= 2;  //58 / 29 = 2
    16'b00111010_00011110 : OUT <= 1;  //58 / 30 = 1
    16'b00111010_00011111 : OUT <= 1;  //58 / 31 = 1
    16'b00111010_00100000 : OUT <= 1;  //58 / 32 = 1
    16'b00111010_00100001 : OUT <= 1;  //58 / 33 = 1
    16'b00111010_00100010 : OUT <= 1;  //58 / 34 = 1
    16'b00111010_00100011 : OUT <= 1;  //58 / 35 = 1
    16'b00111010_00100100 : OUT <= 1;  //58 / 36 = 1
    16'b00111010_00100101 : OUT <= 1;  //58 / 37 = 1
    16'b00111010_00100110 : OUT <= 1;  //58 / 38 = 1
    16'b00111010_00100111 : OUT <= 1;  //58 / 39 = 1
    16'b00111010_00101000 : OUT <= 1;  //58 / 40 = 1
    16'b00111010_00101001 : OUT <= 1;  //58 / 41 = 1
    16'b00111010_00101010 : OUT <= 1;  //58 / 42 = 1
    16'b00111010_00101011 : OUT <= 1;  //58 / 43 = 1
    16'b00111010_00101100 : OUT <= 1;  //58 / 44 = 1
    16'b00111010_00101101 : OUT <= 1;  //58 / 45 = 1
    16'b00111010_00101110 : OUT <= 1;  //58 / 46 = 1
    16'b00111010_00101111 : OUT <= 1;  //58 / 47 = 1
    16'b00111010_00110000 : OUT <= 1;  //58 / 48 = 1
    16'b00111010_00110001 : OUT <= 1;  //58 / 49 = 1
    16'b00111010_00110010 : OUT <= 1;  //58 / 50 = 1
    16'b00111010_00110011 : OUT <= 1;  //58 / 51 = 1
    16'b00111010_00110100 : OUT <= 1;  //58 / 52 = 1
    16'b00111010_00110101 : OUT <= 1;  //58 / 53 = 1
    16'b00111010_00110110 : OUT <= 1;  //58 / 54 = 1
    16'b00111010_00110111 : OUT <= 1;  //58 / 55 = 1
    16'b00111010_00111000 : OUT <= 1;  //58 / 56 = 1
    16'b00111010_00111001 : OUT <= 1;  //58 / 57 = 1
    16'b00111010_00111010 : OUT <= 1;  //58 / 58 = 1
    16'b00111010_00111011 : OUT <= 0;  //58 / 59 = 0
    16'b00111010_00111100 : OUT <= 0;  //58 / 60 = 0
    16'b00111010_00111101 : OUT <= 0;  //58 / 61 = 0
    16'b00111010_00111110 : OUT <= 0;  //58 / 62 = 0
    16'b00111010_00111111 : OUT <= 0;  //58 / 63 = 0
    16'b00111010_01000000 : OUT <= 0;  //58 / 64 = 0
    16'b00111010_01000001 : OUT <= 0;  //58 / 65 = 0
    16'b00111010_01000010 : OUT <= 0;  //58 / 66 = 0
    16'b00111010_01000011 : OUT <= 0;  //58 / 67 = 0
    16'b00111010_01000100 : OUT <= 0;  //58 / 68 = 0
    16'b00111010_01000101 : OUT <= 0;  //58 / 69 = 0
    16'b00111010_01000110 : OUT <= 0;  //58 / 70 = 0
    16'b00111010_01000111 : OUT <= 0;  //58 / 71 = 0
    16'b00111010_01001000 : OUT <= 0;  //58 / 72 = 0
    16'b00111010_01001001 : OUT <= 0;  //58 / 73 = 0
    16'b00111010_01001010 : OUT <= 0;  //58 / 74 = 0
    16'b00111010_01001011 : OUT <= 0;  //58 / 75 = 0
    16'b00111010_01001100 : OUT <= 0;  //58 / 76 = 0
    16'b00111010_01001101 : OUT <= 0;  //58 / 77 = 0
    16'b00111010_01001110 : OUT <= 0;  //58 / 78 = 0
    16'b00111010_01001111 : OUT <= 0;  //58 / 79 = 0
    16'b00111010_01010000 : OUT <= 0;  //58 / 80 = 0
    16'b00111010_01010001 : OUT <= 0;  //58 / 81 = 0
    16'b00111010_01010010 : OUT <= 0;  //58 / 82 = 0
    16'b00111010_01010011 : OUT <= 0;  //58 / 83 = 0
    16'b00111010_01010100 : OUT <= 0;  //58 / 84 = 0
    16'b00111010_01010101 : OUT <= 0;  //58 / 85 = 0
    16'b00111010_01010110 : OUT <= 0;  //58 / 86 = 0
    16'b00111010_01010111 : OUT <= 0;  //58 / 87 = 0
    16'b00111010_01011000 : OUT <= 0;  //58 / 88 = 0
    16'b00111010_01011001 : OUT <= 0;  //58 / 89 = 0
    16'b00111010_01011010 : OUT <= 0;  //58 / 90 = 0
    16'b00111010_01011011 : OUT <= 0;  //58 / 91 = 0
    16'b00111010_01011100 : OUT <= 0;  //58 / 92 = 0
    16'b00111010_01011101 : OUT <= 0;  //58 / 93 = 0
    16'b00111010_01011110 : OUT <= 0;  //58 / 94 = 0
    16'b00111010_01011111 : OUT <= 0;  //58 / 95 = 0
    16'b00111010_01100000 : OUT <= 0;  //58 / 96 = 0
    16'b00111010_01100001 : OUT <= 0;  //58 / 97 = 0
    16'b00111010_01100010 : OUT <= 0;  //58 / 98 = 0
    16'b00111010_01100011 : OUT <= 0;  //58 / 99 = 0
    16'b00111010_01100100 : OUT <= 0;  //58 / 100 = 0
    16'b00111010_01100101 : OUT <= 0;  //58 / 101 = 0
    16'b00111010_01100110 : OUT <= 0;  //58 / 102 = 0
    16'b00111010_01100111 : OUT <= 0;  //58 / 103 = 0
    16'b00111010_01101000 : OUT <= 0;  //58 / 104 = 0
    16'b00111010_01101001 : OUT <= 0;  //58 / 105 = 0
    16'b00111010_01101010 : OUT <= 0;  //58 / 106 = 0
    16'b00111010_01101011 : OUT <= 0;  //58 / 107 = 0
    16'b00111010_01101100 : OUT <= 0;  //58 / 108 = 0
    16'b00111010_01101101 : OUT <= 0;  //58 / 109 = 0
    16'b00111010_01101110 : OUT <= 0;  //58 / 110 = 0
    16'b00111010_01101111 : OUT <= 0;  //58 / 111 = 0
    16'b00111010_01110000 : OUT <= 0;  //58 / 112 = 0
    16'b00111010_01110001 : OUT <= 0;  //58 / 113 = 0
    16'b00111010_01110010 : OUT <= 0;  //58 / 114 = 0
    16'b00111010_01110011 : OUT <= 0;  //58 / 115 = 0
    16'b00111010_01110100 : OUT <= 0;  //58 / 116 = 0
    16'b00111010_01110101 : OUT <= 0;  //58 / 117 = 0
    16'b00111010_01110110 : OUT <= 0;  //58 / 118 = 0
    16'b00111010_01110111 : OUT <= 0;  //58 / 119 = 0
    16'b00111010_01111000 : OUT <= 0;  //58 / 120 = 0
    16'b00111010_01111001 : OUT <= 0;  //58 / 121 = 0
    16'b00111010_01111010 : OUT <= 0;  //58 / 122 = 0
    16'b00111010_01111011 : OUT <= 0;  //58 / 123 = 0
    16'b00111010_01111100 : OUT <= 0;  //58 / 124 = 0
    16'b00111010_01111101 : OUT <= 0;  //58 / 125 = 0
    16'b00111010_01111110 : OUT <= 0;  //58 / 126 = 0
    16'b00111010_01111111 : OUT <= 0;  //58 / 127 = 0
    16'b00111010_10000000 : OUT <= 0;  //58 / 128 = 0
    16'b00111010_10000001 : OUT <= 0;  //58 / 129 = 0
    16'b00111010_10000010 : OUT <= 0;  //58 / 130 = 0
    16'b00111010_10000011 : OUT <= 0;  //58 / 131 = 0
    16'b00111010_10000100 : OUT <= 0;  //58 / 132 = 0
    16'b00111010_10000101 : OUT <= 0;  //58 / 133 = 0
    16'b00111010_10000110 : OUT <= 0;  //58 / 134 = 0
    16'b00111010_10000111 : OUT <= 0;  //58 / 135 = 0
    16'b00111010_10001000 : OUT <= 0;  //58 / 136 = 0
    16'b00111010_10001001 : OUT <= 0;  //58 / 137 = 0
    16'b00111010_10001010 : OUT <= 0;  //58 / 138 = 0
    16'b00111010_10001011 : OUT <= 0;  //58 / 139 = 0
    16'b00111010_10001100 : OUT <= 0;  //58 / 140 = 0
    16'b00111010_10001101 : OUT <= 0;  //58 / 141 = 0
    16'b00111010_10001110 : OUT <= 0;  //58 / 142 = 0
    16'b00111010_10001111 : OUT <= 0;  //58 / 143 = 0
    16'b00111010_10010000 : OUT <= 0;  //58 / 144 = 0
    16'b00111010_10010001 : OUT <= 0;  //58 / 145 = 0
    16'b00111010_10010010 : OUT <= 0;  //58 / 146 = 0
    16'b00111010_10010011 : OUT <= 0;  //58 / 147 = 0
    16'b00111010_10010100 : OUT <= 0;  //58 / 148 = 0
    16'b00111010_10010101 : OUT <= 0;  //58 / 149 = 0
    16'b00111010_10010110 : OUT <= 0;  //58 / 150 = 0
    16'b00111010_10010111 : OUT <= 0;  //58 / 151 = 0
    16'b00111010_10011000 : OUT <= 0;  //58 / 152 = 0
    16'b00111010_10011001 : OUT <= 0;  //58 / 153 = 0
    16'b00111010_10011010 : OUT <= 0;  //58 / 154 = 0
    16'b00111010_10011011 : OUT <= 0;  //58 / 155 = 0
    16'b00111010_10011100 : OUT <= 0;  //58 / 156 = 0
    16'b00111010_10011101 : OUT <= 0;  //58 / 157 = 0
    16'b00111010_10011110 : OUT <= 0;  //58 / 158 = 0
    16'b00111010_10011111 : OUT <= 0;  //58 / 159 = 0
    16'b00111010_10100000 : OUT <= 0;  //58 / 160 = 0
    16'b00111010_10100001 : OUT <= 0;  //58 / 161 = 0
    16'b00111010_10100010 : OUT <= 0;  //58 / 162 = 0
    16'b00111010_10100011 : OUT <= 0;  //58 / 163 = 0
    16'b00111010_10100100 : OUT <= 0;  //58 / 164 = 0
    16'b00111010_10100101 : OUT <= 0;  //58 / 165 = 0
    16'b00111010_10100110 : OUT <= 0;  //58 / 166 = 0
    16'b00111010_10100111 : OUT <= 0;  //58 / 167 = 0
    16'b00111010_10101000 : OUT <= 0;  //58 / 168 = 0
    16'b00111010_10101001 : OUT <= 0;  //58 / 169 = 0
    16'b00111010_10101010 : OUT <= 0;  //58 / 170 = 0
    16'b00111010_10101011 : OUT <= 0;  //58 / 171 = 0
    16'b00111010_10101100 : OUT <= 0;  //58 / 172 = 0
    16'b00111010_10101101 : OUT <= 0;  //58 / 173 = 0
    16'b00111010_10101110 : OUT <= 0;  //58 / 174 = 0
    16'b00111010_10101111 : OUT <= 0;  //58 / 175 = 0
    16'b00111010_10110000 : OUT <= 0;  //58 / 176 = 0
    16'b00111010_10110001 : OUT <= 0;  //58 / 177 = 0
    16'b00111010_10110010 : OUT <= 0;  //58 / 178 = 0
    16'b00111010_10110011 : OUT <= 0;  //58 / 179 = 0
    16'b00111010_10110100 : OUT <= 0;  //58 / 180 = 0
    16'b00111010_10110101 : OUT <= 0;  //58 / 181 = 0
    16'b00111010_10110110 : OUT <= 0;  //58 / 182 = 0
    16'b00111010_10110111 : OUT <= 0;  //58 / 183 = 0
    16'b00111010_10111000 : OUT <= 0;  //58 / 184 = 0
    16'b00111010_10111001 : OUT <= 0;  //58 / 185 = 0
    16'b00111010_10111010 : OUT <= 0;  //58 / 186 = 0
    16'b00111010_10111011 : OUT <= 0;  //58 / 187 = 0
    16'b00111010_10111100 : OUT <= 0;  //58 / 188 = 0
    16'b00111010_10111101 : OUT <= 0;  //58 / 189 = 0
    16'b00111010_10111110 : OUT <= 0;  //58 / 190 = 0
    16'b00111010_10111111 : OUT <= 0;  //58 / 191 = 0
    16'b00111010_11000000 : OUT <= 0;  //58 / 192 = 0
    16'b00111010_11000001 : OUT <= 0;  //58 / 193 = 0
    16'b00111010_11000010 : OUT <= 0;  //58 / 194 = 0
    16'b00111010_11000011 : OUT <= 0;  //58 / 195 = 0
    16'b00111010_11000100 : OUT <= 0;  //58 / 196 = 0
    16'b00111010_11000101 : OUT <= 0;  //58 / 197 = 0
    16'b00111010_11000110 : OUT <= 0;  //58 / 198 = 0
    16'b00111010_11000111 : OUT <= 0;  //58 / 199 = 0
    16'b00111010_11001000 : OUT <= 0;  //58 / 200 = 0
    16'b00111010_11001001 : OUT <= 0;  //58 / 201 = 0
    16'b00111010_11001010 : OUT <= 0;  //58 / 202 = 0
    16'b00111010_11001011 : OUT <= 0;  //58 / 203 = 0
    16'b00111010_11001100 : OUT <= 0;  //58 / 204 = 0
    16'b00111010_11001101 : OUT <= 0;  //58 / 205 = 0
    16'b00111010_11001110 : OUT <= 0;  //58 / 206 = 0
    16'b00111010_11001111 : OUT <= 0;  //58 / 207 = 0
    16'b00111010_11010000 : OUT <= 0;  //58 / 208 = 0
    16'b00111010_11010001 : OUT <= 0;  //58 / 209 = 0
    16'b00111010_11010010 : OUT <= 0;  //58 / 210 = 0
    16'b00111010_11010011 : OUT <= 0;  //58 / 211 = 0
    16'b00111010_11010100 : OUT <= 0;  //58 / 212 = 0
    16'b00111010_11010101 : OUT <= 0;  //58 / 213 = 0
    16'b00111010_11010110 : OUT <= 0;  //58 / 214 = 0
    16'b00111010_11010111 : OUT <= 0;  //58 / 215 = 0
    16'b00111010_11011000 : OUT <= 0;  //58 / 216 = 0
    16'b00111010_11011001 : OUT <= 0;  //58 / 217 = 0
    16'b00111010_11011010 : OUT <= 0;  //58 / 218 = 0
    16'b00111010_11011011 : OUT <= 0;  //58 / 219 = 0
    16'b00111010_11011100 : OUT <= 0;  //58 / 220 = 0
    16'b00111010_11011101 : OUT <= 0;  //58 / 221 = 0
    16'b00111010_11011110 : OUT <= 0;  //58 / 222 = 0
    16'b00111010_11011111 : OUT <= 0;  //58 / 223 = 0
    16'b00111010_11100000 : OUT <= 0;  //58 / 224 = 0
    16'b00111010_11100001 : OUT <= 0;  //58 / 225 = 0
    16'b00111010_11100010 : OUT <= 0;  //58 / 226 = 0
    16'b00111010_11100011 : OUT <= 0;  //58 / 227 = 0
    16'b00111010_11100100 : OUT <= 0;  //58 / 228 = 0
    16'b00111010_11100101 : OUT <= 0;  //58 / 229 = 0
    16'b00111010_11100110 : OUT <= 0;  //58 / 230 = 0
    16'b00111010_11100111 : OUT <= 0;  //58 / 231 = 0
    16'b00111010_11101000 : OUT <= 0;  //58 / 232 = 0
    16'b00111010_11101001 : OUT <= 0;  //58 / 233 = 0
    16'b00111010_11101010 : OUT <= 0;  //58 / 234 = 0
    16'b00111010_11101011 : OUT <= 0;  //58 / 235 = 0
    16'b00111010_11101100 : OUT <= 0;  //58 / 236 = 0
    16'b00111010_11101101 : OUT <= 0;  //58 / 237 = 0
    16'b00111010_11101110 : OUT <= 0;  //58 / 238 = 0
    16'b00111010_11101111 : OUT <= 0;  //58 / 239 = 0
    16'b00111010_11110000 : OUT <= 0;  //58 / 240 = 0
    16'b00111010_11110001 : OUT <= 0;  //58 / 241 = 0
    16'b00111010_11110010 : OUT <= 0;  //58 / 242 = 0
    16'b00111010_11110011 : OUT <= 0;  //58 / 243 = 0
    16'b00111010_11110100 : OUT <= 0;  //58 / 244 = 0
    16'b00111010_11110101 : OUT <= 0;  //58 / 245 = 0
    16'b00111010_11110110 : OUT <= 0;  //58 / 246 = 0
    16'b00111010_11110111 : OUT <= 0;  //58 / 247 = 0
    16'b00111010_11111000 : OUT <= 0;  //58 / 248 = 0
    16'b00111010_11111001 : OUT <= 0;  //58 / 249 = 0
    16'b00111010_11111010 : OUT <= 0;  //58 / 250 = 0
    16'b00111010_11111011 : OUT <= 0;  //58 / 251 = 0
    16'b00111010_11111100 : OUT <= 0;  //58 / 252 = 0
    16'b00111010_11111101 : OUT <= 0;  //58 / 253 = 0
    16'b00111010_11111110 : OUT <= 0;  //58 / 254 = 0
    16'b00111010_11111111 : OUT <= 0;  //58 / 255 = 0
    16'b00111011_00000000 : OUT <= 0;  //59 / 0 = 0
    16'b00111011_00000001 : OUT <= 59;  //59 / 1 = 59
    16'b00111011_00000010 : OUT <= 29;  //59 / 2 = 29
    16'b00111011_00000011 : OUT <= 19;  //59 / 3 = 19
    16'b00111011_00000100 : OUT <= 14;  //59 / 4 = 14
    16'b00111011_00000101 : OUT <= 11;  //59 / 5 = 11
    16'b00111011_00000110 : OUT <= 9;  //59 / 6 = 9
    16'b00111011_00000111 : OUT <= 8;  //59 / 7 = 8
    16'b00111011_00001000 : OUT <= 7;  //59 / 8 = 7
    16'b00111011_00001001 : OUT <= 6;  //59 / 9 = 6
    16'b00111011_00001010 : OUT <= 5;  //59 / 10 = 5
    16'b00111011_00001011 : OUT <= 5;  //59 / 11 = 5
    16'b00111011_00001100 : OUT <= 4;  //59 / 12 = 4
    16'b00111011_00001101 : OUT <= 4;  //59 / 13 = 4
    16'b00111011_00001110 : OUT <= 4;  //59 / 14 = 4
    16'b00111011_00001111 : OUT <= 3;  //59 / 15 = 3
    16'b00111011_00010000 : OUT <= 3;  //59 / 16 = 3
    16'b00111011_00010001 : OUT <= 3;  //59 / 17 = 3
    16'b00111011_00010010 : OUT <= 3;  //59 / 18 = 3
    16'b00111011_00010011 : OUT <= 3;  //59 / 19 = 3
    16'b00111011_00010100 : OUT <= 2;  //59 / 20 = 2
    16'b00111011_00010101 : OUT <= 2;  //59 / 21 = 2
    16'b00111011_00010110 : OUT <= 2;  //59 / 22 = 2
    16'b00111011_00010111 : OUT <= 2;  //59 / 23 = 2
    16'b00111011_00011000 : OUT <= 2;  //59 / 24 = 2
    16'b00111011_00011001 : OUT <= 2;  //59 / 25 = 2
    16'b00111011_00011010 : OUT <= 2;  //59 / 26 = 2
    16'b00111011_00011011 : OUT <= 2;  //59 / 27 = 2
    16'b00111011_00011100 : OUT <= 2;  //59 / 28 = 2
    16'b00111011_00011101 : OUT <= 2;  //59 / 29 = 2
    16'b00111011_00011110 : OUT <= 1;  //59 / 30 = 1
    16'b00111011_00011111 : OUT <= 1;  //59 / 31 = 1
    16'b00111011_00100000 : OUT <= 1;  //59 / 32 = 1
    16'b00111011_00100001 : OUT <= 1;  //59 / 33 = 1
    16'b00111011_00100010 : OUT <= 1;  //59 / 34 = 1
    16'b00111011_00100011 : OUT <= 1;  //59 / 35 = 1
    16'b00111011_00100100 : OUT <= 1;  //59 / 36 = 1
    16'b00111011_00100101 : OUT <= 1;  //59 / 37 = 1
    16'b00111011_00100110 : OUT <= 1;  //59 / 38 = 1
    16'b00111011_00100111 : OUT <= 1;  //59 / 39 = 1
    16'b00111011_00101000 : OUT <= 1;  //59 / 40 = 1
    16'b00111011_00101001 : OUT <= 1;  //59 / 41 = 1
    16'b00111011_00101010 : OUT <= 1;  //59 / 42 = 1
    16'b00111011_00101011 : OUT <= 1;  //59 / 43 = 1
    16'b00111011_00101100 : OUT <= 1;  //59 / 44 = 1
    16'b00111011_00101101 : OUT <= 1;  //59 / 45 = 1
    16'b00111011_00101110 : OUT <= 1;  //59 / 46 = 1
    16'b00111011_00101111 : OUT <= 1;  //59 / 47 = 1
    16'b00111011_00110000 : OUT <= 1;  //59 / 48 = 1
    16'b00111011_00110001 : OUT <= 1;  //59 / 49 = 1
    16'b00111011_00110010 : OUT <= 1;  //59 / 50 = 1
    16'b00111011_00110011 : OUT <= 1;  //59 / 51 = 1
    16'b00111011_00110100 : OUT <= 1;  //59 / 52 = 1
    16'b00111011_00110101 : OUT <= 1;  //59 / 53 = 1
    16'b00111011_00110110 : OUT <= 1;  //59 / 54 = 1
    16'b00111011_00110111 : OUT <= 1;  //59 / 55 = 1
    16'b00111011_00111000 : OUT <= 1;  //59 / 56 = 1
    16'b00111011_00111001 : OUT <= 1;  //59 / 57 = 1
    16'b00111011_00111010 : OUT <= 1;  //59 / 58 = 1
    16'b00111011_00111011 : OUT <= 1;  //59 / 59 = 1
    16'b00111011_00111100 : OUT <= 0;  //59 / 60 = 0
    16'b00111011_00111101 : OUT <= 0;  //59 / 61 = 0
    16'b00111011_00111110 : OUT <= 0;  //59 / 62 = 0
    16'b00111011_00111111 : OUT <= 0;  //59 / 63 = 0
    16'b00111011_01000000 : OUT <= 0;  //59 / 64 = 0
    16'b00111011_01000001 : OUT <= 0;  //59 / 65 = 0
    16'b00111011_01000010 : OUT <= 0;  //59 / 66 = 0
    16'b00111011_01000011 : OUT <= 0;  //59 / 67 = 0
    16'b00111011_01000100 : OUT <= 0;  //59 / 68 = 0
    16'b00111011_01000101 : OUT <= 0;  //59 / 69 = 0
    16'b00111011_01000110 : OUT <= 0;  //59 / 70 = 0
    16'b00111011_01000111 : OUT <= 0;  //59 / 71 = 0
    16'b00111011_01001000 : OUT <= 0;  //59 / 72 = 0
    16'b00111011_01001001 : OUT <= 0;  //59 / 73 = 0
    16'b00111011_01001010 : OUT <= 0;  //59 / 74 = 0
    16'b00111011_01001011 : OUT <= 0;  //59 / 75 = 0
    16'b00111011_01001100 : OUT <= 0;  //59 / 76 = 0
    16'b00111011_01001101 : OUT <= 0;  //59 / 77 = 0
    16'b00111011_01001110 : OUT <= 0;  //59 / 78 = 0
    16'b00111011_01001111 : OUT <= 0;  //59 / 79 = 0
    16'b00111011_01010000 : OUT <= 0;  //59 / 80 = 0
    16'b00111011_01010001 : OUT <= 0;  //59 / 81 = 0
    16'b00111011_01010010 : OUT <= 0;  //59 / 82 = 0
    16'b00111011_01010011 : OUT <= 0;  //59 / 83 = 0
    16'b00111011_01010100 : OUT <= 0;  //59 / 84 = 0
    16'b00111011_01010101 : OUT <= 0;  //59 / 85 = 0
    16'b00111011_01010110 : OUT <= 0;  //59 / 86 = 0
    16'b00111011_01010111 : OUT <= 0;  //59 / 87 = 0
    16'b00111011_01011000 : OUT <= 0;  //59 / 88 = 0
    16'b00111011_01011001 : OUT <= 0;  //59 / 89 = 0
    16'b00111011_01011010 : OUT <= 0;  //59 / 90 = 0
    16'b00111011_01011011 : OUT <= 0;  //59 / 91 = 0
    16'b00111011_01011100 : OUT <= 0;  //59 / 92 = 0
    16'b00111011_01011101 : OUT <= 0;  //59 / 93 = 0
    16'b00111011_01011110 : OUT <= 0;  //59 / 94 = 0
    16'b00111011_01011111 : OUT <= 0;  //59 / 95 = 0
    16'b00111011_01100000 : OUT <= 0;  //59 / 96 = 0
    16'b00111011_01100001 : OUT <= 0;  //59 / 97 = 0
    16'b00111011_01100010 : OUT <= 0;  //59 / 98 = 0
    16'b00111011_01100011 : OUT <= 0;  //59 / 99 = 0
    16'b00111011_01100100 : OUT <= 0;  //59 / 100 = 0
    16'b00111011_01100101 : OUT <= 0;  //59 / 101 = 0
    16'b00111011_01100110 : OUT <= 0;  //59 / 102 = 0
    16'b00111011_01100111 : OUT <= 0;  //59 / 103 = 0
    16'b00111011_01101000 : OUT <= 0;  //59 / 104 = 0
    16'b00111011_01101001 : OUT <= 0;  //59 / 105 = 0
    16'b00111011_01101010 : OUT <= 0;  //59 / 106 = 0
    16'b00111011_01101011 : OUT <= 0;  //59 / 107 = 0
    16'b00111011_01101100 : OUT <= 0;  //59 / 108 = 0
    16'b00111011_01101101 : OUT <= 0;  //59 / 109 = 0
    16'b00111011_01101110 : OUT <= 0;  //59 / 110 = 0
    16'b00111011_01101111 : OUT <= 0;  //59 / 111 = 0
    16'b00111011_01110000 : OUT <= 0;  //59 / 112 = 0
    16'b00111011_01110001 : OUT <= 0;  //59 / 113 = 0
    16'b00111011_01110010 : OUT <= 0;  //59 / 114 = 0
    16'b00111011_01110011 : OUT <= 0;  //59 / 115 = 0
    16'b00111011_01110100 : OUT <= 0;  //59 / 116 = 0
    16'b00111011_01110101 : OUT <= 0;  //59 / 117 = 0
    16'b00111011_01110110 : OUT <= 0;  //59 / 118 = 0
    16'b00111011_01110111 : OUT <= 0;  //59 / 119 = 0
    16'b00111011_01111000 : OUT <= 0;  //59 / 120 = 0
    16'b00111011_01111001 : OUT <= 0;  //59 / 121 = 0
    16'b00111011_01111010 : OUT <= 0;  //59 / 122 = 0
    16'b00111011_01111011 : OUT <= 0;  //59 / 123 = 0
    16'b00111011_01111100 : OUT <= 0;  //59 / 124 = 0
    16'b00111011_01111101 : OUT <= 0;  //59 / 125 = 0
    16'b00111011_01111110 : OUT <= 0;  //59 / 126 = 0
    16'b00111011_01111111 : OUT <= 0;  //59 / 127 = 0
    16'b00111011_10000000 : OUT <= 0;  //59 / 128 = 0
    16'b00111011_10000001 : OUT <= 0;  //59 / 129 = 0
    16'b00111011_10000010 : OUT <= 0;  //59 / 130 = 0
    16'b00111011_10000011 : OUT <= 0;  //59 / 131 = 0
    16'b00111011_10000100 : OUT <= 0;  //59 / 132 = 0
    16'b00111011_10000101 : OUT <= 0;  //59 / 133 = 0
    16'b00111011_10000110 : OUT <= 0;  //59 / 134 = 0
    16'b00111011_10000111 : OUT <= 0;  //59 / 135 = 0
    16'b00111011_10001000 : OUT <= 0;  //59 / 136 = 0
    16'b00111011_10001001 : OUT <= 0;  //59 / 137 = 0
    16'b00111011_10001010 : OUT <= 0;  //59 / 138 = 0
    16'b00111011_10001011 : OUT <= 0;  //59 / 139 = 0
    16'b00111011_10001100 : OUT <= 0;  //59 / 140 = 0
    16'b00111011_10001101 : OUT <= 0;  //59 / 141 = 0
    16'b00111011_10001110 : OUT <= 0;  //59 / 142 = 0
    16'b00111011_10001111 : OUT <= 0;  //59 / 143 = 0
    16'b00111011_10010000 : OUT <= 0;  //59 / 144 = 0
    16'b00111011_10010001 : OUT <= 0;  //59 / 145 = 0
    16'b00111011_10010010 : OUT <= 0;  //59 / 146 = 0
    16'b00111011_10010011 : OUT <= 0;  //59 / 147 = 0
    16'b00111011_10010100 : OUT <= 0;  //59 / 148 = 0
    16'b00111011_10010101 : OUT <= 0;  //59 / 149 = 0
    16'b00111011_10010110 : OUT <= 0;  //59 / 150 = 0
    16'b00111011_10010111 : OUT <= 0;  //59 / 151 = 0
    16'b00111011_10011000 : OUT <= 0;  //59 / 152 = 0
    16'b00111011_10011001 : OUT <= 0;  //59 / 153 = 0
    16'b00111011_10011010 : OUT <= 0;  //59 / 154 = 0
    16'b00111011_10011011 : OUT <= 0;  //59 / 155 = 0
    16'b00111011_10011100 : OUT <= 0;  //59 / 156 = 0
    16'b00111011_10011101 : OUT <= 0;  //59 / 157 = 0
    16'b00111011_10011110 : OUT <= 0;  //59 / 158 = 0
    16'b00111011_10011111 : OUT <= 0;  //59 / 159 = 0
    16'b00111011_10100000 : OUT <= 0;  //59 / 160 = 0
    16'b00111011_10100001 : OUT <= 0;  //59 / 161 = 0
    16'b00111011_10100010 : OUT <= 0;  //59 / 162 = 0
    16'b00111011_10100011 : OUT <= 0;  //59 / 163 = 0
    16'b00111011_10100100 : OUT <= 0;  //59 / 164 = 0
    16'b00111011_10100101 : OUT <= 0;  //59 / 165 = 0
    16'b00111011_10100110 : OUT <= 0;  //59 / 166 = 0
    16'b00111011_10100111 : OUT <= 0;  //59 / 167 = 0
    16'b00111011_10101000 : OUT <= 0;  //59 / 168 = 0
    16'b00111011_10101001 : OUT <= 0;  //59 / 169 = 0
    16'b00111011_10101010 : OUT <= 0;  //59 / 170 = 0
    16'b00111011_10101011 : OUT <= 0;  //59 / 171 = 0
    16'b00111011_10101100 : OUT <= 0;  //59 / 172 = 0
    16'b00111011_10101101 : OUT <= 0;  //59 / 173 = 0
    16'b00111011_10101110 : OUT <= 0;  //59 / 174 = 0
    16'b00111011_10101111 : OUT <= 0;  //59 / 175 = 0
    16'b00111011_10110000 : OUT <= 0;  //59 / 176 = 0
    16'b00111011_10110001 : OUT <= 0;  //59 / 177 = 0
    16'b00111011_10110010 : OUT <= 0;  //59 / 178 = 0
    16'b00111011_10110011 : OUT <= 0;  //59 / 179 = 0
    16'b00111011_10110100 : OUT <= 0;  //59 / 180 = 0
    16'b00111011_10110101 : OUT <= 0;  //59 / 181 = 0
    16'b00111011_10110110 : OUT <= 0;  //59 / 182 = 0
    16'b00111011_10110111 : OUT <= 0;  //59 / 183 = 0
    16'b00111011_10111000 : OUT <= 0;  //59 / 184 = 0
    16'b00111011_10111001 : OUT <= 0;  //59 / 185 = 0
    16'b00111011_10111010 : OUT <= 0;  //59 / 186 = 0
    16'b00111011_10111011 : OUT <= 0;  //59 / 187 = 0
    16'b00111011_10111100 : OUT <= 0;  //59 / 188 = 0
    16'b00111011_10111101 : OUT <= 0;  //59 / 189 = 0
    16'b00111011_10111110 : OUT <= 0;  //59 / 190 = 0
    16'b00111011_10111111 : OUT <= 0;  //59 / 191 = 0
    16'b00111011_11000000 : OUT <= 0;  //59 / 192 = 0
    16'b00111011_11000001 : OUT <= 0;  //59 / 193 = 0
    16'b00111011_11000010 : OUT <= 0;  //59 / 194 = 0
    16'b00111011_11000011 : OUT <= 0;  //59 / 195 = 0
    16'b00111011_11000100 : OUT <= 0;  //59 / 196 = 0
    16'b00111011_11000101 : OUT <= 0;  //59 / 197 = 0
    16'b00111011_11000110 : OUT <= 0;  //59 / 198 = 0
    16'b00111011_11000111 : OUT <= 0;  //59 / 199 = 0
    16'b00111011_11001000 : OUT <= 0;  //59 / 200 = 0
    16'b00111011_11001001 : OUT <= 0;  //59 / 201 = 0
    16'b00111011_11001010 : OUT <= 0;  //59 / 202 = 0
    16'b00111011_11001011 : OUT <= 0;  //59 / 203 = 0
    16'b00111011_11001100 : OUT <= 0;  //59 / 204 = 0
    16'b00111011_11001101 : OUT <= 0;  //59 / 205 = 0
    16'b00111011_11001110 : OUT <= 0;  //59 / 206 = 0
    16'b00111011_11001111 : OUT <= 0;  //59 / 207 = 0
    16'b00111011_11010000 : OUT <= 0;  //59 / 208 = 0
    16'b00111011_11010001 : OUT <= 0;  //59 / 209 = 0
    16'b00111011_11010010 : OUT <= 0;  //59 / 210 = 0
    16'b00111011_11010011 : OUT <= 0;  //59 / 211 = 0
    16'b00111011_11010100 : OUT <= 0;  //59 / 212 = 0
    16'b00111011_11010101 : OUT <= 0;  //59 / 213 = 0
    16'b00111011_11010110 : OUT <= 0;  //59 / 214 = 0
    16'b00111011_11010111 : OUT <= 0;  //59 / 215 = 0
    16'b00111011_11011000 : OUT <= 0;  //59 / 216 = 0
    16'b00111011_11011001 : OUT <= 0;  //59 / 217 = 0
    16'b00111011_11011010 : OUT <= 0;  //59 / 218 = 0
    16'b00111011_11011011 : OUT <= 0;  //59 / 219 = 0
    16'b00111011_11011100 : OUT <= 0;  //59 / 220 = 0
    16'b00111011_11011101 : OUT <= 0;  //59 / 221 = 0
    16'b00111011_11011110 : OUT <= 0;  //59 / 222 = 0
    16'b00111011_11011111 : OUT <= 0;  //59 / 223 = 0
    16'b00111011_11100000 : OUT <= 0;  //59 / 224 = 0
    16'b00111011_11100001 : OUT <= 0;  //59 / 225 = 0
    16'b00111011_11100010 : OUT <= 0;  //59 / 226 = 0
    16'b00111011_11100011 : OUT <= 0;  //59 / 227 = 0
    16'b00111011_11100100 : OUT <= 0;  //59 / 228 = 0
    16'b00111011_11100101 : OUT <= 0;  //59 / 229 = 0
    16'b00111011_11100110 : OUT <= 0;  //59 / 230 = 0
    16'b00111011_11100111 : OUT <= 0;  //59 / 231 = 0
    16'b00111011_11101000 : OUT <= 0;  //59 / 232 = 0
    16'b00111011_11101001 : OUT <= 0;  //59 / 233 = 0
    16'b00111011_11101010 : OUT <= 0;  //59 / 234 = 0
    16'b00111011_11101011 : OUT <= 0;  //59 / 235 = 0
    16'b00111011_11101100 : OUT <= 0;  //59 / 236 = 0
    16'b00111011_11101101 : OUT <= 0;  //59 / 237 = 0
    16'b00111011_11101110 : OUT <= 0;  //59 / 238 = 0
    16'b00111011_11101111 : OUT <= 0;  //59 / 239 = 0
    16'b00111011_11110000 : OUT <= 0;  //59 / 240 = 0
    16'b00111011_11110001 : OUT <= 0;  //59 / 241 = 0
    16'b00111011_11110010 : OUT <= 0;  //59 / 242 = 0
    16'b00111011_11110011 : OUT <= 0;  //59 / 243 = 0
    16'b00111011_11110100 : OUT <= 0;  //59 / 244 = 0
    16'b00111011_11110101 : OUT <= 0;  //59 / 245 = 0
    16'b00111011_11110110 : OUT <= 0;  //59 / 246 = 0
    16'b00111011_11110111 : OUT <= 0;  //59 / 247 = 0
    16'b00111011_11111000 : OUT <= 0;  //59 / 248 = 0
    16'b00111011_11111001 : OUT <= 0;  //59 / 249 = 0
    16'b00111011_11111010 : OUT <= 0;  //59 / 250 = 0
    16'b00111011_11111011 : OUT <= 0;  //59 / 251 = 0
    16'b00111011_11111100 : OUT <= 0;  //59 / 252 = 0
    16'b00111011_11111101 : OUT <= 0;  //59 / 253 = 0
    16'b00111011_11111110 : OUT <= 0;  //59 / 254 = 0
    16'b00111011_11111111 : OUT <= 0;  //59 / 255 = 0
    16'b00111100_00000000 : OUT <= 0;  //60 / 0 = 0
    16'b00111100_00000001 : OUT <= 60;  //60 / 1 = 60
    16'b00111100_00000010 : OUT <= 30;  //60 / 2 = 30
    16'b00111100_00000011 : OUT <= 20;  //60 / 3 = 20
    16'b00111100_00000100 : OUT <= 15;  //60 / 4 = 15
    16'b00111100_00000101 : OUT <= 12;  //60 / 5 = 12
    16'b00111100_00000110 : OUT <= 10;  //60 / 6 = 10
    16'b00111100_00000111 : OUT <= 8;  //60 / 7 = 8
    16'b00111100_00001000 : OUT <= 7;  //60 / 8 = 7
    16'b00111100_00001001 : OUT <= 6;  //60 / 9 = 6
    16'b00111100_00001010 : OUT <= 6;  //60 / 10 = 6
    16'b00111100_00001011 : OUT <= 5;  //60 / 11 = 5
    16'b00111100_00001100 : OUT <= 5;  //60 / 12 = 5
    16'b00111100_00001101 : OUT <= 4;  //60 / 13 = 4
    16'b00111100_00001110 : OUT <= 4;  //60 / 14 = 4
    16'b00111100_00001111 : OUT <= 4;  //60 / 15 = 4
    16'b00111100_00010000 : OUT <= 3;  //60 / 16 = 3
    16'b00111100_00010001 : OUT <= 3;  //60 / 17 = 3
    16'b00111100_00010010 : OUT <= 3;  //60 / 18 = 3
    16'b00111100_00010011 : OUT <= 3;  //60 / 19 = 3
    16'b00111100_00010100 : OUT <= 3;  //60 / 20 = 3
    16'b00111100_00010101 : OUT <= 2;  //60 / 21 = 2
    16'b00111100_00010110 : OUT <= 2;  //60 / 22 = 2
    16'b00111100_00010111 : OUT <= 2;  //60 / 23 = 2
    16'b00111100_00011000 : OUT <= 2;  //60 / 24 = 2
    16'b00111100_00011001 : OUT <= 2;  //60 / 25 = 2
    16'b00111100_00011010 : OUT <= 2;  //60 / 26 = 2
    16'b00111100_00011011 : OUT <= 2;  //60 / 27 = 2
    16'b00111100_00011100 : OUT <= 2;  //60 / 28 = 2
    16'b00111100_00011101 : OUT <= 2;  //60 / 29 = 2
    16'b00111100_00011110 : OUT <= 2;  //60 / 30 = 2
    16'b00111100_00011111 : OUT <= 1;  //60 / 31 = 1
    16'b00111100_00100000 : OUT <= 1;  //60 / 32 = 1
    16'b00111100_00100001 : OUT <= 1;  //60 / 33 = 1
    16'b00111100_00100010 : OUT <= 1;  //60 / 34 = 1
    16'b00111100_00100011 : OUT <= 1;  //60 / 35 = 1
    16'b00111100_00100100 : OUT <= 1;  //60 / 36 = 1
    16'b00111100_00100101 : OUT <= 1;  //60 / 37 = 1
    16'b00111100_00100110 : OUT <= 1;  //60 / 38 = 1
    16'b00111100_00100111 : OUT <= 1;  //60 / 39 = 1
    16'b00111100_00101000 : OUT <= 1;  //60 / 40 = 1
    16'b00111100_00101001 : OUT <= 1;  //60 / 41 = 1
    16'b00111100_00101010 : OUT <= 1;  //60 / 42 = 1
    16'b00111100_00101011 : OUT <= 1;  //60 / 43 = 1
    16'b00111100_00101100 : OUT <= 1;  //60 / 44 = 1
    16'b00111100_00101101 : OUT <= 1;  //60 / 45 = 1
    16'b00111100_00101110 : OUT <= 1;  //60 / 46 = 1
    16'b00111100_00101111 : OUT <= 1;  //60 / 47 = 1
    16'b00111100_00110000 : OUT <= 1;  //60 / 48 = 1
    16'b00111100_00110001 : OUT <= 1;  //60 / 49 = 1
    16'b00111100_00110010 : OUT <= 1;  //60 / 50 = 1
    16'b00111100_00110011 : OUT <= 1;  //60 / 51 = 1
    16'b00111100_00110100 : OUT <= 1;  //60 / 52 = 1
    16'b00111100_00110101 : OUT <= 1;  //60 / 53 = 1
    16'b00111100_00110110 : OUT <= 1;  //60 / 54 = 1
    16'b00111100_00110111 : OUT <= 1;  //60 / 55 = 1
    16'b00111100_00111000 : OUT <= 1;  //60 / 56 = 1
    16'b00111100_00111001 : OUT <= 1;  //60 / 57 = 1
    16'b00111100_00111010 : OUT <= 1;  //60 / 58 = 1
    16'b00111100_00111011 : OUT <= 1;  //60 / 59 = 1
    16'b00111100_00111100 : OUT <= 1;  //60 / 60 = 1
    16'b00111100_00111101 : OUT <= 0;  //60 / 61 = 0
    16'b00111100_00111110 : OUT <= 0;  //60 / 62 = 0
    16'b00111100_00111111 : OUT <= 0;  //60 / 63 = 0
    16'b00111100_01000000 : OUT <= 0;  //60 / 64 = 0
    16'b00111100_01000001 : OUT <= 0;  //60 / 65 = 0
    16'b00111100_01000010 : OUT <= 0;  //60 / 66 = 0
    16'b00111100_01000011 : OUT <= 0;  //60 / 67 = 0
    16'b00111100_01000100 : OUT <= 0;  //60 / 68 = 0
    16'b00111100_01000101 : OUT <= 0;  //60 / 69 = 0
    16'b00111100_01000110 : OUT <= 0;  //60 / 70 = 0
    16'b00111100_01000111 : OUT <= 0;  //60 / 71 = 0
    16'b00111100_01001000 : OUT <= 0;  //60 / 72 = 0
    16'b00111100_01001001 : OUT <= 0;  //60 / 73 = 0
    16'b00111100_01001010 : OUT <= 0;  //60 / 74 = 0
    16'b00111100_01001011 : OUT <= 0;  //60 / 75 = 0
    16'b00111100_01001100 : OUT <= 0;  //60 / 76 = 0
    16'b00111100_01001101 : OUT <= 0;  //60 / 77 = 0
    16'b00111100_01001110 : OUT <= 0;  //60 / 78 = 0
    16'b00111100_01001111 : OUT <= 0;  //60 / 79 = 0
    16'b00111100_01010000 : OUT <= 0;  //60 / 80 = 0
    16'b00111100_01010001 : OUT <= 0;  //60 / 81 = 0
    16'b00111100_01010010 : OUT <= 0;  //60 / 82 = 0
    16'b00111100_01010011 : OUT <= 0;  //60 / 83 = 0
    16'b00111100_01010100 : OUT <= 0;  //60 / 84 = 0
    16'b00111100_01010101 : OUT <= 0;  //60 / 85 = 0
    16'b00111100_01010110 : OUT <= 0;  //60 / 86 = 0
    16'b00111100_01010111 : OUT <= 0;  //60 / 87 = 0
    16'b00111100_01011000 : OUT <= 0;  //60 / 88 = 0
    16'b00111100_01011001 : OUT <= 0;  //60 / 89 = 0
    16'b00111100_01011010 : OUT <= 0;  //60 / 90 = 0
    16'b00111100_01011011 : OUT <= 0;  //60 / 91 = 0
    16'b00111100_01011100 : OUT <= 0;  //60 / 92 = 0
    16'b00111100_01011101 : OUT <= 0;  //60 / 93 = 0
    16'b00111100_01011110 : OUT <= 0;  //60 / 94 = 0
    16'b00111100_01011111 : OUT <= 0;  //60 / 95 = 0
    16'b00111100_01100000 : OUT <= 0;  //60 / 96 = 0
    16'b00111100_01100001 : OUT <= 0;  //60 / 97 = 0
    16'b00111100_01100010 : OUT <= 0;  //60 / 98 = 0
    16'b00111100_01100011 : OUT <= 0;  //60 / 99 = 0
    16'b00111100_01100100 : OUT <= 0;  //60 / 100 = 0
    16'b00111100_01100101 : OUT <= 0;  //60 / 101 = 0
    16'b00111100_01100110 : OUT <= 0;  //60 / 102 = 0
    16'b00111100_01100111 : OUT <= 0;  //60 / 103 = 0
    16'b00111100_01101000 : OUT <= 0;  //60 / 104 = 0
    16'b00111100_01101001 : OUT <= 0;  //60 / 105 = 0
    16'b00111100_01101010 : OUT <= 0;  //60 / 106 = 0
    16'b00111100_01101011 : OUT <= 0;  //60 / 107 = 0
    16'b00111100_01101100 : OUT <= 0;  //60 / 108 = 0
    16'b00111100_01101101 : OUT <= 0;  //60 / 109 = 0
    16'b00111100_01101110 : OUT <= 0;  //60 / 110 = 0
    16'b00111100_01101111 : OUT <= 0;  //60 / 111 = 0
    16'b00111100_01110000 : OUT <= 0;  //60 / 112 = 0
    16'b00111100_01110001 : OUT <= 0;  //60 / 113 = 0
    16'b00111100_01110010 : OUT <= 0;  //60 / 114 = 0
    16'b00111100_01110011 : OUT <= 0;  //60 / 115 = 0
    16'b00111100_01110100 : OUT <= 0;  //60 / 116 = 0
    16'b00111100_01110101 : OUT <= 0;  //60 / 117 = 0
    16'b00111100_01110110 : OUT <= 0;  //60 / 118 = 0
    16'b00111100_01110111 : OUT <= 0;  //60 / 119 = 0
    16'b00111100_01111000 : OUT <= 0;  //60 / 120 = 0
    16'b00111100_01111001 : OUT <= 0;  //60 / 121 = 0
    16'b00111100_01111010 : OUT <= 0;  //60 / 122 = 0
    16'b00111100_01111011 : OUT <= 0;  //60 / 123 = 0
    16'b00111100_01111100 : OUT <= 0;  //60 / 124 = 0
    16'b00111100_01111101 : OUT <= 0;  //60 / 125 = 0
    16'b00111100_01111110 : OUT <= 0;  //60 / 126 = 0
    16'b00111100_01111111 : OUT <= 0;  //60 / 127 = 0
    16'b00111100_10000000 : OUT <= 0;  //60 / 128 = 0
    16'b00111100_10000001 : OUT <= 0;  //60 / 129 = 0
    16'b00111100_10000010 : OUT <= 0;  //60 / 130 = 0
    16'b00111100_10000011 : OUT <= 0;  //60 / 131 = 0
    16'b00111100_10000100 : OUT <= 0;  //60 / 132 = 0
    16'b00111100_10000101 : OUT <= 0;  //60 / 133 = 0
    16'b00111100_10000110 : OUT <= 0;  //60 / 134 = 0
    16'b00111100_10000111 : OUT <= 0;  //60 / 135 = 0
    16'b00111100_10001000 : OUT <= 0;  //60 / 136 = 0
    16'b00111100_10001001 : OUT <= 0;  //60 / 137 = 0
    16'b00111100_10001010 : OUT <= 0;  //60 / 138 = 0
    16'b00111100_10001011 : OUT <= 0;  //60 / 139 = 0
    16'b00111100_10001100 : OUT <= 0;  //60 / 140 = 0
    16'b00111100_10001101 : OUT <= 0;  //60 / 141 = 0
    16'b00111100_10001110 : OUT <= 0;  //60 / 142 = 0
    16'b00111100_10001111 : OUT <= 0;  //60 / 143 = 0
    16'b00111100_10010000 : OUT <= 0;  //60 / 144 = 0
    16'b00111100_10010001 : OUT <= 0;  //60 / 145 = 0
    16'b00111100_10010010 : OUT <= 0;  //60 / 146 = 0
    16'b00111100_10010011 : OUT <= 0;  //60 / 147 = 0
    16'b00111100_10010100 : OUT <= 0;  //60 / 148 = 0
    16'b00111100_10010101 : OUT <= 0;  //60 / 149 = 0
    16'b00111100_10010110 : OUT <= 0;  //60 / 150 = 0
    16'b00111100_10010111 : OUT <= 0;  //60 / 151 = 0
    16'b00111100_10011000 : OUT <= 0;  //60 / 152 = 0
    16'b00111100_10011001 : OUT <= 0;  //60 / 153 = 0
    16'b00111100_10011010 : OUT <= 0;  //60 / 154 = 0
    16'b00111100_10011011 : OUT <= 0;  //60 / 155 = 0
    16'b00111100_10011100 : OUT <= 0;  //60 / 156 = 0
    16'b00111100_10011101 : OUT <= 0;  //60 / 157 = 0
    16'b00111100_10011110 : OUT <= 0;  //60 / 158 = 0
    16'b00111100_10011111 : OUT <= 0;  //60 / 159 = 0
    16'b00111100_10100000 : OUT <= 0;  //60 / 160 = 0
    16'b00111100_10100001 : OUT <= 0;  //60 / 161 = 0
    16'b00111100_10100010 : OUT <= 0;  //60 / 162 = 0
    16'b00111100_10100011 : OUT <= 0;  //60 / 163 = 0
    16'b00111100_10100100 : OUT <= 0;  //60 / 164 = 0
    16'b00111100_10100101 : OUT <= 0;  //60 / 165 = 0
    16'b00111100_10100110 : OUT <= 0;  //60 / 166 = 0
    16'b00111100_10100111 : OUT <= 0;  //60 / 167 = 0
    16'b00111100_10101000 : OUT <= 0;  //60 / 168 = 0
    16'b00111100_10101001 : OUT <= 0;  //60 / 169 = 0
    16'b00111100_10101010 : OUT <= 0;  //60 / 170 = 0
    16'b00111100_10101011 : OUT <= 0;  //60 / 171 = 0
    16'b00111100_10101100 : OUT <= 0;  //60 / 172 = 0
    16'b00111100_10101101 : OUT <= 0;  //60 / 173 = 0
    16'b00111100_10101110 : OUT <= 0;  //60 / 174 = 0
    16'b00111100_10101111 : OUT <= 0;  //60 / 175 = 0
    16'b00111100_10110000 : OUT <= 0;  //60 / 176 = 0
    16'b00111100_10110001 : OUT <= 0;  //60 / 177 = 0
    16'b00111100_10110010 : OUT <= 0;  //60 / 178 = 0
    16'b00111100_10110011 : OUT <= 0;  //60 / 179 = 0
    16'b00111100_10110100 : OUT <= 0;  //60 / 180 = 0
    16'b00111100_10110101 : OUT <= 0;  //60 / 181 = 0
    16'b00111100_10110110 : OUT <= 0;  //60 / 182 = 0
    16'b00111100_10110111 : OUT <= 0;  //60 / 183 = 0
    16'b00111100_10111000 : OUT <= 0;  //60 / 184 = 0
    16'b00111100_10111001 : OUT <= 0;  //60 / 185 = 0
    16'b00111100_10111010 : OUT <= 0;  //60 / 186 = 0
    16'b00111100_10111011 : OUT <= 0;  //60 / 187 = 0
    16'b00111100_10111100 : OUT <= 0;  //60 / 188 = 0
    16'b00111100_10111101 : OUT <= 0;  //60 / 189 = 0
    16'b00111100_10111110 : OUT <= 0;  //60 / 190 = 0
    16'b00111100_10111111 : OUT <= 0;  //60 / 191 = 0
    16'b00111100_11000000 : OUT <= 0;  //60 / 192 = 0
    16'b00111100_11000001 : OUT <= 0;  //60 / 193 = 0
    16'b00111100_11000010 : OUT <= 0;  //60 / 194 = 0
    16'b00111100_11000011 : OUT <= 0;  //60 / 195 = 0
    16'b00111100_11000100 : OUT <= 0;  //60 / 196 = 0
    16'b00111100_11000101 : OUT <= 0;  //60 / 197 = 0
    16'b00111100_11000110 : OUT <= 0;  //60 / 198 = 0
    16'b00111100_11000111 : OUT <= 0;  //60 / 199 = 0
    16'b00111100_11001000 : OUT <= 0;  //60 / 200 = 0
    16'b00111100_11001001 : OUT <= 0;  //60 / 201 = 0
    16'b00111100_11001010 : OUT <= 0;  //60 / 202 = 0
    16'b00111100_11001011 : OUT <= 0;  //60 / 203 = 0
    16'b00111100_11001100 : OUT <= 0;  //60 / 204 = 0
    16'b00111100_11001101 : OUT <= 0;  //60 / 205 = 0
    16'b00111100_11001110 : OUT <= 0;  //60 / 206 = 0
    16'b00111100_11001111 : OUT <= 0;  //60 / 207 = 0
    16'b00111100_11010000 : OUT <= 0;  //60 / 208 = 0
    16'b00111100_11010001 : OUT <= 0;  //60 / 209 = 0
    16'b00111100_11010010 : OUT <= 0;  //60 / 210 = 0
    16'b00111100_11010011 : OUT <= 0;  //60 / 211 = 0
    16'b00111100_11010100 : OUT <= 0;  //60 / 212 = 0
    16'b00111100_11010101 : OUT <= 0;  //60 / 213 = 0
    16'b00111100_11010110 : OUT <= 0;  //60 / 214 = 0
    16'b00111100_11010111 : OUT <= 0;  //60 / 215 = 0
    16'b00111100_11011000 : OUT <= 0;  //60 / 216 = 0
    16'b00111100_11011001 : OUT <= 0;  //60 / 217 = 0
    16'b00111100_11011010 : OUT <= 0;  //60 / 218 = 0
    16'b00111100_11011011 : OUT <= 0;  //60 / 219 = 0
    16'b00111100_11011100 : OUT <= 0;  //60 / 220 = 0
    16'b00111100_11011101 : OUT <= 0;  //60 / 221 = 0
    16'b00111100_11011110 : OUT <= 0;  //60 / 222 = 0
    16'b00111100_11011111 : OUT <= 0;  //60 / 223 = 0
    16'b00111100_11100000 : OUT <= 0;  //60 / 224 = 0
    16'b00111100_11100001 : OUT <= 0;  //60 / 225 = 0
    16'b00111100_11100010 : OUT <= 0;  //60 / 226 = 0
    16'b00111100_11100011 : OUT <= 0;  //60 / 227 = 0
    16'b00111100_11100100 : OUT <= 0;  //60 / 228 = 0
    16'b00111100_11100101 : OUT <= 0;  //60 / 229 = 0
    16'b00111100_11100110 : OUT <= 0;  //60 / 230 = 0
    16'b00111100_11100111 : OUT <= 0;  //60 / 231 = 0
    16'b00111100_11101000 : OUT <= 0;  //60 / 232 = 0
    16'b00111100_11101001 : OUT <= 0;  //60 / 233 = 0
    16'b00111100_11101010 : OUT <= 0;  //60 / 234 = 0
    16'b00111100_11101011 : OUT <= 0;  //60 / 235 = 0
    16'b00111100_11101100 : OUT <= 0;  //60 / 236 = 0
    16'b00111100_11101101 : OUT <= 0;  //60 / 237 = 0
    16'b00111100_11101110 : OUT <= 0;  //60 / 238 = 0
    16'b00111100_11101111 : OUT <= 0;  //60 / 239 = 0
    16'b00111100_11110000 : OUT <= 0;  //60 / 240 = 0
    16'b00111100_11110001 : OUT <= 0;  //60 / 241 = 0
    16'b00111100_11110010 : OUT <= 0;  //60 / 242 = 0
    16'b00111100_11110011 : OUT <= 0;  //60 / 243 = 0
    16'b00111100_11110100 : OUT <= 0;  //60 / 244 = 0
    16'b00111100_11110101 : OUT <= 0;  //60 / 245 = 0
    16'b00111100_11110110 : OUT <= 0;  //60 / 246 = 0
    16'b00111100_11110111 : OUT <= 0;  //60 / 247 = 0
    16'b00111100_11111000 : OUT <= 0;  //60 / 248 = 0
    16'b00111100_11111001 : OUT <= 0;  //60 / 249 = 0
    16'b00111100_11111010 : OUT <= 0;  //60 / 250 = 0
    16'b00111100_11111011 : OUT <= 0;  //60 / 251 = 0
    16'b00111100_11111100 : OUT <= 0;  //60 / 252 = 0
    16'b00111100_11111101 : OUT <= 0;  //60 / 253 = 0
    16'b00111100_11111110 : OUT <= 0;  //60 / 254 = 0
    16'b00111100_11111111 : OUT <= 0;  //60 / 255 = 0
    16'b00111101_00000000 : OUT <= 0;  //61 / 0 = 0
    16'b00111101_00000001 : OUT <= 61;  //61 / 1 = 61
    16'b00111101_00000010 : OUT <= 30;  //61 / 2 = 30
    16'b00111101_00000011 : OUT <= 20;  //61 / 3 = 20
    16'b00111101_00000100 : OUT <= 15;  //61 / 4 = 15
    16'b00111101_00000101 : OUT <= 12;  //61 / 5 = 12
    16'b00111101_00000110 : OUT <= 10;  //61 / 6 = 10
    16'b00111101_00000111 : OUT <= 8;  //61 / 7 = 8
    16'b00111101_00001000 : OUT <= 7;  //61 / 8 = 7
    16'b00111101_00001001 : OUT <= 6;  //61 / 9 = 6
    16'b00111101_00001010 : OUT <= 6;  //61 / 10 = 6
    16'b00111101_00001011 : OUT <= 5;  //61 / 11 = 5
    16'b00111101_00001100 : OUT <= 5;  //61 / 12 = 5
    16'b00111101_00001101 : OUT <= 4;  //61 / 13 = 4
    16'b00111101_00001110 : OUT <= 4;  //61 / 14 = 4
    16'b00111101_00001111 : OUT <= 4;  //61 / 15 = 4
    16'b00111101_00010000 : OUT <= 3;  //61 / 16 = 3
    16'b00111101_00010001 : OUT <= 3;  //61 / 17 = 3
    16'b00111101_00010010 : OUT <= 3;  //61 / 18 = 3
    16'b00111101_00010011 : OUT <= 3;  //61 / 19 = 3
    16'b00111101_00010100 : OUT <= 3;  //61 / 20 = 3
    16'b00111101_00010101 : OUT <= 2;  //61 / 21 = 2
    16'b00111101_00010110 : OUT <= 2;  //61 / 22 = 2
    16'b00111101_00010111 : OUT <= 2;  //61 / 23 = 2
    16'b00111101_00011000 : OUT <= 2;  //61 / 24 = 2
    16'b00111101_00011001 : OUT <= 2;  //61 / 25 = 2
    16'b00111101_00011010 : OUT <= 2;  //61 / 26 = 2
    16'b00111101_00011011 : OUT <= 2;  //61 / 27 = 2
    16'b00111101_00011100 : OUT <= 2;  //61 / 28 = 2
    16'b00111101_00011101 : OUT <= 2;  //61 / 29 = 2
    16'b00111101_00011110 : OUT <= 2;  //61 / 30 = 2
    16'b00111101_00011111 : OUT <= 1;  //61 / 31 = 1
    16'b00111101_00100000 : OUT <= 1;  //61 / 32 = 1
    16'b00111101_00100001 : OUT <= 1;  //61 / 33 = 1
    16'b00111101_00100010 : OUT <= 1;  //61 / 34 = 1
    16'b00111101_00100011 : OUT <= 1;  //61 / 35 = 1
    16'b00111101_00100100 : OUT <= 1;  //61 / 36 = 1
    16'b00111101_00100101 : OUT <= 1;  //61 / 37 = 1
    16'b00111101_00100110 : OUT <= 1;  //61 / 38 = 1
    16'b00111101_00100111 : OUT <= 1;  //61 / 39 = 1
    16'b00111101_00101000 : OUT <= 1;  //61 / 40 = 1
    16'b00111101_00101001 : OUT <= 1;  //61 / 41 = 1
    16'b00111101_00101010 : OUT <= 1;  //61 / 42 = 1
    16'b00111101_00101011 : OUT <= 1;  //61 / 43 = 1
    16'b00111101_00101100 : OUT <= 1;  //61 / 44 = 1
    16'b00111101_00101101 : OUT <= 1;  //61 / 45 = 1
    16'b00111101_00101110 : OUT <= 1;  //61 / 46 = 1
    16'b00111101_00101111 : OUT <= 1;  //61 / 47 = 1
    16'b00111101_00110000 : OUT <= 1;  //61 / 48 = 1
    16'b00111101_00110001 : OUT <= 1;  //61 / 49 = 1
    16'b00111101_00110010 : OUT <= 1;  //61 / 50 = 1
    16'b00111101_00110011 : OUT <= 1;  //61 / 51 = 1
    16'b00111101_00110100 : OUT <= 1;  //61 / 52 = 1
    16'b00111101_00110101 : OUT <= 1;  //61 / 53 = 1
    16'b00111101_00110110 : OUT <= 1;  //61 / 54 = 1
    16'b00111101_00110111 : OUT <= 1;  //61 / 55 = 1
    16'b00111101_00111000 : OUT <= 1;  //61 / 56 = 1
    16'b00111101_00111001 : OUT <= 1;  //61 / 57 = 1
    16'b00111101_00111010 : OUT <= 1;  //61 / 58 = 1
    16'b00111101_00111011 : OUT <= 1;  //61 / 59 = 1
    16'b00111101_00111100 : OUT <= 1;  //61 / 60 = 1
    16'b00111101_00111101 : OUT <= 1;  //61 / 61 = 1
    16'b00111101_00111110 : OUT <= 0;  //61 / 62 = 0
    16'b00111101_00111111 : OUT <= 0;  //61 / 63 = 0
    16'b00111101_01000000 : OUT <= 0;  //61 / 64 = 0
    16'b00111101_01000001 : OUT <= 0;  //61 / 65 = 0
    16'b00111101_01000010 : OUT <= 0;  //61 / 66 = 0
    16'b00111101_01000011 : OUT <= 0;  //61 / 67 = 0
    16'b00111101_01000100 : OUT <= 0;  //61 / 68 = 0
    16'b00111101_01000101 : OUT <= 0;  //61 / 69 = 0
    16'b00111101_01000110 : OUT <= 0;  //61 / 70 = 0
    16'b00111101_01000111 : OUT <= 0;  //61 / 71 = 0
    16'b00111101_01001000 : OUT <= 0;  //61 / 72 = 0
    16'b00111101_01001001 : OUT <= 0;  //61 / 73 = 0
    16'b00111101_01001010 : OUT <= 0;  //61 / 74 = 0
    16'b00111101_01001011 : OUT <= 0;  //61 / 75 = 0
    16'b00111101_01001100 : OUT <= 0;  //61 / 76 = 0
    16'b00111101_01001101 : OUT <= 0;  //61 / 77 = 0
    16'b00111101_01001110 : OUT <= 0;  //61 / 78 = 0
    16'b00111101_01001111 : OUT <= 0;  //61 / 79 = 0
    16'b00111101_01010000 : OUT <= 0;  //61 / 80 = 0
    16'b00111101_01010001 : OUT <= 0;  //61 / 81 = 0
    16'b00111101_01010010 : OUT <= 0;  //61 / 82 = 0
    16'b00111101_01010011 : OUT <= 0;  //61 / 83 = 0
    16'b00111101_01010100 : OUT <= 0;  //61 / 84 = 0
    16'b00111101_01010101 : OUT <= 0;  //61 / 85 = 0
    16'b00111101_01010110 : OUT <= 0;  //61 / 86 = 0
    16'b00111101_01010111 : OUT <= 0;  //61 / 87 = 0
    16'b00111101_01011000 : OUT <= 0;  //61 / 88 = 0
    16'b00111101_01011001 : OUT <= 0;  //61 / 89 = 0
    16'b00111101_01011010 : OUT <= 0;  //61 / 90 = 0
    16'b00111101_01011011 : OUT <= 0;  //61 / 91 = 0
    16'b00111101_01011100 : OUT <= 0;  //61 / 92 = 0
    16'b00111101_01011101 : OUT <= 0;  //61 / 93 = 0
    16'b00111101_01011110 : OUT <= 0;  //61 / 94 = 0
    16'b00111101_01011111 : OUT <= 0;  //61 / 95 = 0
    16'b00111101_01100000 : OUT <= 0;  //61 / 96 = 0
    16'b00111101_01100001 : OUT <= 0;  //61 / 97 = 0
    16'b00111101_01100010 : OUT <= 0;  //61 / 98 = 0
    16'b00111101_01100011 : OUT <= 0;  //61 / 99 = 0
    16'b00111101_01100100 : OUT <= 0;  //61 / 100 = 0
    16'b00111101_01100101 : OUT <= 0;  //61 / 101 = 0
    16'b00111101_01100110 : OUT <= 0;  //61 / 102 = 0
    16'b00111101_01100111 : OUT <= 0;  //61 / 103 = 0
    16'b00111101_01101000 : OUT <= 0;  //61 / 104 = 0
    16'b00111101_01101001 : OUT <= 0;  //61 / 105 = 0
    16'b00111101_01101010 : OUT <= 0;  //61 / 106 = 0
    16'b00111101_01101011 : OUT <= 0;  //61 / 107 = 0
    16'b00111101_01101100 : OUT <= 0;  //61 / 108 = 0
    16'b00111101_01101101 : OUT <= 0;  //61 / 109 = 0
    16'b00111101_01101110 : OUT <= 0;  //61 / 110 = 0
    16'b00111101_01101111 : OUT <= 0;  //61 / 111 = 0
    16'b00111101_01110000 : OUT <= 0;  //61 / 112 = 0
    16'b00111101_01110001 : OUT <= 0;  //61 / 113 = 0
    16'b00111101_01110010 : OUT <= 0;  //61 / 114 = 0
    16'b00111101_01110011 : OUT <= 0;  //61 / 115 = 0
    16'b00111101_01110100 : OUT <= 0;  //61 / 116 = 0
    16'b00111101_01110101 : OUT <= 0;  //61 / 117 = 0
    16'b00111101_01110110 : OUT <= 0;  //61 / 118 = 0
    16'b00111101_01110111 : OUT <= 0;  //61 / 119 = 0
    16'b00111101_01111000 : OUT <= 0;  //61 / 120 = 0
    16'b00111101_01111001 : OUT <= 0;  //61 / 121 = 0
    16'b00111101_01111010 : OUT <= 0;  //61 / 122 = 0
    16'b00111101_01111011 : OUT <= 0;  //61 / 123 = 0
    16'b00111101_01111100 : OUT <= 0;  //61 / 124 = 0
    16'b00111101_01111101 : OUT <= 0;  //61 / 125 = 0
    16'b00111101_01111110 : OUT <= 0;  //61 / 126 = 0
    16'b00111101_01111111 : OUT <= 0;  //61 / 127 = 0
    16'b00111101_10000000 : OUT <= 0;  //61 / 128 = 0
    16'b00111101_10000001 : OUT <= 0;  //61 / 129 = 0
    16'b00111101_10000010 : OUT <= 0;  //61 / 130 = 0
    16'b00111101_10000011 : OUT <= 0;  //61 / 131 = 0
    16'b00111101_10000100 : OUT <= 0;  //61 / 132 = 0
    16'b00111101_10000101 : OUT <= 0;  //61 / 133 = 0
    16'b00111101_10000110 : OUT <= 0;  //61 / 134 = 0
    16'b00111101_10000111 : OUT <= 0;  //61 / 135 = 0
    16'b00111101_10001000 : OUT <= 0;  //61 / 136 = 0
    16'b00111101_10001001 : OUT <= 0;  //61 / 137 = 0
    16'b00111101_10001010 : OUT <= 0;  //61 / 138 = 0
    16'b00111101_10001011 : OUT <= 0;  //61 / 139 = 0
    16'b00111101_10001100 : OUT <= 0;  //61 / 140 = 0
    16'b00111101_10001101 : OUT <= 0;  //61 / 141 = 0
    16'b00111101_10001110 : OUT <= 0;  //61 / 142 = 0
    16'b00111101_10001111 : OUT <= 0;  //61 / 143 = 0
    16'b00111101_10010000 : OUT <= 0;  //61 / 144 = 0
    16'b00111101_10010001 : OUT <= 0;  //61 / 145 = 0
    16'b00111101_10010010 : OUT <= 0;  //61 / 146 = 0
    16'b00111101_10010011 : OUT <= 0;  //61 / 147 = 0
    16'b00111101_10010100 : OUT <= 0;  //61 / 148 = 0
    16'b00111101_10010101 : OUT <= 0;  //61 / 149 = 0
    16'b00111101_10010110 : OUT <= 0;  //61 / 150 = 0
    16'b00111101_10010111 : OUT <= 0;  //61 / 151 = 0
    16'b00111101_10011000 : OUT <= 0;  //61 / 152 = 0
    16'b00111101_10011001 : OUT <= 0;  //61 / 153 = 0
    16'b00111101_10011010 : OUT <= 0;  //61 / 154 = 0
    16'b00111101_10011011 : OUT <= 0;  //61 / 155 = 0
    16'b00111101_10011100 : OUT <= 0;  //61 / 156 = 0
    16'b00111101_10011101 : OUT <= 0;  //61 / 157 = 0
    16'b00111101_10011110 : OUT <= 0;  //61 / 158 = 0
    16'b00111101_10011111 : OUT <= 0;  //61 / 159 = 0
    16'b00111101_10100000 : OUT <= 0;  //61 / 160 = 0
    16'b00111101_10100001 : OUT <= 0;  //61 / 161 = 0
    16'b00111101_10100010 : OUT <= 0;  //61 / 162 = 0
    16'b00111101_10100011 : OUT <= 0;  //61 / 163 = 0
    16'b00111101_10100100 : OUT <= 0;  //61 / 164 = 0
    16'b00111101_10100101 : OUT <= 0;  //61 / 165 = 0
    16'b00111101_10100110 : OUT <= 0;  //61 / 166 = 0
    16'b00111101_10100111 : OUT <= 0;  //61 / 167 = 0
    16'b00111101_10101000 : OUT <= 0;  //61 / 168 = 0
    16'b00111101_10101001 : OUT <= 0;  //61 / 169 = 0
    16'b00111101_10101010 : OUT <= 0;  //61 / 170 = 0
    16'b00111101_10101011 : OUT <= 0;  //61 / 171 = 0
    16'b00111101_10101100 : OUT <= 0;  //61 / 172 = 0
    16'b00111101_10101101 : OUT <= 0;  //61 / 173 = 0
    16'b00111101_10101110 : OUT <= 0;  //61 / 174 = 0
    16'b00111101_10101111 : OUT <= 0;  //61 / 175 = 0
    16'b00111101_10110000 : OUT <= 0;  //61 / 176 = 0
    16'b00111101_10110001 : OUT <= 0;  //61 / 177 = 0
    16'b00111101_10110010 : OUT <= 0;  //61 / 178 = 0
    16'b00111101_10110011 : OUT <= 0;  //61 / 179 = 0
    16'b00111101_10110100 : OUT <= 0;  //61 / 180 = 0
    16'b00111101_10110101 : OUT <= 0;  //61 / 181 = 0
    16'b00111101_10110110 : OUT <= 0;  //61 / 182 = 0
    16'b00111101_10110111 : OUT <= 0;  //61 / 183 = 0
    16'b00111101_10111000 : OUT <= 0;  //61 / 184 = 0
    16'b00111101_10111001 : OUT <= 0;  //61 / 185 = 0
    16'b00111101_10111010 : OUT <= 0;  //61 / 186 = 0
    16'b00111101_10111011 : OUT <= 0;  //61 / 187 = 0
    16'b00111101_10111100 : OUT <= 0;  //61 / 188 = 0
    16'b00111101_10111101 : OUT <= 0;  //61 / 189 = 0
    16'b00111101_10111110 : OUT <= 0;  //61 / 190 = 0
    16'b00111101_10111111 : OUT <= 0;  //61 / 191 = 0
    16'b00111101_11000000 : OUT <= 0;  //61 / 192 = 0
    16'b00111101_11000001 : OUT <= 0;  //61 / 193 = 0
    16'b00111101_11000010 : OUT <= 0;  //61 / 194 = 0
    16'b00111101_11000011 : OUT <= 0;  //61 / 195 = 0
    16'b00111101_11000100 : OUT <= 0;  //61 / 196 = 0
    16'b00111101_11000101 : OUT <= 0;  //61 / 197 = 0
    16'b00111101_11000110 : OUT <= 0;  //61 / 198 = 0
    16'b00111101_11000111 : OUT <= 0;  //61 / 199 = 0
    16'b00111101_11001000 : OUT <= 0;  //61 / 200 = 0
    16'b00111101_11001001 : OUT <= 0;  //61 / 201 = 0
    16'b00111101_11001010 : OUT <= 0;  //61 / 202 = 0
    16'b00111101_11001011 : OUT <= 0;  //61 / 203 = 0
    16'b00111101_11001100 : OUT <= 0;  //61 / 204 = 0
    16'b00111101_11001101 : OUT <= 0;  //61 / 205 = 0
    16'b00111101_11001110 : OUT <= 0;  //61 / 206 = 0
    16'b00111101_11001111 : OUT <= 0;  //61 / 207 = 0
    16'b00111101_11010000 : OUT <= 0;  //61 / 208 = 0
    16'b00111101_11010001 : OUT <= 0;  //61 / 209 = 0
    16'b00111101_11010010 : OUT <= 0;  //61 / 210 = 0
    16'b00111101_11010011 : OUT <= 0;  //61 / 211 = 0
    16'b00111101_11010100 : OUT <= 0;  //61 / 212 = 0
    16'b00111101_11010101 : OUT <= 0;  //61 / 213 = 0
    16'b00111101_11010110 : OUT <= 0;  //61 / 214 = 0
    16'b00111101_11010111 : OUT <= 0;  //61 / 215 = 0
    16'b00111101_11011000 : OUT <= 0;  //61 / 216 = 0
    16'b00111101_11011001 : OUT <= 0;  //61 / 217 = 0
    16'b00111101_11011010 : OUT <= 0;  //61 / 218 = 0
    16'b00111101_11011011 : OUT <= 0;  //61 / 219 = 0
    16'b00111101_11011100 : OUT <= 0;  //61 / 220 = 0
    16'b00111101_11011101 : OUT <= 0;  //61 / 221 = 0
    16'b00111101_11011110 : OUT <= 0;  //61 / 222 = 0
    16'b00111101_11011111 : OUT <= 0;  //61 / 223 = 0
    16'b00111101_11100000 : OUT <= 0;  //61 / 224 = 0
    16'b00111101_11100001 : OUT <= 0;  //61 / 225 = 0
    16'b00111101_11100010 : OUT <= 0;  //61 / 226 = 0
    16'b00111101_11100011 : OUT <= 0;  //61 / 227 = 0
    16'b00111101_11100100 : OUT <= 0;  //61 / 228 = 0
    16'b00111101_11100101 : OUT <= 0;  //61 / 229 = 0
    16'b00111101_11100110 : OUT <= 0;  //61 / 230 = 0
    16'b00111101_11100111 : OUT <= 0;  //61 / 231 = 0
    16'b00111101_11101000 : OUT <= 0;  //61 / 232 = 0
    16'b00111101_11101001 : OUT <= 0;  //61 / 233 = 0
    16'b00111101_11101010 : OUT <= 0;  //61 / 234 = 0
    16'b00111101_11101011 : OUT <= 0;  //61 / 235 = 0
    16'b00111101_11101100 : OUT <= 0;  //61 / 236 = 0
    16'b00111101_11101101 : OUT <= 0;  //61 / 237 = 0
    16'b00111101_11101110 : OUT <= 0;  //61 / 238 = 0
    16'b00111101_11101111 : OUT <= 0;  //61 / 239 = 0
    16'b00111101_11110000 : OUT <= 0;  //61 / 240 = 0
    16'b00111101_11110001 : OUT <= 0;  //61 / 241 = 0
    16'b00111101_11110010 : OUT <= 0;  //61 / 242 = 0
    16'b00111101_11110011 : OUT <= 0;  //61 / 243 = 0
    16'b00111101_11110100 : OUT <= 0;  //61 / 244 = 0
    16'b00111101_11110101 : OUT <= 0;  //61 / 245 = 0
    16'b00111101_11110110 : OUT <= 0;  //61 / 246 = 0
    16'b00111101_11110111 : OUT <= 0;  //61 / 247 = 0
    16'b00111101_11111000 : OUT <= 0;  //61 / 248 = 0
    16'b00111101_11111001 : OUT <= 0;  //61 / 249 = 0
    16'b00111101_11111010 : OUT <= 0;  //61 / 250 = 0
    16'b00111101_11111011 : OUT <= 0;  //61 / 251 = 0
    16'b00111101_11111100 : OUT <= 0;  //61 / 252 = 0
    16'b00111101_11111101 : OUT <= 0;  //61 / 253 = 0
    16'b00111101_11111110 : OUT <= 0;  //61 / 254 = 0
    16'b00111101_11111111 : OUT <= 0;  //61 / 255 = 0
    16'b00111110_00000000 : OUT <= 0;  //62 / 0 = 0
    16'b00111110_00000001 : OUT <= 62;  //62 / 1 = 62
    16'b00111110_00000010 : OUT <= 31;  //62 / 2 = 31
    16'b00111110_00000011 : OUT <= 20;  //62 / 3 = 20
    16'b00111110_00000100 : OUT <= 15;  //62 / 4 = 15
    16'b00111110_00000101 : OUT <= 12;  //62 / 5 = 12
    16'b00111110_00000110 : OUT <= 10;  //62 / 6 = 10
    16'b00111110_00000111 : OUT <= 8;  //62 / 7 = 8
    16'b00111110_00001000 : OUT <= 7;  //62 / 8 = 7
    16'b00111110_00001001 : OUT <= 6;  //62 / 9 = 6
    16'b00111110_00001010 : OUT <= 6;  //62 / 10 = 6
    16'b00111110_00001011 : OUT <= 5;  //62 / 11 = 5
    16'b00111110_00001100 : OUT <= 5;  //62 / 12 = 5
    16'b00111110_00001101 : OUT <= 4;  //62 / 13 = 4
    16'b00111110_00001110 : OUT <= 4;  //62 / 14 = 4
    16'b00111110_00001111 : OUT <= 4;  //62 / 15 = 4
    16'b00111110_00010000 : OUT <= 3;  //62 / 16 = 3
    16'b00111110_00010001 : OUT <= 3;  //62 / 17 = 3
    16'b00111110_00010010 : OUT <= 3;  //62 / 18 = 3
    16'b00111110_00010011 : OUT <= 3;  //62 / 19 = 3
    16'b00111110_00010100 : OUT <= 3;  //62 / 20 = 3
    16'b00111110_00010101 : OUT <= 2;  //62 / 21 = 2
    16'b00111110_00010110 : OUT <= 2;  //62 / 22 = 2
    16'b00111110_00010111 : OUT <= 2;  //62 / 23 = 2
    16'b00111110_00011000 : OUT <= 2;  //62 / 24 = 2
    16'b00111110_00011001 : OUT <= 2;  //62 / 25 = 2
    16'b00111110_00011010 : OUT <= 2;  //62 / 26 = 2
    16'b00111110_00011011 : OUT <= 2;  //62 / 27 = 2
    16'b00111110_00011100 : OUT <= 2;  //62 / 28 = 2
    16'b00111110_00011101 : OUT <= 2;  //62 / 29 = 2
    16'b00111110_00011110 : OUT <= 2;  //62 / 30 = 2
    16'b00111110_00011111 : OUT <= 2;  //62 / 31 = 2
    16'b00111110_00100000 : OUT <= 1;  //62 / 32 = 1
    16'b00111110_00100001 : OUT <= 1;  //62 / 33 = 1
    16'b00111110_00100010 : OUT <= 1;  //62 / 34 = 1
    16'b00111110_00100011 : OUT <= 1;  //62 / 35 = 1
    16'b00111110_00100100 : OUT <= 1;  //62 / 36 = 1
    16'b00111110_00100101 : OUT <= 1;  //62 / 37 = 1
    16'b00111110_00100110 : OUT <= 1;  //62 / 38 = 1
    16'b00111110_00100111 : OUT <= 1;  //62 / 39 = 1
    16'b00111110_00101000 : OUT <= 1;  //62 / 40 = 1
    16'b00111110_00101001 : OUT <= 1;  //62 / 41 = 1
    16'b00111110_00101010 : OUT <= 1;  //62 / 42 = 1
    16'b00111110_00101011 : OUT <= 1;  //62 / 43 = 1
    16'b00111110_00101100 : OUT <= 1;  //62 / 44 = 1
    16'b00111110_00101101 : OUT <= 1;  //62 / 45 = 1
    16'b00111110_00101110 : OUT <= 1;  //62 / 46 = 1
    16'b00111110_00101111 : OUT <= 1;  //62 / 47 = 1
    16'b00111110_00110000 : OUT <= 1;  //62 / 48 = 1
    16'b00111110_00110001 : OUT <= 1;  //62 / 49 = 1
    16'b00111110_00110010 : OUT <= 1;  //62 / 50 = 1
    16'b00111110_00110011 : OUT <= 1;  //62 / 51 = 1
    16'b00111110_00110100 : OUT <= 1;  //62 / 52 = 1
    16'b00111110_00110101 : OUT <= 1;  //62 / 53 = 1
    16'b00111110_00110110 : OUT <= 1;  //62 / 54 = 1
    16'b00111110_00110111 : OUT <= 1;  //62 / 55 = 1
    16'b00111110_00111000 : OUT <= 1;  //62 / 56 = 1
    16'b00111110_00111001 : OUT <= 1;  //62 / 57 = 1
    16'b00111110_00111010 : OUT <= 1;  //62 / 58 = 1
    16'b00111110_00111011 : OUT <= 1;  //62 / 59 = 1
    16'b00111110_00111100 : OUT <= 1;  //62 / 60 = 1
    16'b00111110_00111101 : OUT <= 1;  //62 / 61 = 1
    16'b00111110_00111110 : OUT <= 1;  //62 / 62 = 1
    16'b00111110_00111111 : OUT <= 0;  //62 / 63 = 0
    16'b00111110_01000000 : OUT <= 0;  //62 / 64 = 0
    16'b00111110_01000001 : OUT <= 0;  //62 / 65 = 0
    16'b00111110_01000010 : OUT <= 0;  //62 / 66 = 0
    16'b00111110_01000011 : OUT <= 0;  //62 / 67 = 0
    16'b00111110_01000100 : OUT <= 0;  //62 / 68 = 0
    16'b00111110_01000101 : OUT <= 0;  //62 / 69 = 0
    16'b00111110_01000110 : OUT <= 0;  //62 / 70 = 0
    16'b00111110_01000111 : OUT <= 0;  //62 / 71 = 0
    16'b00111110_01001000 : OUT <= 0;  //62 / 72 = 0
    16'b00111110_01001001 : OUT <= 0;  //62 / 73 = 0
    16'b00111110_01001010 : OUT <= 0;  //62 / 74 = 0
    16'b00111110_01001011 : OUT <= 0;  //62 / 75 = 0
    16'b00111110_01001100 : OUT <= 0;  //62 / 76 = 0
    16'b00111110_01001101 : OUT <= 0;  //62 / 77 = 0
    16'b00111110_01001110 : OUT <= 0;  //62 / 78 = 0
    16'b00111110_01001111 : OUT <= 0;  //62 / 79 = 0
    16'b00111110_01010000 : OUT <= 0;  //62 / 80 = 0
    16'b00111110_01010001 : OUT <= 0;  //62 / 81 = 0
    16'b00111110_01010010 : OUT <= 0;  //62 / 82 = 0
    16'b00111110_01010011 : OUT <= 0;  //62 / 83 = 0
    16'b00111110_01010100 : OUT <= 0;  //62 / 84 = 0
    16'b00111110_01010101 : OUT <= 0;  //62 / 85 = 0
    16'b00111110_01010110 : OUT <= 0;  //62 / 86 = 0
    16'b00111110_01010111 : OUT <= 0;  //62 / 87 = 0
    16'b00111110_01011000 : OUT <= 0;  //62 / 88 = 0
    16'b00111110_01011001 : OUT <= 0;  //62 / 89 = 0
    16'b00111110_01011010 : OUT <= 0;  //62 / 90 = 0
    16'b00111110_01011011 : OUT <= 0;  //62 / 91 = 0
    16'b00111110_01011100 : OUT <= 0;  //62 / 92 = 0
    16'b00111110_01011101 : OUT <= 0;  //62 / 93 = 0
    16'b00111110_01011110 : OUT <= 0;  //62 / 94 = 0
    16'b00111110_01011111 : OUT <= 0;  //62 / 95 = 0
    16'b00111110_01100000 : OUT <= 0;  //62 / 96 = 0
    16'b00111110_01100001 : OUT <= 0;  //62 / 97 = 0
    16'b00111110_01100010 : OUT <= 0;  //62 / 98 = 0
    16'b00111110_01100011 : OUT <= 0;  //62 / 99 = 0
    16'b00111110_01100100 : OUT <= 0;  //62 / 100 = 0
    16'b00111110_01100101 : OUT <= 0;  //62 / 101 = 0
    16'b00111110_01100110 : OUT <= 0;  //62 / 102 = 0
    16'b00111110_01100111 : OUT <= 0;  //62 / 103 = 0
    16'b00111110_01101000 : OUT <= 0;  //62 / 104 = 0
    16'b00111110_01101001 : OUT <= 0;  //62 / 105 = 0
    16'b00111110_01101010 : OUT <= 0;  //62 / 106 = 0
    16'b00111110_01101011 : OUT <= 0;  //62 / 107 = 0
    16'b00111110_01101100 : OUT <= 0;  //62 / 108 = 0
    16'b00111110_01101101 : OUT <= 0;  //62 / 109 = 0
    16'b00111110_01101110 : OUT <= 0;  //62 / 110 = 0
    16'b00111110_01101111 : OUT <= 0;  //62 / 111 = 0
    16'b00111110_01110000 : OUT <= 0;  //62 / 112 = 0
    16'b00111110_01110001 : OUT <= 0;  //62 / 113 = 0
    16'b00111110_01110010 : OUT <= 0;  //62 / 114 = 0
    16'b00111110_01110011 : OUT <= 0;  //62 / 115 = 0
    16'b00111110_01110100 : OUT <= 0;  //62 / 116 = 0
    16'b00111110_01110101 : OUT <= 0;  //62 / 117 = 0
    16'b00111110_01110110 : OUT <= 0;  //62 / 118 = 0
    16'b00111110_01110111 : OUT <= 0;  //62 / 119 = 0
    16'b00111110_01111000 : OUT <= 0;  //62 / 120 = 0
    16'b00111110_01111001 : OUT <= 0;  //62 / 121 = 0
    16'b00111110_01111010 : OUT <= 0;  //62 / 122 = 0
    16'b00111110_01111011 : OUT <= 0;  //62 / 123 = 0
    16'b00111110_01111100 : OUT <= 0;  //62 / 124 = 0
    16'b00111110_01111101 : OUT <= 0;  //62 / 125 = 0
    16'b00111110_01111110 : OUT <= 0;  //62 / 126 = 0
    16'b00111110_01111111 : OUT <= 0;  //62 / 127 = 0
    16'b00111110_10000000 : OUT <= 0;  //62 / 128 = 0
    16'b00111110_10000001 : OUT <= 0;  //62 / 129 = 0
    16'b00111110_10000010 : OUT <= 0;  //62 / 130 = 0
    16'b00111110_10000011 : OUT <= 0;  //62 / 131 = 0
    16'b00111110_10000100 : OUT <= 0;  //62 / 132 = 0
    16'b00111110_10000101 : OUT <= 0;  //62 / 133 = 0
    16'b00111110_10000110 : OUT <= 0;  //62 / 134 = 0
    16'b00111110_10000111 : OUT <= 0;  //62 / 135 = 0
    16'b00111110_10001000 : OUT <= 0;  //62 / 136 = 0
    16'b00111110_10001001 : OUT <= 0;  //62 / 137 = 0
    16'b00111110_10001010 : OUT <= 0;  //62 / 138 = 0
    16'b00111110_10001011 : OUT <= 0;  //62 / 139 = 0
    16'b00111110_10001100 : OUT <= 0;  //62 / 140 = 0
    16'b00111110_10001101 : OUT <= 0;  //62 / 141 = 0
    16'b00111110_10001110 : OUT <= 0;  //62 / 142 = 0
    16'b00111110_10001111 : OUT <= 0;  //62 / 143 = 0
    16'b00111110_10010000 : OUT <= 0;  //62 / 144 = 0
    16'b00111110_10010001 : OUT <= 0;  //62 / 145 = 0
    16'b00111110_10010010 : OUT <= 0;  //62 / 146 = 0
    16'b00111110_10010011 : OUT <= 0;  //62 / 147 = 0
    16'b00111110_10010100 : OUT <= 0;  //62 / 148 = 0
    16'b00111110_10010101 : OUT <= 0;  //62 / 149 = 0
    16'b00111110_10010110 : OUT <= 0;  //62 / 150 = 0
    16'b00111110_10010111 : OUT <= 0;  //62 / 151 = 0
    16'b00111110_10011000 : OUT <= 0;  //62 / 152 = 0
    16'b00111110_10011001 : OUT <= 0;  //62 / 153 = 0
    16'b00111110_10011010 : OUT <= 0;  //62 / 154 = 0
    16'b00111110_10011011 : OUT <= 0;  //62 / 155 = 0
    16'b00111110_10011100 : OUT <= 0;  //62 / 156 = 0
    16'b00111110_10011101 : OUT <= 0;  //62 / 157 = 0
    16'b00111110_10011110 : OUT <= 0;  //62 / 158 = 0
    16'b00111110_10011111 : OUT <= 0;  //62 / 159 = 0
    16'b00111110_10100000 : OUT <= 0;  //62 / 160 = 0
    16'b00111110_10100001 : OUT <= 0;  //62 / 161 = 0
    16'b00111110_10100010 : OUT <= 0;  //62 / 162 = 0
    16'b00111110_10100011 : OUT <= 0;  //62 / 163 = 0
    16'b00111110_10100100 : OUT <= 0;  //62 / 164 = 0
    16'b00111110_10100101 : OUT <= 0;  //62 / 165 = 0
    16'b00111110_10100110 : OUT <= 0;  //62 / 166 = 0
    16'b00111110_10100111 : OUT <= 0;  //62 / 167 = 0
    16'b00111110_10101000 : OUT <= 0;  //62 / 168 = 0
    16'b00111110_10101001 : OUT <= 0;  //62 / 169 = 0
    16'b00111110_10101010 : OUT <= 0;  //62 / 170 = 0
    16'b00111110_10101011 : OUT <= 0;  //62 / 171 = 0
    16'b00111110_10101100 : OUT <= 0;  //62 / 172 = 0
    16'b00111110_10101101 : OUT <= 0;  //62 / 173 = 0
    16'b00111110_10101110 : OUT <= 0;  //62 / 174 = 0
    16'b00111110_10101111 : OUT <= 0;  //62 / 175 = 0
    16'b00111110_10110000 : OUT <= 0;  //62 / 176 = 0
    16'b00111110_10110001 : OUT <= 0;  //62 / 177 = 0
    16'b00111110_10110010 : OUT <= 0;  //62 / 178 = 0
    16'b00111110_10110011 : OUT <= 0;  //62 / 179 = 0
    16'b00111110_10110100 : OUT <= 0;  //62 / 180 = 0
    16'b00111110_10110101 : OUT <= 0;  //62 / 181 = 0
    16'b00111110_10110110 : OUT <= 0;  //62 / 182 = 0
    16'b00111110_10110111 : OUT <= 0;  //62 / 183 = 0
    16'b00111110_10111000 : OUT <= 0;  //62 / 184 = 0
    16'b00111110_10111001 : OUT <= 0;  //62 / 185 = 0
    16'b00111110_10111010 : OUT <= 0;  //62 / 186 = 0
    16'b00111110_10111011 : OUT <= 0;  //62 / 187 = 0
    16'b00111110_10111100 : OUT <= 0;  //62 / 188 = 0
    16'b00111110_10111101 : OUT <= 0;  //62 / 189 = 0
    16'b00111110_10111110 : OUT <= 0;  //62 / 190 = 0
    16'b00111110_10111111 : OUT <= 0;  //62 / 191 = 0
    16'b00111110_11000000 : OUT <= 0;  //62 / 192 = 0
    16'b00111110_11000001 : OUT <= 0;  //62 / 193 = 0
    16'b00111110_11000010 : OUT <= 0;  //62 / 194 = 0
    16'b00111110_11000011 : OUT <= 0;  //62 / 195 = 0
    16'b00111110_11000100 : OUT <= 0;  //62 / 196 = 0
    16'b00111110_11000101 : OUT <= 0;  //62 / 197 = 0
    16'b00111110_11000110 : OUT <= 0;  //62 / 198 = 0
    16'b00111110_11000111 : OUT <= 0;  //62 / 199 = 0
    16'b00111110_11001000 : OUT <= 0;  //62 / 200 = 0
    16'b00111110_11001001 : OUT <= 0;  //62 / 201 = 0
    16'b00111110_11001010 : OUT <= 0;  //62 / 202 = 0
    16'b00111110_11001011 : OUT <= 0;  //62 / 203 = 0
    16'b00111110_11001100 : OUT <= 0;  //62 / 204 = 0
    16'b00111110_11001101 : OUT <= 0;  //62 / 205 = 0
    16'b00111110_11001110 : OUT <= 0;  //62 / 206 = 0
    16'b00111110_11001111 : OUT <= 0;  //62 / 207 = 0
    16'b00111110_11010000 : OUT <= 0;  //62 / 208 = 0
    16'b00111110_11010001 : OUT <= 0;  //62 / 209 = 0
    16'b00111110_11010010 : OUT <= 0;  //62 / 210 = 0
    16'b00111110_11010011 : OUT <= 0;  //62 / 211 = 0
    16'b00111110_11010100 : OUT <= 0;  //62 / 212 = 0
    16'b00111110_11010101 : OUT <= 0;  //62 / 213 = 0
    16'b00111110_11010110 : OUT <= 0;  //62 / 214 = 0
    16'b00111110_11010111 : OUT <= 0;  //62 / 215 = 0
    16'b00111110_11011000 : OUT <= 0;  //62 / 216 = 0
    16'b00111110_11011001 : OUT <= 0;  //62 / 217 = 0
    16'b00111110_11011010 : OUT <= 0;  //62 / 218 = 0
    16'b00111110_11011011 : OUT <= 0;  //62 / 219 = 0
    16'b00111110_11011100 : OUT <= 0;  //62 / 220 = 0
    16'b00111110_11011101 : OUT <= 0;  //62 / 221 = 0
    16'b00111110_11011110 : OUT <= 0;  //62 / 222 = 0
    16'b00111110_11011111 : OUT <= 0;  //62 / 223 = 0
    16'b00111110_11100000 : OUT <= 0;  //62 / 224 = 0
    16'b00111110_11100001 : OUT <= 0;  //62 / 225 = 0
    16'b00111110_11100010 : OUT <= 0;  //62 / 226 = 0
    16'b00111110_11100011 : OUT <= 0;  //62 / 227 = 0
    16'b00111110_11100100 : OUT <= 0;  //62 / 228 = 0
    16'b00111110_11100101 : OUT <= 0;  //62 / 229 = 0
    16'b00111110_11100110 : OUT <= 0;  //62 / 230 = 0
    16'b00111110_11100111 : OUT <= 0;  //62 / 231 = 0
    16'b00111110_11101000 : OUT <= 0;  //62 / 232 = 0
    16'b00111110_11101001 : OUT <= 0;  //62 / 233 = 0
    16'b00111110_11101010 : OUT <= 0;  //62 / 234 = 0
    16'b00111110_11101011 : OUT <= 0;  //62 / 235 = 0
    16'b00111110_11101100 : OUT <= 0;  //62 / 236 = 0
    16'b00111110_11101101 : OUT <= 0;  //62 / 237 = 0
    16'b00111110_11101110 : OUT <= 0;  //62 / 238 = 0
    16'b00111110_11101111 : OUT <= 0;  //62 / 239 = 0
    16'b00111110_11110000 : OUT <= 0;  //62 / 240 = 0
    16'b00111110_11110001 : OUT <= 0;  //62 / 241 = 0
    16'b00111110_11110010 : OUT <= 0;  //62 / 242 = 0
    16'b00111110_11110011 : OUT <= 0;  //62 / 243 = 0
    16'b00111110_11110100 : OUT <= 0;  //62 / 244 = 0
    16'b00111110_11110101 : OUT <= 0;  //62 / 245 = 0
    16'b00111110_11110110 : OUT <= 0;  //62 / 246 = 0
    16'b00111110_11110111 : OUT <= 0;  //62 / 247 = 0
    16'b00111110_11111000 : OUT <= 0;  //62 / 248 = 0
    16'b00111110_11111001 : OUT <= 0;  //62 / 249 = 0
    16'b00111110_11111010 : OUT <= 0;  //62 / 250 = 0
    16'b00111110_11111011 : OUT <= 0;  //62 / 251 = 0
    16'b00111110_11111100 : OUT <= 0;  //62 / 252 = 0
    16'b00111110_11111101 : OUT <= 0;  //62 / 253 = 0
    16'b00111110_11111110 : OUT <= 0;  //62 / 254 = 0
    16'b00111110_11111111 : OUT <= 0;  //62 / 255 = 0
    16'b00111111_00000000 : OUT <= 0;  //63 / 0 = 0
    16'b00111111_00000001 : OUT <= 63;  //63 / 1 = 63
    16'b00111111_00000010 : OUT <= 31;  //63 / 2 = 31
    16'b00111111_00000011 : OUT <= 21;  //63 / 3 = 21
    16'b00111111_00000100 : OUT <= 15;  //63 / 4 = 15
    16'b00111111_00000101 : OUT <= 12;  //63 / 5 = 12
    16'b00111111_00000110 : OUT <= 10;  //63 / 6 = 10
    16'b00111111_00000111 : OUT <= 9;  //63 / 7 = 9
    16'b00111111_00001000 : OUT <= 7;  //63 / 8 = 7
    16'b00111111_00001001 : OUT <= 7;  //63 / 9 = 7
    16'b00111111_00001010 : OUT <= 6;  //63 / 10 = 6
    16'b00111111_00001011 : OUT <= 5;  //63 / 11 = 5
    16'b00111111_00001100 : OUT <= 5;  //63 / 12 = 5
    16'b00111111_00001101 : OUT <= 4;  //63 / 13 = 4
    16'b00111111_00001110 : OUT <= 4;  //63 / 14 = 4
    16'b00111111_00001111 : OUT <= 4;  //63 / 15 = 4
    16'b00111111_00010000 : OUT <= 3;  //63 / 16 = 3
    16'b00111111_00010001 : OUT <= 3;  //63 / 17 = 3
    16'b00111111_00010010 : OUT <= 3;  //63 / 18 = 3
    16'b00111111_00010011 : OUT <= 3;  //63 / 19 = 3
    16'b00111111_00010100 : OUT <= 3;  //63 / 20 = 3
    16'b00111111_00010101 : OUT <= 3;  //63 / 21 = 3
    16'b00111111_00010110 : OUT <= 2;  //63 / 22 = 2
    16'b00111111_00010111 : OUT <= 2;  //63 / 23 = 2
    16'b00111111_00011000 : OUT <= 2;  //63 / 24 = 2
    16'b00111111_00011001 : OUT <= 2;  //63 / 25 = 2
    16'b00111111_00011010 : OUT <= 2;  //63 / 26 = 2
    16'b00111111_00011011 : OUT <= 2;  //63 / 27 = 2
    16'b00111111_00011100 : OUT <= 2;  //63 / 28 = 2
    16'b00111111_00011101 : OUT <= 2;  //63 / 29 = 2
    16'b00111111_00011110 : OUT <= 2;  //63 / 30 = 2
    16'b00111111_00011111 : OUT <= 2;  //63 / 31 = 2
    16'b00111111_00100000 : OUT <= 1;  //63 / 32 = 1
    16'b00111111_00100001 : OUT <= 1;  //63 / 33 = 1
    16'b00111111_00100010 : OUT <= 1;  //63 / 34 = 1
    16'b00111111_00100011 : OUT <= 1;  //63 / 35 = 1
    16'b00111111_00100100 : OUT <= 1;  //63 / 36 = 1
    16'b00111111_00100101 : OUT <= 1;  //63 / 37 = 1
    16'b00111111_00100110 : OUT <= 1;  //63 / 38 = 1
    16'b00111111_00100111 : OUT <= 1;  //63 / 39 = 1
    16'b00111111_00101000 : OUT <= 1;  //63 / 40 = 1
    16'b00111111_00101001 : OUT <= 1;  //63 / 41 = 1
    16'b00111111_00101010 : OUT <= 1;  //63 / 42 = 1
    16'b00111111_00101011 : OUT <= 1;  //63 / 43 = 1
    16'b00111111_00101100 : OUT <= 1;  //63 / 44 = 1
    16'b00111111_00101101 : OUT <= 1;  //63 / 45 = 1
    16'b00111111_00101110 : OUT <= 1;  //63 / 46 = 1
    16'b00111111_00101111 : OUT <= 1;  //63 / 47 = 1
    16'b00111111_00110000 : OUT <= 1;  //63 / 48 = 1
    16'b00111111_00110001 : OUT <= 1;  //63 / 49 = 1
    16'b00111111_00110010 : OUT <= 1;  //63 / 50 = 1
    16'b00111111_00110011 : OUT <= 1;  //63 / 51 = 1
    16'b00111111_00110100 : OUT <= 1;  //63 / 52 = 1
    16'b00111111_00110101 : OUT <= 1;  //63 / 53 = 1
    16'b00111111_00110110 : OUT <= 1;  //63 / 54 = 1
    16'b00111111_00110111 : OUT <= 1;  //63 / 55 = 1
    16'b00111111_00111000 : OUT <= 1;  //63 / 56 = 1
    16'b00111111_00111001 : OUT <= 1;  //63 / 57 = 1
    16'b00111111_00111010 : OUT <= 1;  //63 / 58 = 1
    16'b00111111_00111011 : OUT <= 1;  //63 / 59 = 1
    16'b00111111_00111100 : OUT <= 1;  //63 / 60 = 1
    16'b00111111_00111101 : OUT <= 1;  //63 / 61 = 1
    16'b00111111_00111110 : OUT <= 1;  //63 / 62 = 1
    16'b00111111_00111111 : OUT <= 1;  //63 / 63 = 1
    16'b00111111_01000000 : OUT <= 0;  //63 / 64 = 0
    16'b00111111_01000001 : OUT <= 0;  //63 / 65 = 0
    16'b00111111_01000010 : OUT <= 0;  //63 / 66 = 0
    16'b00111111_01000011 : OUT <= 0;  //63 / 67 = 0
    16'b00111111_01000100 : OUT <= 0;  //63 / 68 = 0
    16'b00111111_01000101 : OUT <= 0;  //63 / 69 = 0
    16'b00111111_01000110 : OUT <= 0;  //63 / 70 = 0
    16'b00111111_01000111 : OUT <= 0;  //63 / 71 = 0
    16'b00111111_01001000 : OUT <= 0;  //63 / 72 = 0
    16'b00111111_01001001 : OUT <= 0;  //63 / 73 = 0
    16'b00111111_01001010 : OUT <= 0;  //63 / 74 = 0
    16'b00111111_01001011 : OUT <= 0;  //63 / 75 = 0
    16'b00111111_01001100 : OUT <= 0;  //63 / 76 = 0
    16'b00111111_01001101 : OUT <= 0;  //63 / 77 = 0
    16'b00111111_01001110 : OUT <= 0;  //63 / 78 = 0
    16'b00111111_01001111 : OUT <= 0;  //63 / 79 = 0
    16'b00111111_01010000 : OUT <= 0;  //63 / 80 = 0
    16'b00111111_01010001 : OUT <= 0;  //63 / 81 = 0
    16'b00111111_01010010 : OUT <= 0;  //63 / 82 = 0
    16'b00111111_01010011 : OUT <= 0;  //63 / 83 = 0
    16'b00111111_01010100 : OUT <= 0;  //63 / 84 = 0
    16'b00111111_01010101 : OUT <= 0;  //63 / 85 = 0
    16'b00111111_01010110 : OUT <= 0;  //63 / 86 = 0
    16'b00111111_01010111 : OUT <= 0;  //63 / 87 = 0
    16'b00111111_01011000 : OUT <= 0;  //63 / 88 = 0
    16'b00111111_01011001 : OUT <= 0;  //63 / 89 = 0
    16'b00111111_01011010 : OUT <= 0;  //63 / 90 = 0
    16'b00111111_01011011 : OUT <= 0;  //63 / 91 = 0
    16'b00111111_01011100 : OUT <= 0;  //63 / 92 = 0
    16'b00111111_01011101 : OUT <= 0;  //63 / 93 = 0
    16'b00111111_01011110 : OUT <= 0;  //63 / 94 = 0
    16'b00111111_01011111 : OUT <= 0;  //63 / 95 = 0
    16'b00111111_01100000 : OUT <= 0;  //63 / 96 = 0
    16'b00111111_01100001 : OUT <= 0;  //63 / 97 = 0
    16'b00111111_01100010 : OUT <= 0;  //63 / 98 = 0
    16'b00111111_01100011 : OUT <= 0;  //63 / 99 = 0
    16'b00111111_01100100 : OUT <= 0;  //63 / 100 = 0
    16'b00111111_01100101 : OUT <= 0;  //63 / 101 = 0
    16'b00111111_01100110 : OUT <= 0;  //63 / 102 = 0
    16'b00111111_01100111 : OUT <= 0;  //63 / 103 = 0
    16'b00111111_01101000 : OUT <= 0;  //63 / 104 = 0
    16'b00111111_01101001 : OUT <= 0;  //63 / 105 = 0
    16'b00111111_01101010 : OUT <= 0;  //63 / 106 = 0
    16'b00111111_01101011 : OUT <= 0;  //63 / 107 = 0
    16'b00111111_01101100 : OUT <= 0;  //63 / 108 = 0
    16'b00111111_01101101 : OUT <= 0;  //63 / 109 = 0
    16'b00111111_01101110 : OUT <= 0;  //63 / 110 = 0
    16'b00111111_01101111 : OUT <= 0;  //63 / 111 = 0
    16'b00111111_01110000 : OUT <= 0;  //63 / 112 = 0
    16'b00111111_01110001 : OUT <= 0;  //63 / 113 = 0
    16'b00111111_01110010 : OUT <= 0;  //63 / 114 = 0
    16'b00111111_01110011 : OUT <= 0;  //63 / 115 = 0
    16'b00111111_01110100 : OUT <= 0;  //63 / 116 = 0
    16'b00111111_01110101 : OUT <= 0;  //63 / 117 = 0
    16'b00111111_01110110 : OUT <= 0;  //63 / 118 = 0
    16'b00111111_01110111 : OUT <= 0;  //63 / 119 = 0
    16'b00111111_01111000 : OUT <= 0;  //63 / 120 = 0
    16'b00111111_01111001 : OUT <= 0;  //63 / 121 = 0
    16'b00111111_01111010 : OUT <= 0;  //63 / 122 = 0
    16'b00111111_01111011 : OUT <= 0;  //63 / 123 = 0
    16'b00111111_01111100 : OUT <= 0;  //63 / 124 = 0
    16'b00111111_01111101 : OUT <= 0;  //63 / 125 = 0
    16'b00111111_01111110 : OUT <= 0;  //63 / 126 = 0
    16'b00111111_01111111 : OUT <= 0;  //63 / 127 = 0
    16'b00111111_10000000 : OUT <= 0;  //63 / 128 = 0
    16'b00111111_10000001 : OUT <= 0;  //63 / 129 = 0
    16'b00111111_10000010 : OUT <= 0;  //63 / 130 = 0
    16'b00111111_10000011 : OUT <= 0;  //63 / 131 = 0
    16'b00111111_10000100 : OUT <= 0;  //63 / 132 = 0
    16'b00111111_10000101 : OUT <= 0;  //63 / 133 = 0
    16'b00111111_10000110 : OUT <= 0;  //63 / 134 = 0
    16'b00111111_10000111 : OUT <= 0;  //63 / 135 = 0
    16'b00111111_10001000 : OUT <= 0;  //63 / 136 = 0
    16'b00111111_10001001 : OUT <= 0;  //63 / 137 = 0
    16'b00111111_10001010 : OUT <= 0;  //63 / 138 = 0
    16'b00111111_10001011 : OUT <= 0;  //63 / 139 = 0
    16'b00111111_10001100 : OUT <= 0;  //63 / 140 = 0
    16'b00111111_10001101 : OUT <= 0;  //63 / 141 = 0
    16'b00111111_10001110 : OUT <= 0;  //63 / 142 = 0
    16'b00111111_10001111 : OUT <= 0;  //63 / 143 = 0
    16'b00111111_10010000 : OUT <= 0;  //63 / 144 = 0
    16'b00111111_10010001 : OUT <= 0;  //63 / 145 = 0
    16'b00111111_10010010 : OUT <= 0;  //63 / 146 = 0
    16'b00111111_10010011 : OUT <= 0;  //63 / 147 = 0
    16'b00111111_10010100 : OUT <= 0;  //63 / 148 = 0
    16'b00111111_10010101 : OUT <= 0;  //63 / 149 = 0
    16'b00111111_10010110 : OUT <= 0;  //63 / 150 = 0
    16'b00111111_10010111 : OUT <= 0;  //63 / 151 = 0
    16'b00111111_10011000 : OUT <= 0;  //63 / 152 = 0
    16'b00111111_10011001 : OUT <= 0;  //63 / 153 = 0
    16'b00111111_10011010 : OUT <= 0;  //63 / 154 = 0
    16'b00111111_10011011 : OUT <= 0;  //63 / 155 = 0
    16'b00111111_10011100 : OUT <= 0;  //63 / 156 = 0
    16'b00111111_10011101 : OUT <= 0;  //63 / 157 = 0
    16'b00111111_10011110 : OUT <= 0;  //63 / 158 = 0
    16'b00111111_10011111 : OUT <= 0;  //63 / 159 = 0
    16'b00111111_10100000 : OUT <= 0;  //63 / 160 = 0
    16'b00111111_10100001 : OUT <= 0;  //63 / 161 = 0
    16'b00111111_10100010 : OUT <= 0;  //63 / 162 = 0
    16'b00111111_10100011 : OUT <= 0;  //63 / 163 = 0
    16'b00111111_10100100 : OUT <= 0;  //63 / 164 = 0
    16'b00111111_10100101 : OUT <= 0;  //63 / 165 = 0
    16'b00111111_10100110 : OUT <= 0;  //63 / 166 = 0
    16'b00111111_10100111 : OUT <= 0;  //63 / 167 = 0
    16'b00111111_10101000 : OUT <= 0;  //63 / 168 = 0
    16'b00111111_10101001 : OUT <= 0;  //63 / 169 = 0
    16'b00111111_10101010 : OUT <= 0;  //63 / 170 = 0
    16'b00111111_10101011 : OUT <= 0;  //63 / 171 = 0
    16'b00111111_10101100 : OUT <= 0;  //63 / 172 = 0
    16'b00111111_10101101 : OUT <= 0;  //63 / 173 = 0
    16'b00111111_10101110 : OUT <= 0;  //63 / 174 = 0
    16'b00111111_10101111 : OUT <= 0;  //63 / 175 = 0
    16'b00111111_10110000 : OUT <= 0;  //63 / 176 = 0
    16'b00111111_10110001 : OUT <= 0;  //63 / 177 = 0
    16'b00111111_10110010 : OUT <= 0;  //63 / 178 = 0
    16'b00111111_10110011 : OUT <= 0;  //63 / 179 = 0
    16'b00111111_10110100 : OUT <= 0;  //63 / 180 = 0
    16'b00111111_10110101 : OUT <= 0;  //63 / 181 = 0
    16'b00111111_10110110 : OUT <= 0;  //63 / 182 = 0
    16'b00111111_10110111 : OUT <= 0;  //63 / 183 = 0
    16'b00111111_10111000 : OUT <= 0;  //63 / 184 = 0
    16'b00111111_10111001 : OUT <= 0;  //63 / 185 = 0
    16'b00111111_10111010 : OUT <= 0;  //63 / 186 = 0
    16'b00111111_10111011 : OUT <= 0;  //63 / 187 = 0
    16'b00111111_10111100 : OUT <= 0;  //63 / 188 = 0
    16'b00111111_10111101 : OUT <= 0;  //63 / 189 = 0
    16'b00111111_10111110 : OUT <= 0;  //63 / 190 = 0
    16'b00111111_10111111 : OUT <= 0;  //63 / 191 = 0
    16'b00111111_11000000 : OUT <= 0;  //63 / 192 = 0
    16'b00111111_11000001 : OUT <= 0;  //63 / 193 = 0
    16'b00111111_11000010 : OUT <= 0;  //63 / 194 = 0
    16'b00111111_11000011 : OUT <= 0;  //63 / 195 = 0
    16'b00111111_11000100 : OUT <= 0;  //63 / 196 = 0
    16'b00111111_11000101 : OUT <= 0;  //63 / 197 = 0
    16'b00111111_11000110 : OUT <= 0;  //63 / 198 = 0
    16'b00111111_11000111 : OUT <= 0;  //63 / 199 = 0
    16'b00111111_11001000 : OUT <= 0;  //63 / 200 = 0
    16'b00111111_11001001 : OUT <= 0;  //63 / 201 = 0
    16'b00111111_11001010 : OUT <= 0;  //63 / 202 = 0
    16'b00111111_11001011 : OUT <= 0;  //63 / 203 = 0
    16'b00111111_11001100 : OUT <= 0;  //63 / 204 = 0
    16'b00111111_11001101 : OUT <= 0;  //63 / 205 = 0
    16'b00111111_11001110 : OUT <= 0;  //63 / 206 = 0
    16'b00111111_11001111 : OUT <= 0;  //63 / 207 = 0
    16'b00111111_11010000 : OUT <= 0;  //63 / 208 = 0
    16'b00111111_11010001 : OUT <= 0;  //63 / 209 = 0
    16'b00111111_11010010 : OUT <= 0;  //63 / 210 = 0
    16'b00111111_11010011 : OUT <= 0;  //63 / 211 = 0
    16'b00111111_11010100 : OUT <= 0;  //63 / 212 = 0
    16'b00111111_11010101 : OUT <= 0;  //63 / 213 = 0
    16'b00111111_11010110 : OUT <= 0;  //63 / 214 = 0
    16'b00111111_11010111 : OUT <= 0;  //63 / 215 = 0
    16'b00111111_11011000 : OUT <= 0;  //63 / 216 = 0
    16'b00111111_11011001 : OUT <= 0;  //63 / 217 = 0
    16'b00111111_11011010 : OUT <= 0;  //63 / 218 = 0
    16'b00111111_11011011 : OUT <= 0;  //63 / 219 = 0
    16'b00111111_11011100 : OUT <= 0;  //63 / 220 = 0
    16'b00111111_11011101 : OUT <= 0;  //63 / 221 = 0
    16'b00111111_11011110 : OUT <= 0;  //63 / 222 = 0
    16'b00111111_11011111 : OUT <= 0;  //63 / 223 = 0
    16'b00111111_11100000 : OUT <= 0;  //63 / 224 = 0
    16'b00111111_11100001 : OUT <= 0;  //63 / 225 = 0
    16'b00111111_11100010 : OUT <= 0;  //63 / 226 = 0
    16'b00111111_11100011 : OUT <= 0;  //63 / 227 = 0
    16'b00111111_11100100 : OUT <= 0;  //63 / 228 = 0
    16'b00111111_11100101 : OUT <= 0;  //63 / 229 = 0
    16'b00111111_11100110 : OUT <= 0;  //63 / 230 = 0
    16'b00111111_11100111 : OUT <= 0;  //63 / 231 = 0
    16'b00111111_11101000 : OUT <= 0;  //63 / 232 = 0
    16'b00111111_11101001 : OUT <= 0;  //63 / 233 = 0
    16'b00111111_11101010 : OUT <= 0;  //63 / 234 = 0
    16'b00111111_11101011 : OUT <= 0;  //63 / 235 = 0
    16'b00111111_11101100 : OUT <= 0;  //63 / 236 = 0
    16'b00111111_11101101 : OUT <= 0;  //63 / 237 = 0
    16'b00111111_11101110 : OUT <= 0;  //63 / 238 = 0
    16'b00111111_11101111 : OUT <= 0;  //63 / 239 = 0
    16'b00111111_11110000 : OUT <= 0;  //63 / 240 = 0
    16'b00111111_11110001 : OUT <= 0;  //63 / 241 = 0
    16'b00111111_11110010 : OUT <= 0;  //63 / 242 = 0
    16'b00111111_11110011 : OUT <= 0;  //63 / 243 = 0
    16'b00111111_11110100 : OUT <= 0;  //63 / 244 = 0
    16'b00111111_11110101 : OUT <= 0;  //63 / 245 = 0
    16'b00111111_11110110 : OUT <= 0;  //63 / 246 = 0
    16'b00111111_11110111 : OUT <= 0;  //63 / 247 = 0
    16'b00111111_11111000 : OUT <= 0;  //63 / 248 = 0
    16'b00111111_11111001 : OUT <= 0;  //63 / 249 = 0
    16'b00111111_11111010 : OUT <= 0;  //63 / 250 = 0
    16'b00111111_11111011 : OUT <= 0;  //63 / 251 = 0
    16'b00111111_11111100 : OUT <= 0;  //63 / 252 = 0
    16'b00111111_11111101 : OUT <= 0;  //63 / 253 = 0
    16'b00111111_11111110 : OUT <= 0;  //63 / 254 = 0
    16'b00111111_11111111 : OUT <= 0;  //63 / 255 = 0
    16'b01000000_00000000 : OUT <= 0;  //64 / 0 = 0
    16'b01000000_00000001 : OUT <= 64;  //64 / 1 = 64
    16'b01000000_00000010 : OUT <= 32;  //64 / 2 = 32
    16'b01000000_00000011 : OUT <= 21;  //64 / 3 = 21
    16'b01000000_00000100 : OUT <= 16;  //64 / 4 = 16
    16'b01000000_00000101 : OUT <= 12;  //64 / 5 = 12
    16'b01000000_00000110 : OUT <= 10;  //64 / 6 = 10
    16'b01000000_00000111 : OUT <= 9;  //64 / 7 = 9
    16'b01000000_00001000 : OUT <= 8;  //64 / 8 = 8
    16'b01000000_00001001 : OUT <= 7;  //64 / 9 = 7
    16'b01000000_00001010 : OUT <= 6;  //64 / 10 = 6
    16'b01000000_00001011 : OUT <= 5;  //64 / 11 = 5
    16'b01000000_00001100 : OUT <= 5;  //64 / 12 = 5
    16'b01000000_00001101 : OUT <= 4;  //64 / 13 = 4
    16'b01000000_00001110 : OUT <= 4;  //64 / 14 = 4
    16'b01000000_00001111 : OUT <= 4;  //64 / 15 = 4
    16'b01000000_00010000 : OUT <= 4;  //64 / 16 = 4
    16'b01000000_00010001 : OUT <= 3;  //64 / 17 = 3
    16'b01000000_00010010 : OUT <= 3;  //64 / 18 = 3
    16'b01000000_00010011 : OUT <= 3;  //64 / 19 = 3
    16'b01000000_00010100 : OUT <= 3;  //64 / 20 = 3
    16'b01000000_00010101 : OUT <= 3;  //64 / 21 = 3
    16'b01000000_00010110 : OUT <= 2;  //64 / 22 = 2
    16'b01000000_00010111 : OUT <= 2;  //64 / 23 = 2
    16'b01000000_00011000 : OUT <= 2;  //64 / 24 = 2
    16'b01000000_00011001 : OUT <= 2;  //64 / 25 = 2
    16'b01000000_00011010 : OUT <= 2;  //64 / 26 = 2
    16'b01000000_00011011 : OUT <= 2;  //64 / 27 = 2
    16'b01000000_00011100 : OUT <= 2;  //64 / 28 = 2
    16'b01000000_00011101 : OUT <= 2;  //64 / 29 = 2
    16'b01000000_00011110 : OUT <= 2;  //64 / 30 = 2
    16'b01000000_00011111 : OUT <= 2;  //64 / 31 = 2
    16'b01000000_00100000 : OUT <= 2;  //64 / 32 = 2
    16'b01000000_00100001 : OUT <= 1;  //64 / 33 = 1
    16'b01000000_00100010 : OUT <= 1;  //64 / 34 = 1
    16'b01000000_00100011 : OUT <= 1;  //64 / 35 = 1
    16'b01000000_00100100 : OUT <= 1;  //64 / 36 = 1
    16'b01000000_00100101 : OUT <= 1;  //64 / 37 = 1
    16'b01000000_00100110 : OUT <= 1;  //64 / 38 = 1
    16'b01000000_00100111 : OUT <= 1;  //64 / 39 = 1
    16'b01000000_00101000 : OUT <= 1;  //64 / 40 = 1
    16'b01000000_00101001 : OUT <= 1;  //64 / 41 = 1
    16'b01000000_00101010 : OUT <= 1;  //64 / 42 = 1
    16'b01000000_00101011 : OUT <= 1;  //64 / 43 = 1
    16'b01000000_00101100 : OUT <= 1;  //64 / 44 = 1
    16'b01000000_00101101 : OUT <= 1;  //64 / 45 = 1
    16'b01000000_00101110 : OUT <= 1;  //64 / 46 = 1
    16'b01000000_00101111 : OUT <= 1;  //64 / 47 = 1
    16'b01000000_00110000 : OUT <= 1;  //64 / 48 = 1
    16'b01000000_00110001 : OUT <= 1;  //64 / 49 = 1
    16'b01000000_00110010 : OUT <= 1;  //64 / 50 = 1
    16'b01000000_00110011 : OUT <= 1;  //64 / 51 = 1
    16'b01000000_00110100 : OUT <= 1;  //64 / 52 = 1
    16'b01000000_00110101 : OUT <= 1;  //64 / 53 = 1
    16'b01000000_00110110 : OUT <= 1;  //64 / 54 = 1
    16'b01000000_00110111 : OUT <= 1;  //64 / 55 = 1
    16'b01000000_00111000 : OUT <= 1;  //64 / 56 = 1
    16'b01000000_00111001 : OUT <= 1;  //64 / 57 = 1
    16'b01000000_00111010 : OUT <= 1;  //64 / 58 = 1
    16'b01000000_00111011 : OUT <= 1;  //64 / 59 = 1
    16'b01000000_00111100 : OUT <= 1;  //64 / 60 = 1
    16'b01000000_00111101 : OUT <= 1;  //64 / 61 = 1
    16'b01000000_00111110 : OUT <= 1;  //64 / 62 = 1
    16'b01000000_00111111 : OUT <= 1;  //64 / 63 = 1
    16'b01000000_01000000 : OUT <= 1;  //64 / 64 = 1
    16'b01000000_01000001 : OUT <= 0;  //64 / 65 = 0
    16'b01000000_01000010 : OUT <= 0;  //64 / 66 = 0
    16'b01000000_01000011 : OUT <= 0;  //64 / 67 = 0
    16'b01000000_01000100 : OUT <= 0;  //64 / 68 = 0
    16'b01000000_01000101 : OUT <= 0;  //64 / 69 = 0
    16'b01000000_01000110 : OUT <= 0;  //64 / 70 = 0
    16'b01000000_01000111 : OUT <= 0;  //64 / 71 = 0
    16'b01000000_01001000 : OUT <= 0;  //64 / 72 = 0
    16'b01000000_01001001 : OUT <= 0;  //64 / 73 = 0
    16'b01000000_01001010 : OUT <= 0;  //64 / 74 = 0
    16'b01000000_01001011 : OUT <= 0;  //64 / 75 = 0
    16'b01000000_01001100 : OUT <= 0;  //64 / 76 = 0
    16'b01000000_01001101 : OUT <= 0;  //64 / 77 = 0
    16'b01000000_01001110 : OUT <= 0;  //64 / 78 = 0
    16'b01000000_01001111 : OUT <= 0;  //64 / 79 = 0
    16'b01000000_01010000 : OUT <= 0;  //64 / 80 = 0
    16'b01000000_01010001 : OUT <= 0;  //64 / 81 = 0
    16'b01000000_01010010 : OUT <= 0;  //64 / 82 = 0
    16'b01000000_01010011 : OUT <= 0;  //64 / 83 = 0
    16'b01000000_01010100 : OUT <= 0;  //64 / 84 = 0
    16'b01000000_01010101 : OUT <= 0;  //64 / 85 = 0
    16'b01000000_01010110 : OUT <= 0;  //64 / 86 = 0
    16'b01000000_01010111 : OUT <= 0;  //64 / 87 = 0
    16'b01000000_01011000 : OUT <= 0;  //64 / 88 = 0
    16'b01000000_01011001 : OUT <= 0;  //64 / 89 = 0
    16'b01000000_01011010 : OUT <= 0;  //64 / 90 = 0
    16'b01000000_01011011 : OUT <= 0;  //64 / 91 = 0
    16'b01000000_01011100 : OUT <= 0;  //64 / 92 = 0
    16'b01000000_01011101 : OUT <= 0;  //64 / 93 = 0
    16'b01000000_01011110 : OUT <= 0;  //64 / 94 = 0
    16'b01000000_01011111 : OUT <= 0;  //64 / 95 = 0
    16'b01000000_01100000 : OUT <= 0;  //64 / 96 = 0
    16'b01000000_01100001 : OUT <= 0;  //64 / 97 = 0
    16'b01000000_01100010 : OUT <= 0;  //64 / 98 = 0
    16'b01000000_01100011 : OUT <= 0;  //64 / 99 = 0
    16'b01000000_01100100 : OUT <= 0;  //64 / 100 = 0
    16'b01000000_01100101 : OUT <= 0;  //64 / 101 = 0
    16'b01000000_01100110 : OUT <= 0;  //64 / 102 = 0
    16'b01000000_01100111 : OUT <= 0;  //64 / 103 = 0
    16'b01000000_01101000 : OUT <= 0;  //64 / 104 = 0
    16'b01000000_01101001 : OUT <= 0;  //64 / 105 = 0
    16'b01000000_01101010 : OUT <= 0;  //64 / 106 = 0
    16'b01000000_01101011 : OUT <= 0;  //64 / 107 = 0
    16'b01000000_01101100 : OUT <= 0;  //64 / 108 = 0
    16'b01000000_01101101 : OUT <= 0;  //64 / 109 = 0
    16'b01000000_01101110 : OUT <= 0;  //64 / 110 = 0
    16'b01000000_01101111 : OUT <= 0;  //64 / 111 = 0
    16'b01000000_01110000 : OUT <= 0;  //64 / 112 = 0
    16'b01000000_01110001 : OUT <= 0;  //64 / 113 = 0
    16'b01000000_01110010 : OUT <= 0;  //64 / 114 = 0
    16'b01000000_01110011 : OUT <= 0;  //64 / 115 = 0
    16'b01000000_01110100 : OUT <= 0;  //64 / 116 = 0
    16'b01000000_01110101 : OUT <= 0;  //64 / 117 = 0
    16'b01000000_01110110 : OUT <= 0;  //64 / 118 = 0
    16'b01000000_01110111 : OUT <= 0;  //64 / 119 = 0
    16'b01000000_01111000 : OUT <= 0;  //64 / 120 = 0
    16'b01000000_01111001 : OUT <= 0;  //64 / 121 = 0
    16'b01000000_01111010 : OUT <= 0;  //64 / 122 = 0
    16'b01000000_01111011 : OUT <= 0;  //64 / 123 = 0
    16'b01000000_01111100 : OUT <= 0;  //64 / 124 = 0
    16'b01000000_01111101 : OUT <= 0;  //64 / 125 = 0
    16'b01000000_01111110 : OUT <= 0;  //64 / 126 = 0
    16'b01000000_01111111 : OUT <= 0;  //64 / 127 = 0
    16'b01000000_10000000 : OUT <= 0;  //64 / 128 = 0
    16'b01000000_10000001 : OUT <= 0;  //64 / 129 = 0
    16'b01000000_10000010 : OUT <= 0;  //64 / 130 = 0
    16'b01000000_10000011 : OUT <= 0;  //64 / 131 = 0
    16'b01000000_10000100 : OUT <= 0;  //64 / 132 = 0
    16'b01000000_10000101 : OUT <= 0;  //64 / 133 = 0
    16'b01000000_10000110 : OUT <= 0;  //64 / 134 = 0
    16'b01000000_10000111 : OUT <= 0;  //64 / 135 = 0
    16'b01000000_10001000 : OUT <= 0;  //64 / 136 = 0
    16'b01000000_10001001 : OUT <= 0;  //64 / 137 = 0
    16'b01000000_10001010 : OUT <= 0;  //64 / 138 = 0
    16'b01000000_10001011 : OUT <= 0;  //64 / 139 = 0
    16'b01000000_10001100 : OUT <= 0;  //64 / 140 = 0
    16'b01000000_10001101 : OUT <= 0;  //64 / 141 = 0
    16'b01000000_10001110 : OUT <= 0;  //64 / 142 = 0
    16'b01000000_10001111 : OUT <= 0;  //64 / 143 = 0
    16'b01000000_10010000 : OUT <= 0;  //64 / 144 = 0
    16'b01000000_10010001 : OUT <= 0;  //64 / 145 = 0
    16'b01000000_10010010 : OUT <= 0;  //64 / 146 = 0
    16'b01000000_10010011 : OUT <= 0;  //64 / 147 = 0
    16'b01000000_10010100 : OUT <= 0;  //64 / 148 = 0
    16'b01000000_10010101 : OUT <= 0;  //64 / 149 = 0
    16'b01000000_10010110 : OUT <= 0;  //64 / 150 = 0
    16'b01000000_10010111 : OUT <= 0;  //64 / 151 = 0
    16'b01000000_10011000 : OUT <= 0;  //64 / 152 = 0
    16'b01000000_10011001 : OUT <= 0;  //64 / 153 = 0
    16'b01000000_10011010 : OUT <= 0;  //64 / 154 = 0
    16'b01000000_10011011 : OUT <= 0;  //64 / 155 = 0
    16'b01000000_10011100 : OUT <= 0;  //64 / 156 = 0
    16'b01000000_10011101 : OUT <= 0;  //64 / 157 = 0
    16'b01000000_10011110 : OUT <= 0;  //64 / 158 = 0
    16'b01000000_10011111 : OUT <= 0;  //64 / 159 = 0
    16'b01000000_10100000 : OUT <= 0;  //64 / 160 = 0
    16'b01000000_10100001 : OUT <= 0;  //64 / 161 = 0
    16'b01000000_10100010 : OUT <= 0;  //64 / 162 = 0
    16'b01000000_10100011 : OUT <= 0;  //64 / 163 = 0
    16'b01000000_10100100 : OUT <= 0;  //64 / 164 = 0
    16'b01000000_10100101 : OUT <= 0;  //64 / 165 = 0
    16'b01000000_10100110 : OUT <= 0;  //64 / 166 = 0
    16'b01000000_10100111 : OUT <= 0;  //64 / 167 = 0
    16'b01000000_10101000 : OUT <= 0;  //64 / 168 = 0
    16'b01000000_10101001 : OUT <= 0;  //64 / 169 = 0
    16'b01000000_10101010 : OUT <= 0;  //64 / 170 = 0
    16'b01000000_10101011 : OUT <= 0;  //64 / 171 = 0
    16'b01000000_10101100 : OUT <= 0;  //64 / 172 = 0
    16'b01000000_10101101 : OUT <= 0;  //64 / 173 = 0
    16'b01000000_10101110 : OUT <= 0;  //64 / 174 = 0
    16'b01000000_10101111 : OUT <= 0;  //64 / 175 = 0
    16'b01000000_10110000 : OUT <= 0;  //64 / 176 = 0
    16'b01000000_10110001 : OUT <= 0;  //64 / 177 = 0
    16'b01000000_10110010 : OUT <= 0;  //64 / 178 = 0
    16'b01000000_10110011 : OUT <= 0;  //64 / 179 = 0
    16'b01000000_10110100 : OUT <= 0;  //64 / 180 = 0
    16'b01000000_10110101 : OUT <= 0;  //64 / 181 = 0
    16'b01000000_10110110 : OUT <= 0;  //64 / 182 = 0
    16'b01000000_10110111 : OUT <= 0;  //64 / 183 = 0
    16'b01000000_10111000 : OUT <= 0;  //64 / 184 = 0
    16'b01000000_10111001 : OUT <= 0;  //64 / 185 = 0
    16'b01000000_10111010 : OUT <= 0;  //64 / 186 = 0
    16'b01000000_10111011 : OUT <= 0;  //64 / 187 = 0
    16'b01000000_10111100 : OUT <= 0;  //64 / 188 = 0
    16'b01000000_10111101 : OUT <= 0;  //64 / 189 = 0
    16'b01000000_10111110 : OUT <= 0;  //64 / 190 = 0
    16'b01000000_10111111 : OUT <= 0;  //64 / 191 = 0
    16'b01000000_11000000 : OUT <= 0;  //64 / 192 = 0
    16'b01000000_11000001 : OUT <= 0;  //64 / 193 = 0
    16'b01000000_11000010 : OUT <= 0;  //64 / 194 = 0
    16'b01000000_11000011 : OUT <= 0;  //64 / 195 = 0
    16'b01000000_11000100 : OUT <= 0;  //64 / 196 = 0
    16'b01000000_11000101 : OUT <= 0;  //64 / 197 = 0
    16'b01000000_11000110 : OUT <= 0;  //64 / 198 = 0
    16'b01000000_11000111 : OUT <= 0;  //64 / 199 = 0
    16'b01000000_11001000 : OUT <= 0;  //64 / 200 = 0
    16'b01000000_11001001 : OUT <= 0;  //64 / 201 = 0
    16'b01000000_11001010 : OUT <= 0;  //64 / 202 = 0
    16'b01000000_11001011 : OUT <= 0;  //64 / 203 = 0
    16'b01000000_11001100 : OUT <= 0;  //64 / 204 = 0
    16'b01000000_11001101 : OUT <= 0;  //64 / 205 = 0
    16'b01000000_11001110 : OUT <= 0;  //64 / 206 = 0
    16'b01000000_11001111 : OUT <= 0;  //64 / 207 = 0
    16'b01000000_11010000 : OUT <= 0;  //64 / 208 = 0
    16'b01000000_11010001 : OUT <= 0;  //64 / 209 = 0
    16'b01000000_11010010 : OUT <= 0;  //64 / 210 = 0
    16'b01000000_11010011 : OUT <= 0;  //64 / 211 = 0
    16'b01000000_11010100 : OUT <= 0;  //64 / 212 = 0
    16'b01000000_11010101 : OUT <= 0;  //64 / 213 = 0
    16'b01000000_11010110 : OUT <= 0;  //64 / 214 = 0
    16'b01000000_11010111 : OUT <= 0;  //64 / 215 = 0
    16'b01000000_11011000 : OUT <= 0;  //64 / 216 = 0
    16'b01000000_11011001 : OUT <= 0;  //64 / 217 = 0
    16'b01000000_11011010 : OUT <= 0;  //64 / 218 = 0
    16'b01000000_11011011 : OUT <= 0;  //64 / 219 = 0
    16'b01000000_11011100 : OUT <= 0;  //64 / 220 = 0
    16'b01000000_11011101 : OUT <= 0;  //64 / 221 = 0
    16'b01000000_11011110 : OUT <= 0;  //64 / 222 = 0
    16'b01000000_11011111 : OUT <= 0;  //64 / 223 = 0
    16'b01000000_11100000 : OUT <= 0;  //64 / 224 = 0
    16'b01000000_11100001 : OUT <= 0;  //64 / 225 = 0
    16'b01000000_11100010 : OUT <= 0;  //64 / 226 = 0
    16'b01000000_11100011 : OUT <= 0;  //64 / 227 = 0
    16'b01000000_11100100 : OUT <= 0;  //64 / 228 = 0
    16'b01000000_11100101 : OUT <= 0;  //64 / 229 = 0
    16'b01000000_11100110 : OUT <= 0;  //64 / 230 = 0
    16'b01000000_11100111 : OUT <= 0;  //64 / 231 = 0
    16'b01000000_11101000 : OUT <= 0;  //64 / 232 = 0
    16'b01000000_11101001 : OUT <= 0;  //64 / 233 = 0
    16'b01000000_11101010 : OUT <= 0;  //64 / 234 = 0
    16'b01000000_11101011 : OUT <= 0;  //64 / 235 = 0
    16'b01000000_11101100 : OUT <= 0;  //64 / 236 = 0
    16'b01000000_11101101 : OUT <= 0;  //64 / 237 = 0
    16'b01000000_11101110 : OUT <= 0;  //64 / 238 = 0
    16'b01000000_11101111 : OUT <= 0;  //64 / 239 = 0
    16'b01000000_11110000 : OUT <= 0;  //64 / 240 = 0
    16'b01000000_11110001 : OUT <= 0;  //64 / 241 = 0
    16'b01000000_11110010 : OUT <= 0;  //64 / 242 = 0
    16'b01000000_11110011 : OUT <= 0;  //64 / 243 = 0
    16'b01000000_11110100 : OUT <= 0;  //64 / 244 = 0
    16'b01000000_11110101 : OUT <= 0;  //64 / 245 = 0
    16'b01000000_11110110 : OUT <= 0;  //64 / 246 = 0
    16'b01000000_11110111 : OUT <= 0;  //64 / 247 = 0
    16'b01000000_11111000 : OUT <= 0;  //64 / 248 = 0
    16'b01000000_11111001 : OUT <= 0;  //64 / 249 = 0
    16'b01000000_11111010 : OUT <= 0;  //64 / 250 = 0
    16'b01000000_11111011 : OUT <= 0;  //64 / 251 = 0
    16'b01000000_11111100 : OUT <= 0;  //64 / 252 = 0
    16'b01000000_11111101 : OUT <= 0;  //64 / 253 = 0
    16'b01000000_11111110 : OUT <= 0;  //64 / 254 = 0
    16'b01000000_11111111 : OUT <= 0;  //64 / 255 = 0
    16'b01000001_00000000 : OUT <= 0;  //65 / 0 = 0
    16'b01000001_00000001 : OUT <= 65;  //65 / 1 = 65
    16'b01000001_00000010 : OUT <= 32;  //65 / 2 = 32
    16'b01000001_00000011 : OUT <= 21;  //65 / 3 = 21
    16'b01000001_00000100 : OUT <= 16;  //65 / 4 = 16
    16'b01000001_00000101 : OUT <= 13;  //65 / 5 = 13
    16'b01000001_00000110 : OUT <= 10;  //65 / 6 = 10
    16'b01000001_00000111 : OUT <= 9;  //65 / 7 = 9
    16'b01000001_00001000 : OUT <= 8;  //65 / 8 = 8
    16'b01000001_00001001 : OUT <= 7;  //65 / 9 = 7
    16'b01000001_00001010 : OUT <= 6;  //65 / 10 = 6
    16'b01000001_00001011 : OUT <= 5;  //65 / 11 = 5
    16'b01000001_00001100 : OUT <= 5;  //65 / 12 = 5
    16'b01000001_00001101 : OUT <= 5;  //65 / 13 = 5
    16'b01000001_00001110 : OUT <= 4;  //65 / 14 = 4
    16'b01000001_00001111 : OUT <= 4;  //65 / 15 = 4
    16'b01000001_00010000 : OUT <= 4;  //65 / 16 = 4
    16'b01000001_00010001 : OUT <= 3;  //65 / 17 = 3
    16'b01000001_00010010 : OUT <= 3;  //65 / 18 = 3
    16'b01000001_00010011 : OUT <= 3;  //65 / 19 = 3
    16'b01000001_00010100 : OUT <= 3;  //65 / 20 = 3
    16'b01000001_00010101 : OUT <= 3;  //65 / 21 = 3
    16'b01000001_00010110 : OUT <= 2;  //65 / 22 = 2
    16'b01000001_00010111 : OUT <= 2;  //65 / 23 = 2
    16'b01000001_00011000 : OUT <= 2;  //65 / 24 = 2
    16'b01000001_00011001 : OUT <= 2;  //65 / 25 = 2
    16'b01000001_00011010 : OUT <= 2;  //65 / 26 = 2
    16'b01000001_00011011 : OUT <= 2;  //65 / 27 = 2
    16'b01000001_00011100 : OUT <= 2;  //65 / 28 = 2
    16'b01000001_00011101 : OUT <= 2;  //65 / 29 = 2
    16'b01000001_00011110 : OUT <= 2;  //65 / 30 = 2
    16'b01000001_00011111 : OUT <= 2;  //65 / 31 = 2
    16'b01000001_00100000 : OUT <= 2;  //65 / 32 = 2
    16'b01000001_00100001 : OUT <= 1;  //65 / 33 = 1
    16'b01000001_00100010 : OUT <= 1;  //65 / 34 = 1
    16'b01000001_00100011 : OUT <= 1;  //65 / 35 = 1
    16'b01000001_00100100 : OUT <= 1;  //65 / 36 = 1
    16'b01000001_00100101 : OUT <= 1;  //65 / 37 = 1
    16'b01000001_00100110 : OUT <= 1;  //65 / 38 = 1
    16'b01000001_00100111 : OUT <= 1;  //65 / 39 = 1
    16'b01000001_00101000 : OUT <= 1;  //65 / 40 = 1
    16'b01000001_00101001 : OUT <= 1;  //65 / 41 = 1
    16'b01000001_00101010 : OUT <= 1;  //65 / 42 = 1
    16'b01000001_00101011 : OUT <= 1;  //65 / 43 = 1
    16'b01000001_00101100 : OUT <= 1;  //65 / 44 = 1
    16'b01000001_00101101 : OUT <= 1;  //65 / 45 = 1
    16'b01000001_00101110 : OUT <= 1;  //65 / 46 = 1
    16'b01000001_00101111 : OUT <= 1;  //65 / 47 = 1
    16'b01000001_00110000 : OUT <= 1;  //65 / 48 = 1
    16'b01000001_00110001 : OUT <= 1;  //65 / 49 = 1
    16'b01000001_00110010 : OUT <= 1;  //65 / 50 = 1
    16'b01000001_00110011 : OUT <= 1;  //65 / 51 = 1
    16'b01000001_00110100 : OUT <= 1;  //65 / 52 = 1
    16'b01000001_00110101 : OUT <= 1;  //65 / 53 = 1
    16'b01000001_00110110 : OUT <= 1;  //65 / 54 = 1
    16'b01000001_00110111 : OUT <= 1;  //65 / 55 = 1
    16'b01000001_00111000 : OUT <= 1;  //65 / 56 = 1
    16'b01000001_00111001 : OUT <= 1;  //65 / 57 = 1
    16'b01000001_00111010 : OUT <= 1;  //65 / 58 = 1
    16'b01000001_00111011 : OUT <= 1;  //65 / 59 = 1
    16'b01000001_00111100 : OUT <= 1;  //65 / 60 = 1
    16'b01000001_00111101 : OUT <= 1;  //65 / 61 = 1
    16'b01000001_00111110 : OUT <= 1;  //65 / 62 = 1
    16'b01000001_00111111 : OUT <= 1;  //65 / 63 = 1
    16'b01000001_01000000 : OUT <= 1;  //65 / 64 = 1
    16'b01000001_01000001 : OUT <= 1;  //65 / 65 = 1
    16'b01000001_01000010 : OUT <= 0;  //65 / 66 = 0
    16'b01000001_01000011 : OUT <= 0;  //65 / 67 = 0
    16'b01000001_01000100 : OUT <= 0;  //65 / 68 = 0
    16'b01000001_01000101 : OUT <= 0;  //65 / 69 = 0
    16'b01000001_01000110 : OUT <= 0;  //65 / 70 = 0
    16'b01000001_01000111 : OUT <= 0;  //65 / 71 = 0
    16'b01000001_01001000 : OUT <= 0;  //65 / 72 = 0
    16'b01000001_01001001 : OUT <= 0;  //65 / 73 = 0
    16'b01000001_01001010 : OUT <= 0;  //65 / 74 = 0
    16'b01000001_01001011 : OUT <= 0;  //65 / 75 = 0
    16'b01000001_01001100 : OUT <= 0;  //65 / 76 = 0
    16'b01000001_01001101 : OUT <= 0;  //65 / 77 = 0
    16'b01000001_01001110 : OUT <= 0;  //65 / 78 = 0
    16'b01000001_01001111 : OUT <= 0;  //65 / 79 = 0
    16'b01000001_01010000 : OUT <= 0;  //65 / 80 = 0
    16'b01000001_01010001 : OUT <= 0;  //65 / 81 = 0
    16'b01000001_01010010 : OUT <= 0;  //65 / 82 = 0
    16'b01000001_01010011 : OUT <= 0;  //65 / 83 = 0
    16'b01000001_01010100 : OUT <= 0;  //65 / 84 = 0
    16'b01000001_01010101 : OUT <= 0;  //65 / 85 = 0
    16'b01000001_01010110 : OUT <= 0;  //65 / 86 = 0
    16'b01000001_01010111 : OUT <= 0;  //65 / 87 = 0
    16'b01000001_01011000 : OUT <= 0;  //65 / 88 = 0
    16'b01000001_01011001 : OUT <= 0;  //65 / 89 = 0
    16'b01000001_01011010 : OUT <= 0;  //65 / 90 = 0
    16'b01000001_01011011 : OUT <= 0;  //65 / 91 = 0
    16'b01000001_01011100 : OUT <= 0;  //65 / 92 = 0
    16'b01000001_01011101 : OUT <= 0;  //65 / 93 = 0
    16'b01000001_01011110 : OUT <= 0;  //65 / 94 = 0
    16'b01000001_01011111 : OUT <= 0;  //65 / 95 = 0
    16'b01000001_01100000 : OUT <= 0;  //65 / 96 = 0
    16'b01000001_01100001 : OUT <= 0;  //65 / 97 = 0
    16'b01000001_01100010 : OUT <= 0;  //65 / 98 = 0
    16'b01000001_01100011 : OUT <= 0;  //65 / 99 = 0
    16'b01000001_01100100 : OUT <= 0;  //65 / 100 = 0
    16'b01000001_01100101 : OUT <= 0;  //65 / 101 = 0
    16'b01000001_01100110 : OUT <= 0;  //65 / 102 = 0
    16'b01000001_01100111 : OUT <= 0;  //65 / 103 = 0
    16'b01000001_01101000 : OUT <= 0;  //65 / 104 = 0
    16'b01000001_01101001 : OUT <= 0;  //65 / 105 = 0
    16'b01000001_01101010 : OUT <= 0;  //65 / 106 = 0
    16'b01000001_01101011 : OUT <= 0;  //65 / 107 = 0
    16'b01000001_01101100 : OUT <= 0;  //65 / 108 = 0
    16'b01000001_01101101 : OUT <= 0;  //65 / 109 = 0
    16'b01000001_01101110 : OUT <= 0;  //65 / 110 = 0
    16'b01000001_01101111 : OUT <= 0;  //65 / 111 = 0
    16'b01000001_01110000 : OUT <= 0;  //65 / 112 = 0
    16'b01000001_01110001 : OUT <= 0;  //65 / 113 = 0
    16'b01000001_01110010 : OUT <= 0;  //65 / 114 = 0
    16'b01000001_01110011 : OUT <= 0;  //65 / 115 = 0
    16'b01000001_01110100 : OUT <= 0;  //65 / 116 = 0
    16'b01000001_01110101 : OUT <= 0;  //65 / 117 = 0
    16'b01000001_01110110 : OUT <= 0;  //65 / 118 = 0
    16'b01000001_01110111 : OUT <= 0;  //65 / 119 = 0
    16'b01000001_01111000 : OUT <= 0;  //65 / 120 = 0
    16'b01000001_01111001 : OUT <= 0;  //65 / 121 = 0
    16'b01000001_01111010 : OUT <= 0;  //65 / 122 = 0
    16'b01000001_01111011 : OUT <= 0;  //65 / 123 = 0
    16'b01000001_01111100 : OUT <= 0;  //65 / 124 = 0
    16'b01000001_01111101 : OUT <= 0;  //65 / 125 = 0
    16'b01000001_01111110 : OUT <= 0;  //65 / 126 = 0
    16'b01000001_01111111 : OUT <= 0;  //65 / 127 = 0
    16'b01000001_10000000 : OUT <= 0;  //65 / 128 = 0
    16'b01000001_10000001 : OUT <= 0;  //65 / 129 = 0
    16'b01000001_10000010 : OUT <= 0;  //65 / 130 = 0
    16'b01000001_10000011 : OUT <= 0;  //65 / 131 = 0
    16'b01000001_10000100 : OUT <= 0;  //65 / 132 = 0
    16'b01000001_10000101 : OUT <= 0;  //65 / 133 = 0
    16'b01000001_10000110 : OUT <= 0;  //65 / 134 = 0
    16'b01000001_10000111 : OUT <= 0;  //65 / 135 = 0
    16'b01000001_10001000 : OUT <= 0;  //65 / 136 = 0
    16'b01000001_10001001 : OUT <= 0;  //65 / 137 = 0
    16'b01000001_10001010 : OUT <= 0;  //65 / 138 = 0
    16'b01000001_10001011 : OUT <= 0;  //65 / 139 = 0
    16'b01000001_10001100 : OUT <= 0;  //65 / 140 = 0
    16'b01000001_10001101 : OUT <= 0;  //65 / 141 = 0
    16'b01000001_10001110 : OUT <= 0;  //65 / 142 = 0
    16'b01000001_10001111 : OUT <= 0;  //65 / 143 = 0
    16'b01000001_10010000 : OUT <= 0;  //65 / 144 = 0
    16'b01000001_10010001 : OUT <= 0;  //65 / 145 = 0
    16'b01000001_10010010 : OUT <= 0;  //65 / 146 = 0
    16'b01000001_10010011 : OUT <= 0;  //65 / 147 = 0
    16'b01000001_10010100 : OUT <= 0;  //65 / 148 = 0
    16'b01000001_10010101 : OUT <= 0;  //65 / 149 = 0
    16'b01000001_10010110 : OUT <= 0;  //65 / 150 = 0
    16'b01000001_10010111 : OUT <= 0;  //65 / 151 = 0
    16'b01000001_10011000 : OUT <= 0;  //65 / 152 = 0
    16'b01000001_10011001 : OUT <= 0;  //65 / 153 = 0
    16'b01000001_10011010 : OUT <= 0;  //65 / 154 = 0
    16'b01000001_10011011 : OUT <= 0;  //65 / 155 = 0
    16'b01000001_10011100 : OUT <= 0;  //65 / 156 = 0
    16'b01000001_10011101 : OUT <= 0;  //65 / 157 = 0
    16'b01000001_10011110 : OUT <= 0;  //65 / 158 = 0
    16'b01000001_10011111 : OUT <= 0;  //65 / 159 = 0
    16'b01000001_10100000 : OUT <= 0;  //65 / 160 = 0
    16'b01000001_10100001 : OUT <= 0;  //65 / 161 = 0
    16'b01000001_10100010 : OUT <= 0;  //65 / 162 = 0
    16'b01000001_10100011 : OUT <= 0;  //65 / 163 = 0
    16'b01000001_10100100 : OUT <= 0;  //65 / 164 = 0
    16'b01000001_10100101 : OUT <= 0;  //65 / 165 = 0
    16'b01000001_10100110 : OUT <= 0;  //65 / 166 = 0
    16'b01000001_10100111 : OUT <= 0;  //65 / 167 = 0
    16'b01000001_10101000 : OUT <= 0;  //65 / 168 = 0
    16'b01000001_10101001 : OUT <= 0;  //65 / 169 = 0
    16'b01000001_10101010 : OUT <= 0;  //65 / 170 = 0
    16'b01000001_10101011 : OUT <= 0;  //65 / 171 = 0
    16'b01000001_10101100 : OUT <= 0;  //65 / 172 = 0
    16'b01000001_10101101 : OUT <= 0;  //65 / 173 = 0
    16'b01000001_10101110 : OUT <= 0;  //65 / 174 = 0
    16'b01000001_10101111 : OUT <= 0;  //65 / 175 = 0
    16'b01000001_10110000 : OUT <= 0;  //65 / 176 = 0
    16'b01000001_10110001 : OUT <= 0;  //65 / 177 = 0
    16'b01000001_10110010 : OUT <= 0;  //65 / 178 = 0
    16'b01000001_10110011 : OUT <= 0;  //65 / 179 = 0
    16'b01000001_10110100 : OUT <= 0;  //65 / 180 = 0
    16'b01000001_10110101 : OUT <= 0;  //65 / 181 = 0
    16'b01000001_10110110 : OUT <= 0;  //65 / 182 = 0
    16'b01000001_10110111 : OUT <= 0;  //65 / 183 = 0
    16'b01000001_10111000 : OUT <= 0;  //65 / 184 = 0
    16'b01000001_10111001 : OUT <= 0;  //65 / 185 = 0
    16'b01000001_10111010 : OUT <= 0;  //65 / 186 = 0
    16'b01000001_10111011 : OUT <= 0;  //65 / 187 = 0
    16'b01000001_10111100 : OUT <= 0;  //65 / 188 = 0
    16'b01000001_10111101 : OUT <= 0;  //65 / 189 = 0
    16'b01000001_10111110 : OUT <= 0;  //65 / 190 = 0
    16'b01000001_10111111 : OUT <= 0;  //65 / 191 = 0
    16'b01000001_11000000 : OUT <= 0;  //65 / 192 = 0
    16'b01000001_11000001 : OUT <= 0;  //65 / 193 = 0
    16'b01000001_11000010 : OUT <= 0;  //65 / 194 = 0
    16'b01000001_11000011 : OUT <= 0;  //65 / 195 = 0
    16'b01000001_11000100 : OUT <= 0;  //65 / 196 = 0
    16'b01000001_11000101 : OUT <= 0;  //65 / 197 = 0
    16'b01000001_11000110 : OUT <= 0;  //65 / 198 = 0
    16'b01000001_11000111 : OUT <= 0;  //65 / 199 = 0
    16'b01000001_11001000 : OUT <= 0;  //65 / 200 = 0
    16'b01000001_11001001 : OUT <= 0;  //65 / 201 = 0
    16'b01000001_11001010 : OUT <= 0;  //65 / 202 = 0
    16'b01000001_11001011 : OUT <= 0;  //65 / 203 = 0
    16'b01000001_11001100 : OUT <= 0;  //65 / 204 = 0
    16'b01000001_11001101 : OUT <= 0;  //65 / 205 = 0
    16'b01000001_11001110 : OUT <= 0;  //65 / 206 = 0
    16'b01000001_11001111 : OUT <= 0;  //65 / 207 = 0
    16'b01000001_11010000 : OUT <= 0;  //65 / 208 = 0
    16'b01000001_11010001 : OUT <= 0;  //65 / 209 = 0
    16'b01000001_11010010 : OUT <= 0;  //65 / 210 = 0
    16'b01000001_11010011 : OUT <= 0;  //65 / 211 = 0
    16'b01000001_11010100 : OUT <= 0;  //65 / 212 = 0
    16'b01000001_11010101 : OUT <= 0;  //65 / 213 = 0
    16'b01000001_11010110 : OUT <= 0;  //65 / 214 = 0
    16'b01000001_11010111 : OUT <= 0;  //65 / 215 = 0
    16'b01000001_11011000 : OUT <= 0;  //65 / 216 = 0
    16'b01000001_11011001 : OUT <= 0;  //65 / 217 = 0
    16'b01000001_11011010 : OUT <= 0;  //65 / 218 = 0
    16'b01000001_11011011 : OUT <= 0;  //65 / 219 = 0
    16'b01000001_11011100 : OUT <= 0;  //65 / 220 = 0
    16'b01000001_11011101 : OUT <= 0;  //65 / 221 = 0
    16'b01000001_11011110 : OUT <= 0;  //65 / 222 = 0
    16'b01000001_11011111 : OUT <= 0;  //65 / 223 = 0
    16'b01000001_11100000 : OUT <= 0;  //65 / 224 = 0
    16'b01000001_11100001 : OUT <= 0;  //65 / 225 = 0
    16'b01000001_11100010 : OUT <= 0;  //65 / 226 = 0
    16'b01000001_11100011 : OUT <= 0;  //65 / 227 = 0
    16'b01000001_11100100 : OUT <= 0;  //65 / 228 = 0
    16'b01000001_11100101 : OUT <= 0;  //65 / 229 = 0
    16'b01000001_11100110 : OUT <= 0;  //65 / 230 = 0
    16'b01000001_11100111 : OUT <= 0;  //65 / 231 = 0
    16'b01000001_11101000 : OUT <= 0;  //65 / 232 = 0
    16'b01000001_11101001 : OUT <= 0;  //65 / 233 = 0
    16'b01000001_11101010 : OUT <= 0;  //65 / 234 = 0
    16'b01000001_11101011 : OUT <= 0;  //65 / 235 = 0
    16'b01000001_11101100 : OUT <= 0;  //65 / 236 = 0
    16'b01000001_11101101 : OUT <= 0;  //65 / 237 = 0
    16'b01000001_11101110 : OUT <= 0;  //65 / 238 = 0
    16'b01000001_11101111 : OUT <= 0;  //65 / 239 = 0
    16'b01000001_11110000 : OUT <= 0;  //65 / 240 = 0
    16'b01000001_11110001 : OUT <= 0;  //65 / 241 = 0
    16'b01000001_11110010 : OUT <= 0;  //65 / 242 = 0
    16'b01000001_11110011 : OUT <= 0;  //65 / 243 = 0
    16'b01000001_11110100 : OUT <= 0;  //65 / 244 = 0
    16'b01000001_11110101 : OUT <= 0;  //65 / 245 = 0
    16'b01000001_11110110 : OUT <= 0;  //65 / 246 = 0
    16'b01000001_11110111 : OUT <= 0;  //65 / 247 = 0
    16'b01000001_11111000 : OUT <= 0;  //65 / 248 = 0
    16'b01000001_11111001 : OUT <= 0;  //65 / 249 = 0
    16'b01000001_11111010 : OUT <= 0;  //65 / 250 = 0
    16'b01000001_11111011 : OUT <= 0;  //65 / 251 = 0
    16'b01000001_11111100 : OUT <= 0;  //65 / 252 = 0
    16'b01000001_11111101 : OUT <= 0;  //65 / 253 = 0
    16'b01000001_11111110 : OUT <= 0;  //65 / 254 = 0
    16'b01000001_11111111 : OUT <= 0;  //65 / 255 = 0
    16'b01000010_00000000 : OUT <= 0;  //66 / 0 = 0
    16'b01000010_00000001 : OUT <= 66;  //66 / 1 = 66
    16'b01000010_00000010 : OUT <= 33;  //66 / 2 = 33
    16'b01000010_00000011 : OUT <= 22;  //66 / 3 = 22
    16'b01000010_00000100 : OUT <= 16;  //66 / 4 = 16
    16'b01000010_00000101 : OUT <= 13;  //66 / 5 = 13
    16'b01000010_00000110 : OUT <= 11;  //66 / 6 = 11
    16'b01000010_00000111 : OUT <= 9;  //66 / 7 = 9
    16'b01000010_00001000 : OUT <= 8;  //66 / 8 = 8
    16'b01000010_00001001 : OUT <= 7;  //66 / 9 = 7
    16'b01000010_00001010 : OUT <= 6;  //66 / 10 = 6
    16'b01000010_00001011 : OUT <= 6;  //66 / 11 = 6
    16'b01000010_00001100 : OUT <= 5;  //66 / 12 = 5
    16'b01000010_00001101 : OUT <= 5;  //66 / 13 = 5
    16'b01000010_00001110 : OUT <= 4;  //66 / 14 = 4
    16'b01000010_00001111 : OUT <= 4;  //66 / 15 = 4
    16'b01000010_00010000 : OUT <= 4;  //66 / 16 = 4
    16'b01000010_00010001 : OUT <= 3;  //66 / 17 = 3
    16'b01000010_00010010 : OUT <= 3;  //66 / 18 = 3
    16'b01000010_00010011 : OUT <= 3;  //66 / 19 = 3
    16'b01000010_00010100 : OUT <= 3;  //66 / 20 = 3
    16'b01000010_00010101 : OUT <= 3;  //66 / 21 = 3
    16'b01000010_00010110 : OUT <= 3;  //66 / 22 = 3
    16'b01000010_00010111 : OUT <= 2;  //66 / 23 = 2
    16'b01000010_00011000 : OUT <= 2;  //66 / 24 = 2
    16'b01000010_00011001 : OUT <= 2;  //66 / 25 = 2
    16'b01000010_00011010 : OUT <= 2;  //66 / 26 = 2
    16'b01000010_00011011 : OUT <= 2;  //66 / 27 = 2
    16'b01000010_00011100 : OUT <= 2;  //66 / 28 = 2
    16'b01000010_00011101 : OUT <= 2;  //66 / 29 = 2
    16'b01000010_00011110 : OUT <= 2;  //66 / 30 = 2
    16'b01000010_00011111 : OUT <= 2;  //66 / 31 = 2
    16'b01000010_00100000 : OUT <= 2;  //66 / 32 = 2
    16'b01000010_00100001 : OUT <= 2;  //66 / 33 = 2
    16'b01000010_00100010 : OUT <= 1;  //66 / 34 = 1
    16'b01000010_00100011 : OUT <= 1;  //66 / 35 = 1
    16'b01000010_00100100 : OUT <= 1;  //66 / 36 = 1
    16'b01000010_00100101 : OUT <= 1;  //66 / 37 = 1
    16'b01000010_00100110 : OUT <= 1;  //66 / 38 = 1
    16'b01000010_00100111 : OUT <= 1;  //66 / 39 = 1
    16'b01000010_00101000 : OUT <= 1;  //66 / 40 = 1
    16'b01000010_00101001 : OUT <= 1;  //66 / 41 = 1
    16'b01000010_00101010 : OUT <= 1;  //66 / 42 = 1
    16'b01000010_00101011 : OUT <= 1;  //66 / 43 = 1
    16'b01000010_00101100 : OUT <= 1;  //66 / 44 = 1
    16'b01000010_00101101 : OUT <= 1;  //66 / 45 = 1
    16'b01000010_00101110 : OUT <= 1;  //66 / 46 = 1
    16'b01000010_00101111 : OUT <= 1;  //66 / 47 = 1
    16'b01000010_00110000 : OUT <= 1;  //66 / 48 = 1
    16'b01000010_00110001 : OUT <= 1;  //66 / 49 = 1
    16'b01000010_00110010 : OUT <= 1;  //66 / 50 = 1
    16'b01000010_00110011 : OUT <= 1;  //66 / 51 = 1
    16'b01000010_00110100 : OUT <= 1;  //66 / 52 = 1
    16'b01000010_00110101 : OUT <= 1;  //66 / 53 = 1
    16'b01000010_00110110 : OUT <= 1;  //66 / 54 = 1
    16'b01000010_00110111 : OUT <= 1;  //66 / 55 = 1
    16'b01000010_00111000 : OUT <= 1;  //66 / 56 = 1
    16'b01000010_00111001 : OUT <= 1;  //66 / 57 = 1
    16'b01000010_00111010 : OUT <= 1;  //66 / 58 = 1
    16'b01000010_00111011 : OUT <= 1;  //66 / 59 = 1
    16'b01000010_00111100 : OUT <= 1;  //66 / 60 = 1
    16'b01000010_00111101 : OUT <= 1;  //66 / 61 = 1
    16'b01000010_00111110 : OUT <= 1;  //66 / 62 = 1
    16'b01000010_00111111 : OUT <= 1;  //66 / 63 = 1
    16'b01000010_01000000 : OUT <= 1;  //66 / 64 = 1
    16'b01000010_01000001 : OUT <= 1;  //66 / 65 = 1
    16'b01000010_01000010 : OUT <= 1;  //66 / 66 = 1
    16'b01000010_01000011 : OUT <= 0;  //66 / 67 = 0
    16'b01000010_01000100 : OUT <= 0;  //66 / 68 = 0
    16'b01000010_01000101 : OUT <= 0;  //66 / 69 = 0
    16'b01000010_01000110 : OUT <= 0;  //66 / 70 = 0
    16'b01000010_01000111 : OUT <= 0;  //66 / 71 = 0
    16'b01000010_01001000 : OUT <= 0;  //66 / 72 = 0
    16'b01000010_01001001 : OUT <= 0;  //66 / 73 = 0
    16'b01000010_01001010 : OUT <= 0;  //66 / 74 = 0
    16'b01000010_01001011 : OUT <= 0;  //66 / 75 = 0
    16'b01000010_01001100 : OUT <= 0;  //66 / 76 = 0
    16'b01000010_01001101 : OUT <= 0;  //66 / 77 = 0
    16'b01000010_01001110 : OUT <= 0;  //66 / 78 = 0
    16'b01000010_01001111 : OUT <= 0;  //66 / 79 = 0
    16'b01000010_01010000 : OUT <= 0;  //66 / 80 = 0
    16'b01000010_01010001 : OUT <= 0;  //66 / 81 = 0
    16'b01000010_01010010 : OUT <= 0;  //66 / 82 = 0
    16'b01000010_01010011 : OUT <= 0;  //66 / 83 = 0
    16'b01000010_01010100 : OUT <= 0;  //66 / 84 = 0
    16'b01000010_01010101 : OUT <= 0;  //66 / 85 = 0
    16'b01000010_01010110 : OUT <= 0;  //66 / 86 = 0
    16'b01000010_01010111 : OUT <= 0;  //66 / 87 = 0
    16'b01000010_01011000 : OUT <= 0;  //66 / 88 = 0
    16'b01000010_01011001 : OUT <= 0;  //66 / 89 = 0
    16'b01000010_01011010 : OUT <= 0;  //66 / 90 = 0
    16'b01000010_01011011 : OUT <= 0;  //66 / 91 = 0
    16'b01000010_01011100 : OUT <= 0;  //66 / 92 = 0
    16'b01000010_01011101 : OUT <= 0;  //66 / 93 = 0
    16'b01000010_01011110 : OUT <= 0;  //66 / 94 = 0
    16'b01000010_01011111 : OUT <= 0;  //66 / 95 = 0
    16'b01000010_01100000 : OUT <= 0;  //66 / 96 = 0
    16'b01000010_01100001 : OUT <= 0;  //66 / 97 = 0
    16'b01000010_01100010 : OUT <= 0;  //66 / 98 = 0
    16'b01000010_01100011 : OUT <= 0;  //66 / 99 = 0
    16'b01000010_01100100 : OUT <= 0;  //66 / 100 = 0
    16'b01000010_01100101 : OUT <= 0;  //66 / 101 = 0
    16'b01000010_01100110 : OUT <= 0;  //66 / 102 = 0
    16'b01000010_01100111 : OUT <= 0;  //66 / 103 = 0
    16'b01000010_01101000 : OUT <= 0;  //66 / 104 = 0
    16'b01000010_01101001 : OUT <= 0;  //66 / 105 = 0
    16'b01000010_01101010 : OUT <= 0;  //66 / 106 = 0
    16'b01000010_01101011 : OUT <= 0;  //66 / 107 = 0
    16'b01000010_01101100 : OUT <= 0;  //66 / 108 = 0
    16'b01000010_01101101 : OUT <= 0;  //66 / 109 = 0
    16'b01000010_01101110 : OUT <= 0;  //66 / 110 = 0
    16'b01000010_01101111 : OUT <= 0;  //66 / 111 = 0
    16'b01000010_01110000 : OUT <= 0;  //66 / 112 = 0
    16'b01000010_01110001 : OUT <= 0;  //66 / 113 = 0
    16'b01000010_01110010 : OUT <= 0;  //66 / 114 = 0
    16'b01000010_01110011 : OUT <= 0;  //66 / 115 = 0
    16'b01000010_01110100 : OUT <= 0;  //66 / 116 = 0
    16'b01000010_01110101 : OUT <= 0;  //66 / 117 = 0
    16'b01000010_01110110 : OUT <= 0;  //66 / 118 = 0
    16'b01000010_01110111 : OUT <= 0;  //66 / 119 = 0
    16'b01000010_01111000 : OUT <= 0;  //66 / 120 = 0
    16'b01000010_01111001 : OUT <= 0;  //66 / 121 = 0
    16'b01000010_01111010 : OUT <= 0;  //66 / 122 = 0
    16'b01000010_01111011 : OUT <= 0;  //66 / 123 = 0
    16'b01000010_01111100 : OUT <= 0;  //66 / 124 = 0
    16'b01000010_01111101 : OUT <= 0;  //66 / 125 = 0
    16'b01000010_01111110 : OUT <= 0;  //66 / 126 = 0
    16'b01000010_01111111 : OUT <= 0;  //66 / 127 = 0
    16'b01000010_10000000 : OUT <= 0;  //66 / 128 = 0
    16'b01000010_10000001 : OUT <= 0;  //66 / 129 = 0
    16'b01000010_10000010 : OUT <= 0;  //66 / 130 = 0
    16'b01000010_10000011 : OUT <= 0;  //66 / 131 = 0
    16'b01000010_10000100 : OUT <= 0;  //66 / 132 = 0
    16'b01000010_10000101 : OUT <= 0;  //66 / 133 = 0
    16'b01000010_10000110 : OUT <= 0;  //66 / 134 = 0
    16'b01000010_10000111 : OUT <= 0;  //66 / 135 = 0
    16'b01000010_10001000 : OUT <= 0;  //66 / 136 = 0
    16'b01000010_10001001 : OUT <= 0;  //66 / 137 = 0
    16'b01000010_10001010 : OUT <= 0;  //66 / 138 = 0
    16'b01000010_10001011 : OUT <= 0;  //66 / 139 = 0
    16'b01000010_10001100 : OUT <= 0;  //66 / 140 = 0
    16'b01000010_10001101 : OUT <= 0;  //66 / 141 = 0
    16'b01000010_10001110 : OUT <= 0;  //66 / 142 = 0
    16'b01000010_10001111 : OUT <= 0;  //66 / 143 = 0
    16'b01000010_10010000 : OUT <= 0;  //66 / 144 = 0
    16'b01000010_10010001 : OUT <= 0;  //66 / 145 = 0
    16'b01000010_10010010 : OUT <= 0;  //66 / 146 = 0
    16'b01000010_10010011 : OUT <= 0;  //66 / 147 = 0
    16'b01000010_10010100 : OUT <= 0;  //66 / 148 = 0
    16'b01000010_10010101 : OUT <= 0;  //66 / 149 = 0
    16'b01000010_10010110 : OUT <= 0;  //66 / 150 = 0
    16'b01000010_10010111 : OUT <= 0;  //66 / 151 = 0
    16'b01000010_10011000 : OUT <= 0;  //66 / 152 = 0
    16'b01000010_10011001 : OUT <= 0;  //66 / 153 = 0
    16'b01000010_10011010 : OUT <= 0;  //66 / 154 = 0
    16'b01000010_10011011 : OUT <= 0;  //66 / 155 = 0
    16'b01000010_10011100 : OUT <= 0;  //66 / 156 = 0
    16'b01000010_10011101 : OUT <= 0;  //66 / 157 = 0
    16'b01000010_10011110 : OUT <= 0;  //66 / 158 = 0
    16'b01000010_10011111 : OUT <= 0;  //66 / 159 = 0
    16'b01000010_10100000 : OUT <= 0;  //66 / 160 = 0
    16'b01000010_10100001 : OUT <= 0;  //66 / 161 = 0
    16'b01000010_10100010 : OUT <= 0;  //66 / 162 = 0
    16'b01000010_10100011 : OUT <= 0;  //66 / 163 = 0
    16'b01000010_10100100 : OUT <= 0;  //66 / 164 = 0
    16'b01000010_10100101 : OUT <= 0;  //66 / 165 = 0
    16'b01000010_10100110 : OUT <= 0;  //66 / 166 = 0
    16'b01000010_10100111 : OUT <= 0;  //66 / 167 = 0
    16'b01000010_10101000 : OUT <= 0;  //66 / 168 = 0
    16'b01000010_10101001 : OUT <= 0;  //66 / 169 = 0
    16'b01000010_10101010 : OUT <= 0;  //66 / 170 = 0
    16'b01000010_10101011 : OUT <= 0;  //66 / 171 = 0
    16'b01000010_10101100 : OUT <= 0;  //66 / 172 = 0
    16'b01000010_10101101 : OUT <= 0;  //66 / 173 = 0
    16'b01000010_10101110 : OUT <= 0;  //66 / 174 = 0
    16'b01000010_10101111 : OUT <= 0;  //66 / 175 = 0
    16'b01000010_10110000 : OUT <= 0;  //66 / 176 = 0
    16'b01000010_10110001 : OUT <= 0;  //66 / 177 = 0
    16'b01000010_10110010 : OUT <= 0;  //66 / 178 = 0
    16'b01000010_10110011 : OUT <= 0;  //66 / 179 = 0
    16'b01000010_10110100 : OUT <= 0;  //66 / 180 = 0
    16'b01000010_10110101 : OUT <= 0;  //66 / 181 = 0
    16'b01000010_10110110 : OUT <= 0;  //66 / 182 = 0
    16'b01000010_10110111 : OUT <= 0;  //66 / 183 = 0
    16'b01000010_10111000 : OUT <= 0;  //66 / 184 = 0
    16'b01000010_10111001 : OUT <= 0;  //66 / 185 = 0
    16'b01000010_10111010 : OUT <= 0;  //66 / 186 = 0
    16'b01000010_10111011 : OUT <= 0;  //66 / 187 = 0
    16'b01000010_10111100 : OUT <= 0;  //66 / 188 = 0
    16'b01000010_10111101 : OUT <= 0;  //66 / 189 = 0
    16'b01000010_10111110 : OUT <= 0;  //66 / 190 = 0
    16'b01000010_10111111 : OUT <= 0;  //66 / 191 = 0
    16'b01000010_11000000 : OUT <= 0;  //66 / 192 = 0
    16'b01000010_11000001 : OUT <= 0;  //66 / 193 = 0
    16'b01000010_11000010 : OUT <= 0;  //66 / 194 = 0
    16'b01000010_11000011 : OUT <= 0;  //66 / 195 = 0
    16'b01000010_11000100 : OUT <= 0;  //66 / 196 = 0
    16'b01000010_11000101 : OUT <= 0;  //66 / 197 = 0
    16'b01000010_11000110 : OUT <= 0;  //66 / 198 = 0
    16'b01000010_11000111 : OUT <= 0;  //66 / 199 = 0
    16'b01000010_11001000 : OUT <= 0;  //66 / 200 = 0
    16'b01000010_11001001 : OUT <= 0;  //66 / 201 = 0
    16'b01000010_11001010 : OUT <= 0;  //66 / 202 = 0
    16'b01000010_11001011 : OUT <= 0;  //66 / 203 = 0
    16'b01000010_11001100 : OUT <= 0;  //66 / 204 = 0
    16'b01000010_11001101 : OUT <= 0;  //66 / 205 = 0
    16'b01000010_11001110 : OUT <= 0;  //66 / 206 = 0
    16'b01000010_11001111 : OUT <= 0;  //66 / 207 = 0
    16'b01000010_11010000 : OUT <= 0;  //66 / 208 = 0
    16'b01000010_11010001 : OUT <= 0;  //66 / 209 = 0
    16'b01000010_11010010 : OUT <= 0;  //66 / 210 = 0
    16'b01000010_11010011 : OUT <= 0;  //66 / 211 = 0
    16'b01000010_11010100 : OUT <= 0;  //66 / 212 = 0
    16'b01000010_11010101 : OUT <= 0;  //66 / 213 = 0
    16'b01000010_11010110 : OUT <= 0;  //66 / 214 = 0
    16'b01000010_11010111 : OUT <= 0;  //66 / 215 = 0
    16'b01000010_11011000 : OUT <= 0;  //66 / 216 = 0
    16'b01000010_11011001 : OUT <= 0;  //66 / 217 = 0
    16'b01000010_11011010 : OUT <= 0;  //66 / 218 = 0
    16'b01000010_11011011 : OUT <= 0;  //66 / 219 = 0
    16'b01000010_11011100 : OUT <= 0;  //66 / 220 = 0
    16'b01000010_11011101 : OUT <= 0;  //66 / 221 = 0
    16'b01000010_11011110 : OUT <= 0;  //66 / 222 = 0
    16'b01000010_11011111 : OUT <= 0;  //66 / 223 = 0
    16'b01000010_11100000 : OUT <= 0;  //66 / 224 = 0
    16'b01000010_11100001 : OUT <= 0;  //66 / 225 = 0
    16'b01000010_11100010 : OUT <= 0;  //66 / 226 = 0
    16'b01000010_11100011 : OUT <= 0;  //66 / 227 = 0
    16'b01000010_11100100 : OUT <= 0;  //66 / 228 = 0
    16'b01000010_11100101 : OUT <= 0;  //66 / 229 = 0
    16'b01000010_11100110 : OUT <= 0;  //66 / 230 = 0
    16'b01000010_11100111 : OUT <= 0;  //66 / 231 = 0
    16'b01000010_11101000 : OUT <= 0;  //66 / 232 = 0
    16'b01000010_11101001 : OUT <= 0;  //66 / 233 = 0
    16'b01000010_11101010 : OUT <= 0;  //66 / 234 = 0
    16'b01000010_11101011 : OUT <= 0;  //66 / 235 = 0
    16'b01000010_11101100 : OUT <= 0;  //66 / 236 = 0
    16'b01000010_11101101 : OUT <= 0;  //66 / 237 = 0
    16'b01000010_11101110 : OUT <= 0;  //66 / 238 = 0
    16'b01000010_11101111 : OUT <= 0;  //66 / 239 = 0
    16'b01000010_11110000 : OUT <= 0;  //66 / 240 = 0
    16'b01000010_11110001 : OUT <= 0;  //66 / 241 = 0
    16'b01000010_11110010 : OUT <= 0;  //66 / 242 = 0
    16'b01000010_11110011 : OUT <= 0;  //66 / 243 = 0
    16'b01000010_11110100 : OUT <= 0;  //66 / 244 = 0
    16'b01000010_11110101 : OUT <= 0;  //66 / 245 = 0
    16'b01000010_11110110 : OUT <= 0;  //66 / 246 = 0
    16'b01000010_11110111 : OUT <= 0;  //66 / 247 = 0
    16'b01000010_11111000 : OUT <= 0;  //66 / 248 = 0
    16'b01000010_11111001 : OUT <= 0;  //66 / 249 = 0
    16'b01000010_11111010 : OUT <= 0;  //66 / 250 = 0
    16'b01000010_11111011 : OUT <= 0;  //66 / 251 = 0
    16'b01000010_11111100 : OUT <= 0;  //66 / 252 = 0
    16'b01000010_11111101 : OUT <= 0;  //66 / 253 = 0
    16'b01000010_11111110 : OUT <= 0;  //66 / 254 = 0
    16'b01000010_11111111 : OUT <= 0;  //66 / 255 = 0
    16'b01000011_00000000 : OUT <= 0;  //67 / 0 = 0
    16'b01000011_00000001 : OUT <= 67;  //67 / 1 = 67
    16'b01000011_00000010 : OUT <= 33;  //67 / 2 = 33
    16'b01000011_00000011 : OUT <= 22;  //67 / 3 = 22
    16'b01000011_00000100 : OUT <= 16;  //67 / 4 = 16
    16'b01000011_00000101 : OUT <= 13;  //67 / 5 = 13
    16'b01000011_00000110 : OUT <= 11;  //67 / 6 = 11
    16'b01000011_00000111 : OUT <= 9;  //67 / 7 = 9
    16'b01000011_00001000 : OUT <= 8;  //67 / 8 = 8
    16'b01000011_00001001 : OUT <= 7;  //67 / 9 = 7
    16'b01000011_00001010 : OUT <= 6;  //67 / 10 = 6
    16'b01000011_00001011 : OUT <= 6;  //67 / 11 = 6
    16'b01000011_00001100 : OUT <= 5;  //67 / 12 = 5
    16'b01000011_00001101 : OUT <= 5;  //67 / 13 = 5
    16'b01000011_00001110 : OUT <= 4;  //67 / 14 = 4
    16'b01000011_00001111 : OUT <= 4;  //67 / 15 = 4
    16'b01000011_00010000 : OUT <= 4;  //67 / 16 = 4
    16'b01000011_00010001 : OUT <= 3;  //67 / 17 = 3
    16'b01000011_00010010 : OUT <= 3;  //67 / 18 = 3
    16'b01000011_00010011 : OUT <= 3;  //67 / 19 = 3
    16'b01000011_00010100 : OUT <= 3;  //67 / 20 = 3
    16'b01000011_00010101 : OUT <= 3;  //67 / 21 = 3
    16'b01000011_00010110 : OUT <= 3;  //67 / 22 = 3
    16'b01000011_00010111 : OUT <= 2;  //67 / 23 = 2
    16'b01000011_00011000 : OUT <= 2;  //67 / 24 = 2
    16'b01000011_00011001 : OUT <= 2;  //67 / 25 = 2
    16'b01000011_00011010 : OUT <= 2;  //67 / 26 = 2
    16'b01000011_00011011 : OUT <= 2;  //67 / 27 = 2
    16'b01000011_00011100 : OUT <= 2;  //67 / 28 = 2
    16'b01000011_00011101 : OUT <= 2;  //67 / 29 = 2
    16'b01000011_00011110 : OUT <= 2;  //67 / 30 = 2
    16'b01000011_00011111 : OUT <= 2;  //67 / 31 = 2
    16'b01000011_00100000 : OUT <= 2;  //67 / 32 = 2
    16'b01000011_00100001 : OUT <= 2;  //67 / 33 = 2
    16'b01000011_00100010 : OUT <= 1;  //67 / 34 = 1
    16'b01000011_00100011 : OUT <= 1;  //67 / 35 = 1
    16'b01000011_00100100 : OUT <= 1;  //67 / 36 = 1
    16'b01000011_00100101 : OUT <= 1;  //67 / 37 = 1
    16'b01000011_00100110 : OUT <= 1;  //67 / 38 = 1
    16'b01000011_00100111 : OUT <= 1;  //67 / 39 = 1
    16'b01000011_00101000 : OUT <= 1;  //67 / 40 = 1
    16'b01000011_00101001 : OUT <= 1;  //67 / 41 = 1
    16'b01000011_00101010 : OUT <= 1;  //67 / 42 = 1
    16'b01000011_00101011 : OUT <= 1;  //67 / 43 = 1
    16'b01000011_00101100 : OUT <= 1;  //67 / 44 = 1
    16'b01000011_00101101 : OUT <= 1;  //67 / 45 = 1
    16'b01000011_00101110 : OUT <= 1;  //67 / 46 = 1
    16'b01000011_00101111 : OUT <= 1;  //67 / 47 = 1
    16'b01000011_00110000 : OUT <= 1;  //67 / 48 = 1
    16'b01000011_00110001 : OUT <= 1;  //67 / 49 = 1
    16'b01000011_00110010 : OUT <= 1;  //67 / 50 = 1
    16'b01000011_00110011 : OUT <= 1;  //67 / 51 = 1
    16'b01000011_00110100 : OUT <= 1;  //67 / 52 = 1
    16'b01000011_00110101 : OUT <= 1;  //67 / 53 = 1
    16'b01000011_00110110 : OUT <= 1;  //67 / 54 = 1
    16'b01000011_00110111 : OUT <= 1;  //67 / 55 = 1
    16'b01000011_00111000 : OUT <= 1;  //67 / 56 = 1
    16'b01000011_00111001 : OUT <= 1;  //67 / 57 = 1
    16'b01000011_00111010 : OUT <= 1;  //67 / 58 = 1
    16'b01000011_00111011 : OUT <= 1;  //67 / 59 = 1
    16'b01000011_00111100 : OUT <= 1;  //67 / 60 = 1
    16'b01000011_00111101 : OUT <= 1;  //67 / 61 = 1
    16'b01000011_00111110 : OUT <= 1;  //67 / 62 = 1
    16'b01000011_00111111 : OUT <= 1;  //67 / 63 = 1
    16'b01000011_01000000 : OUT <= 1;  //67 / 64 = 1
    16'b01000011_01000001 : OUT <= 1;  //67 / 65 = 1
    16'b01000011_01000010 : OUT <= 1;  //67 / 66 = 1
    16'b01000011_01000011 : OUT <= 1;  //67 / 67 = 1
    16'b01000011_01000100 : OUT <= 0;  //67 / 68 = 0
    16'b01000011_01000101 : OUT <= 0;  //67 / 69 = 0
    16'b01000011_01000110 : OUT <= 0;  //67 / 70 = 0
    16'b01000011_01000111 : OUT <= 0;  //67 / 71 = 0
    16'b01000011_01001000 : OUT <= 0;  //67 / 72 = 0
    16'b01000011_01001001 : OUT <= 0;  //67 / 73 = 0
    16'b01000011_01001010 : OUT <= 0;  //67 / 74 = 0
    16'b01000011_01001011 : OUT <= 0;  //67 / 75 = 0
    16'b01000011_01001100 : OUT <= 0;  //67 / 76 = 0
    16'b01000011_01001101 : OUT <= 0;  //67 / 77 = 0
    16'b01000011_01001110 : OUT <= 0;  //67 / 78 = 0
    16'b01000011_01001111 : OUT <= 0;  //67 / 79 = 0
    16'b01000011_01010000 : OUT <= 0;  //67 / 80 = 0
    16'b01000011_01010001 : OUT <= 0;  //67 / 81 = 0
    16'b01000011_01010010 : OUT <= 0;  //67 / 82 = 0
    16'b01000011_01010011 : OUT <= 0;  //67 / 83 = 0
    16'b01000011_01010100 : OUT <= 0;  //67 / 84 = 0
    16'b01000011_01010101 : OUT <= 0;  //67 / 85 = 0
    16'b01000011_01010110 : OUT <= 0;  //67 / 86 = 0
    16'b01000011_01010111 : OUT <= 0;  //67 / 87 = 0
    16'b01000011_01011000 : OUT <= 0;  //67 / 88 = 0
    16'b01000011_01011001 : OUT <= 0;  //67 / 89 = 0
    16'b01000011_01011010 : OUT <= 0;  //67 / 90 = 0
    16'b01000011_01011011 : OUT <= 0;  //67 / 91 = 0
    16'b01000011_01011100 : OUT <= 0;  //67 / 92 = 0
    16'b01000011_01011101 : OUT <= 0;  //67 / 93 = 0
    16'b01000011_01011110 : OUT <= 0;  //67 / 94 = 0
    16'b01000011_01011111 : OUT <= 0;  //67 / 95 = 0
    16'b01000011_01100000 : OUT <= 0;  //67 / 96 = 0
    16'b01000011_01100001 : OUT <= 0;  //67 / 97 = 0
    16'b01000011_01100010 : OUT <= 0;  //67 / 98 = 0
    16'b01000011_01100011 : OUT <= 0;  //67 / 99 = 0
    16'b01000011_01100100 : OUT <= 0;  //67 / 100 = 0
    16'b01000011_01100101 : OUT <= 0;  //67 / 101 = 0
    16'b01000011_01100110 : OUT <= 0;  //67 / 102 = 0
    16'b01000011_01100111 : OUT <= 0;  //67 / 103 = 0
    16'b01000011_01101000 : OUT <= 0;  //67 / 104 = 0
    16'b01000011_01101001 : OUT <= 0;  //67 / 105 = 0
    16'b01000011_01101010 : OUT <= 0;  //67 / 106 = 0
    16'b01000011_01101011 : OUT <= 0;  //67 / 107 = 0
    16'b01000011_01101100 : OUT <= 0;  //67 / 108 = 0
    16'b01000011_01101101 : OUT <= 0;  //67 / 109 = 0
    16'b01000011_01101110 : OUT <= 0;  //67 / 110 = 0
    16'b01000011_01101111 : OUT <= 0;  //67 / 111 = 0
    16'b01000011_01110000 : OUT <= 0;  //67 / 112 = 0
    16'b01000011_01110001 : OUT <= 0;  //67 / 113 = 0
    16'b01000011_01110010 : OUT <= 0;  //67 / 114 = 0
    16'b01000011_01110011 : OUT <= 0;  //67 / 115 = 0
    16'b01000011_01110100 : OUT <= 0;  //67 / 116 = 0
    16'b01000011_01110101 : OUT <= 0;  //67 / 117 = 0
    16'b01000011_01110110 : OUT <= 0;  //67 / 118 = 0
    16'b01000011_01110111 : OUT <= 0;  //67 / 119 = 0
    16'b01000011_01111000 : OUT <= 0;  //67 / 120 = 0
    16'b01000011_01111001 : OUT <= 0;  //67 / 121 = 0
    16'b01000011_01111010 : OUT <= 0;  //67 / 122 = 0
    16'b01000011_01111011 : OUT <= 0;  //67 / 123 = 0
    16'b01000011_01111100 : OUT <= 0;  //67 / 124 = 0
    16'b01000011_01111101 : OUT <= 0;  //67 / 125 = 0
    16'b01000011_01111110 : OUT <= 0;  //67 / 126 = 0
    16'b01000011_01111111 : OUT <= 0;  //67 / 127 = 0
    16'b01000011_10000000 : OUT <= 0;  //67 / 128 = 0
    16'b01000011_10000001 : OUT <= 0;  //67 / 129 = 0
    16'b01000011_10000010 : OUT <= 0;  //67 / 130 = 0
    16'b01000011_10000011 : OUT <= 0;  //67 / 131 = 0
    16'b01000011_10000100 : OUT <= 0;  //67 / 132 = 0
    16'b01000011_10000101 : OUT <= 0;  //67 / 133 = 0
    16'b01000011_10000110 : OUT <= 0;  //67 / 134 = 0
    16'b01000011_10000111 : OUT <= 0;  //67 / 135 = 0
    16'b01000011_10001000 : OUT <= 0;  //67 / 136 = 0
    16'b01000011_10001001 : OUT <= 0;  //67 / 137 = 0
    16'b01000011_10001010 : OUT <= 0;  //67 / 138 = 0
    16'b01000011_10001011 : OUT <= 0;  //67 / 139 = 0
    16'b01000011_10001100 : OUT <= 0;  //67 / 140 = 0
    16'b01000011_10001101 : OUT <= 0;  //67 / 141 = 0
    16'b01000011_10001110 : OUT <= 0;  //67 / 142 = 0
    16'b01000011_10001111 : OUT <= 0;  //67 / 143 = 0
    16'b01000011_10010000 : OUT <= 0;  //67 / 144 = 0
    16'b01000011_10010001 : OUT <= 0;  //67 / 145 = 0
    16'b01000011_10010010 : OUT <= 0;  //67 / 146 = 0
    16'b01000011_10010011 : OUT <= 0;  //67 / 147 = 0
    16'b01000011_10010100 : OUT <= 0;  //67 / 148 = 0
    16'b01000011_10010101 : OUT <= 0;  //67 / 149 = 0
    16'b01000011_10010110 : OUT <= 0;  //67 / 150 = 0
    16'b01000011_10010111 : OUT <= 0;  //67 / 151 = 0
    16'b01000011_10011000 : OUT <= 0;  //67 / 152 = 0
    16'b01000011_10011001 : OUT <= 0;  //67 / 153 = 0
    16'b01000011_10011010 : OUT <= 0;  //67 / 154 = 0
    16'b01000011_10011011 : OUT <= 0;  //67 / 155 = 0
    16'b01000011_10011100 : OUT <= 0;  //67 / 156 = 0
    16'b01000011_10011101 : OUT <= 0;  //67 / 157 = 0
    16'b01000011_10011110 : OUT <= 0;  //67 / 158 = 0
    16'b01000011_10011111 : OUT <= 0;  //67 / 159 = 0
    16'b01000011_10100000 : OUT <= 0;  //67 / 160 = 0
    16'b01000011_10100001 : OUT <= 0;  //67 / 161 = 0
    16'b01000011_10100010 : OUT <= 0;  //67 / 162 = 0
    16'b01000011_10100011 : OUT <= 0;  //67 / 163 = 0
    16'b01000011_10100100 : OUT <= 0;  //67 / 164 = 0
    16'b01000011_10100101 : OUT <= 0;  //67 / 165 = 0
    16'b01000011_10100110 : OUT <= 0;  //67 / 166 = 0
    16'b01000011_10100111 : OUT <= 0;  //67 / 167 = 0
    16'b01000011_10101000 : OUT <= 0;  //67 / 168 = 0
    16'b01000011_10101001 : OUT <= 0;  //67 / 169 = 0
    16'b01000011_10101010 : OUT <= 0;  //67 / 170 = 0
    16'b01000011_10101011 : OUT <= 0;  //67 / 171 = 0
    16'b01000011_10101100 : OUT <= 0;  //67 / 172 = 0
    16'b01000011_10101101 : OUT <= 0;  //67 / 173 = 0
    16'b01000011_10101110 : OUT <= 0;  //67 / 174 = 0
    16'b01000011_10101111 : OUT <= 0;  //67 / 175 = 0
    16'b01000011_10110000 : OUT <= 0;  //67 / 176 = 0
    16'b01000011_10110001 : OUT <= 0;  //67 / 177 = 0
    16'b01000011_10110010 : OUT <= 0;  //67 / 178 = 0
    16'b01000011_10110011 : OUT <= 0;  //67 / 179 = 0
    16'b01000011_10110100 : OUT <= 0;  //67 / 180 = 0
    16'b01000011_10110101 : OUT <= 0;  //67 / 181 = 0
    16'b01000011_10110110 : OUT <= 0;  //67 / 182 = 0
    16'b01000011_10110111 : OUT <= 0;  //67 / 183 = 0
    16'b01000011_10111000 : OUT <= 0;  //67 / 184 = 0
    16'b01000011_10111001 : OUT <= 0;  //67 / 185 = 0
    16'b01000011_10111010 : OUT <= 0;  //67 / 186 = 0
    16'b01000011_10111011 : OUT <= 0;  //67 / 187 = 0
    16'b01000011_10111100 : OUT <= 0;  //67 / 188 = 0
    16'b01000011_10111101 : OUT <= 0;  //67 / 189 = 0
    16'b01000011_10111110 : OUT <= 0;  //67 / 190 = 0
    16'b01000011_10111111 : OUT <= 0;  //67 / 191 = 0
    16'b01000011_11000000 : OUT <= 0;  //67 / 192 = 0
    16'b01000011_11000001 : OUT <= 0;  //67 / 193 = 0
    16'b01000011_11000010 : OUT <= 0;  //67 / 194 = 0
    16'b01000011_11000011 : OUT <= 0;  //67 / 195 = 0
    16'b01000011_11000100 : OUT <= 0;  //67 / 196 = 0
    16'b01000011_11000101 : OUT <= 0;  //67 / 197 = 0
    16'b01000011_11000110 : OUT <= 0;  //67 / 198 = 0
    16'b01000011_11000111 : OUT <= 0;  //67 / 199 = 0
    16'b01000011_11001000 : OUT <= 0;  //67 / 200 = 0
    16'b01000011_11001001 : OUT <= 0;  //67 / 201 = 0
    16'b01000011_11001010 : OUT <= 0;  //67 / 202 = 0
    16'b01000011_11001011 : OUT <= 0;  //67 / 203 = 0
    16'b01000011_11001100 : OUT <= 0;  //67 / 204 = 0
    16'b01000011_11001101 : OUT <= 0;  //67 / 205 = 0
    16'b01000011_11001110 : OUT <= 0;  //67 / 206 = 0
    16'b01000011_11001111 : OUT <= 0;  //67 / 207 = 0
    16'b01000011_11010000 : OUT <= 0;  //67 / 208 = 0
    16'b01000011_11010001 : OUT <= 0;  //67 / 209 = 0
    16'b01000011_11010010 : OUT <= 0;  //67 / 210 = 0
    16'b01000011_11010011 : OUT <= 0;  //67 / 211 = 0
    16'b01000011_11010100 : OUT <= 0;  //67 / 212 = 0
    16'b01000011_11010101 : OUT <= 0;  //67 / 213 = 0
    16'b01000011_11010110 : OUT <= 0;  //67 / 214 = 0
    16'b01000011_11010111 : OUT <= 0;  //67 / 215 = 0
    16'b01000011_11011000 : OUT <= 0;  //67 / 216 = 0
    16'b01000011_11011001 : OUT <= 0;  //67 / 217 = 0
    16'b01000011_11011010 : OUT <= 0;  //67 / 218 = 0
    16'b01000011_11011011 : OUT <= 0;  //67 / 219 = 0
    16'b01000011_11011100 : OUT <= 0;  //67 / 220 = 0
    16'b01000011_11011101 : OUT <= 0;  //67 / 221 = 0
    16'b01000011_11011110 : OUT <= 0;  //67 / 222 = 0
    16'b01000011_11011111 : OUT <= 0;  //67 / 223 = 0
    16'b01000011_11100000 : OUT <= 0;  //67 / 224 = 0
    16'b01000011_11100001 : OUT <= 0;  //67 / 225 = 0
    16'b01000011_11100010 : OUT <= 0;  //67 / 226 = 0
    16'b01000011_11100011 : OUT <= 0;  //67 / 227 = 0
    16'b01000011_11100100 : OUT <= 0;  //67 / 228 = 0
    16'b01000011_11100101 : OUT <= 0;  //67 / 229 = 0
    16'b01000011_11100110 : OUT <= 0;  //67 / 230 = 0
    16'b01000011_11100111 : OUT <= 0;  //67 / 231 = 0
    16'b01000011_11101000 : OUT <= 0;  //67 / 232 = 0
    16'b01000011_11101001 : OUT <= 0;  //67 / 233 = 0
    16'b01000011_11101010 : OUT <= 0;  //67 / 234 = 0
    16'b01000011_11101011 : OUT <= 0;  //67 / 235 = 0
    16'b01000011_11101100 : OUT <= 0;  //67 / 236 = 0
    16'b01000011_11101101 : OUT <= 0;  //67 / 237 = 0
    16'b01000011_11101110 : OUT <= 0;  //67 / 238 = 0
    16'b01000011_11101111 : OUT <= 0;  //67 / 239 = 0
    16'b01000011_11110000 : OUT <= 0;  //67 / 240 = 0
    16'b01000011_11110001 : OUT <= 0;  //67 / 241 = 0
    16'b01000011_11110010 : OUT <= 0;  //67 / 242 = 0
    16'b01000011_11110011 : OUT <= 0;  //67 / 243 = 0
    16'b01000011_11110100 : OUT <= 0;  //67 / 244 = 0
    16'b01000011_11110101 : OUT <= 0;  //67 / 245 = 0
    16'b01000011_11110110 : OUT <= 0;  //67 / 246 = 0
    16'b01000011_11110111 : OUT <= 0;  //67 / 247 = 0
    16'b01000011_11111000 : OUT <= 0;  //67 / 248 = 0
    16'b01000011_11111001 : OUT <= 0;  //67 / 249 = 0
    16'b01000011_11111010 : OUT <= 0;  //67 / 250 = 0
    16'b01000011_11111011 : OUT <= 0;  //67 / 251 = 0
    16'b01000011_11111100 : OUT <= 0;  //67 / 252 = 0
    16'b01000011_11111101 : OUT <= 0;  //67 / 253 = 0
    16'b01000011_11111110 : OUT <= 0;  //67 / 254 = 0
    16'b01000011_11111111 : OUT <= 0;  //67 / 255 = 0
    16'b01000100_00000000 : OUT <= 0;  //68 / 0 = 0
    16'b01000100_00000001 : OUT <= 68;  //68 / 1 = 68
    16'b01000100_00000010 : OUT <= 34;  //68 / 2 = 34
    16'b01000100_00000011 : OUT <= 22;  //68 / 3 = 22
    16'b01000100_00000100 : OUT <= 17;  //68 / 4 = 17
    16'b01000100_00000101 : OUT <= 13;  //68 / 5 = 13
    16'b01000100_00000110 : OUT <= 11;  //68 / 6 = 11
    16'b01000100_00000111 : OUT <= 9;  //68 / 7 = 9
    16'b01000100_00001000 : OUT <= 8;  //68 / 8 = 8
    16'b01000100_00001001 : OUT <= 7;  //68 / 9 = 7
    16'b01000100_00001010 : OUT <= 6;  //68 / 10 = 6
    16'b01000100_00001011 : OUT <= 6;  //68 / 11 = 6
    16'b01000100_00001100 : OUT <= 5;  //68 / 12 = 5
    16'b01000100_00001101 : OUT <= 5;  //68 / 13 = 5
    16'b01000100_00001110 : OUT <= 4;  //68 / 14 = 4
    16'b01000100_00001111 : OUT <= 4;  //68 / 15 = 4
    16'b01000100_00010000 : OUT <= 4;  //68 / 16 = 4
    16'b01000100_00010001 : OUT <= 4;  //68 / 17 = 4
    16'b01000100_00010010 : OUT <= 3;  //68 / 18 = 3
    16'b01000100_00010011 : OUT <= 3;  //68 / 19 = 3
    16'b01000100_00010100 : OUT <= 3;  //68 / 20 = 3
    16'b01000100_00010101 : OUT <= 3;  //68 / 21 = 3
    16'b01000100_00010110 : OUT <= 3;  //68 / 22 = 3
    16'b01000100_00010111 : OUT <= 2;  //68 / 23 = 2
    16'b01000100_00011000 : OUT <= 2;  //68 / 24 = 2
    16'b01000100_00011001 : OUT <= 2;  //68 / 25 = 2
    16'b01000100_00011010 : OUT <= 2;  //68 / 26 = 2
    16'b01000100_00011011 : OUT <= 2;  //68 / 27 = 2
    16'b01000100_00011100 : OUT <= 2;  //68 / 28 = 2
    16'b01000100_00011101 : OUT <= 2;  //68 / 29 = 2
    16'b01000100_00011110 : OUT <= 2;  //68 / 30 = 2
    16'b01000100_00011111 : OUT <= 2;  //68 / 31 = 2
    16'b01000100_00100000 : OUT <= 2;  //68 / 32 = 2
    16'b01000100_00100001 : OUT <= 2;  //68 / 33 = 2
    16'b01000100_00100010 : OUT <= 2;  //68 / 34 = 2
    16'b01000100_00100011 : OUT <= 1;  //68 / 35 = 1
    16'b01000100_00100100 : OUT <= 1;  //68 / 36 = 1
    16'b01000100_00100101 : OUT <= 1;  //68 / 37 = 1
    16'b01000100_00100110 : OUT <= 1;  //68 / 38 = 1
    16'b01000100_00100111 : OUT <= 1;  //68 / 39 = 1
    16'b01000100_00101000 : OUT <= 1;  //68 / 40 = 1
    16'b01000100_00101001 : OUT <= 1;  //68 / 41 = 1
    16'b01000100_00101010 : OUT <= 1;  //68 / 42 = 1
    16'b01000100_00101011 : OUT <= 1;  //68 / 43 = 1
    16'b01000100_00101100 : OUT <= 1;  //68 / 44 = 1
    16'b01000100_00101101 : OUT <= 1;  //68 / 45 = 1
    16'b01000100_00101110 : OUT <= 1;  //68 / 46 = 1
    16'b01000100_00101111 : OUT <= 1;  //68 / 47 = 1
    16'b01000100_00110000 : OUT <= 1;  //68 / 48 = 1
    16'b01000100_00110001 : OUT <= 1;  //68 / 49 = 1
    16'b01000100_00110010 : OUT <= 1;  //68 / 50 = 1
    16'b01000100_00110011 : OUT <= 1;  //68 / 51 = 1
    16'b01000100_00110100 : OUT <= 1;  //68 / 52 = 1
    16'b01000100_00110101 : OUT <= 1;  //68 / 53 = 1
    16'b01000100_00110110 : OUT <= 1;  //68 / 54 = 1
    16'b01000100_00110111 : OUT <= 1;  //68 / 55 = 1
    16'b01000100_00111000 : OUT <= 1;  //68 / 56 = 1
    16'b01000100_00111001 : OUT <= 1;  //68 / 57 = 1
    16'b01000100_00111010 : OUT <= 1;  //68 / 58 = 1
    16'b01000100_00111011 : OUT <= 1;  //68 / 59 = 1
    16'b01000100_00111100 : OUT <= 1;  //68 / 60 = 1
    16'b01000100_00111101 : OUT <= 1;  //68 / 61 = 1
    16'b01000100_00111110 : OUT <= 1;  //68 / 62 = 1
    16'b01000100_00111111 : OUT <= 1;  //68 / 63 = 1
    16'b01000100_01000000 : OUT <= 1;  //68 / 64 = 1
    16'b01000100_01000001 : OUT <= 1;  //68 / 65 = 1
    16'b01000100_01000010 : OUT <= 1;  //68 / 66 = 1
    16'b01000100_01000011 : OUT <= 1;  //68 / 67 = 1
    16'b01000100_01000100 : OUT <= 1;  //68 / 68 = 1
    16'b01000100_01000101 : OUT <= 0;  //68 / 69 = 0
    16'b01000100_01000110 : OUT <= 0;  //68 / 70 = 0
    16'b01000100_01000111 : OUT <= 0;  //68 / 71 = 0
    16'b01000100_01001000 : OUT <= 0;  //68 / 72 = 0
    16'b01000100_01001001 : OUT <= 0;  //68 / 73 = 0
    16'b01000100_01001010 : OUT <= 0;  //68 / 74 = 0
    16'b01000100_01001011 : OUT <= 0;  //68 / 75 = 0
    16'b01000100_01001100 : OUT <= 0;  //68 / 76 = 0
    16'b01000100_01001101 : OUT <= 0;  //68 / 77 = 0
    16'b01000100_01001110 : OUT <= 0;  //68 / 78 = 0
    16'b01000100_01001111 : OUT <= 0;  //68 / 79 = 0
    16'b01000100_01010000 : OUT <= 0;  //68 / 80 = 0
    16'b01000100_01010001 : OUT <= 0;  //68 / 81 = 0
    16'b01000100_01010010 : OUT <= 0;  //68 / 82 = 0
    16'b01000100_01010011 : OUT <= 0;  //68 / 83 = 0
    16'b01000100_01010100 : OUT <= 0;  //68 / 84 = 0
    16'b01000100_01010101 : OUT <= 0;  //68 / 85 = 0
    16'b01000100_01010110 : OUT <= 0;  //68 / 86 = 0
    16'b01000100_01010111 : OUT <= 0;  //68 / 87 = 0
    16'b01000100_01011000 : OUT <= 0;  //68 / 88 = 0
    16'b01000100_01011001 : OUT <= 0;  //68 / 89 = 0
    16'b01000100_01011010 : OUT <= 0;  //68 / 90 = 0
    16'b01000100_01011011 : OUT <= 0;  //68 / 91 = 0
    16'b01000100_01011100 : OUT <= 0;  //68 / 92 = 0
    16'b01000100_01011101 : OUT <= 0;  //68 / 93 = 0
    16'b01000100_01011110 : OUT <= 0;  //68 / 94 = 0
    16'b01000100_01011111 : OUT <= 0;  //68 / 95 = 0
    16'b01000100_01100000 : OUT <= 0;  //68 / 96 = 0
    16'b01000100_01100001 : OUT <= 0;  //68 / 97 = 0
    16'b01000100_01100010 : OUT <= 0;  //68 / 98 = 0
    16'b01000100_01100011 : OUT <= 0;  //68 / 99 = 0
    16'b01000100_01100100 : OUT <= 0;  //68 / 100 = 0
    16'b01000100_01100101 : OUT <= 0;  //68 / 101 = 0
    16'b01000100_01100110 : OUT <= 0;  //68 / 102 = 0
    16'b01000100_01100111 : OUT <= 0;  //68 / 103 = 0
    16'b01000100_01101000 : OUT <= 0;  //68 / 104 = 0
    16'b01000100_01101001 : OUT <= 0;  //68 / 105 = 0
    16'b01000100_01101010 : OUT <= 0;  //68 / 106 = 0
    16'b01000100_01101011 : OUT <= 0;  //68 / 107 = 0
    16'b01000100_01101100 : OUT <= 0;  //68 / 108 = 0
    16'b01000100_01101101 : OUT <= 0;  //68 / 109 = 0
    16'b01000100_01101110 : OUT <= 0;  //68 / 110 = 0
    16'b01000100_01101111 : OUT <= 0;  //68 / 111 = 0
    16'b01000100_01110000 : OUT <= 0;  //68 / 112 = 0
    16'b01000100_01110001 : OUT <= 0;  //68 / 113 = 0
    16'b01000100_01110010 : OUT <= 0;  //68 / 114 = 0
    16'b01000100_01110011 : OUT <= 0;  //68 / 115 = 0
    16'b01000100_01110100 : OUT <= 0;  //68 / 116 = 0
    16'b01000100_01110101 : OUT <= 0;  //68 / 117 = 0
    16'b01000100_01110110 : OUT <= 0;  //68 / 118 = 0
    16'b01000100_01110111 : OUT <= 0;  //68 / 119 = 0
    16'b01000100_01111000 : OUT <= 0;  //68 / 120 = 0
    16'b01000100_01111001 : OUT <= 0;  //68 / 121 = 0
    16'b01000100_01111010 : OUT <= 0;  //68 / 122 = 0
    16'b01000100_01111011 : OUT <= 0;  //68 / 123 = 0
    16'b01000100_01111100 : OUT <= 0;  //68 / 124 = 0
    16'b01000100_01111101 : OUT <= 0;  //68 / 125 = 0
    16'b01000100_01111110 : OUT <= 0;  //68 / 126 = 0
    16'b01000100_01111111 : OUT <= 0;  //68 / 127 = 0
    16'b01000100_10000000 : OUT <= 0;  //68 / 128 = 0
    16'b01000100_10000001 : OUT <= 0;  //68 / 129 = 0
    16'b01000100_10000010 : OUT <= 0;  //68 / 130 = 0
    16'b01000100_10000011 : OUT <= 0;  //68 / 131 = 0
    16'b01000100_10000100 : OUT <= 0;  //68 / 132 = 0
    16'b01000100_10000101 : OUT <= 0;  //68 / 133 = 0
    16'b01000100_10000110 : OUT <= 0;  //68 / 134 = 0
    16'b01000100_10000111 : OUT <= 0;  //68 / 135 = 0
    16'b01000100_10001000 : OUT <= 0;  //68 / 136 = 0
    16'b01000100_10001001 : OUT <= 0;  //68 / 137 = 0
    16'b01000100_10001010 : OUT <= 0;  //68 / 138 = 0
    16'b01000100_10001011 : OUT <= 0;  //68 / 139 = 0
    16'b01000100_10001100 : OUT <= 0;  //68 / 140 = 0
    16'b01000100_10001101 : OUT <= 0;  //68 / 141 = 0
    16'b01000100_10001110 : OUT <= 0;  //68 / 142 = 0
    16'b01000100_10001111 : OUT <= 0;  //68 / 143 = 0
    16'b01000100_10010000 : OUT <= 0;  //68 / 144 = 0
    16'b01000100_10010001 : OUT <= 0;  //68 / 145 = 0
    16'b01000100_10010010 : OUT <= 0;  //68 / 146 = 0
    16'b01000100_10010011 : OUT <= 0;  //68 / 147 = 0
    16'b01000100_10010100 : OUT <= 0;  //68 / 148 = 0
    16'b01000100_10010101 : OUT <= 0;  //68 / 149 = 0
    16'b01000100_10010110 : OUT <= 0;  //68 / 150 = 0
    16'b01000100_10010111 : OUT <= 0;  //68 / 151 = 0
    16'b01000100_10011000 : OUT <= 0;  //68 / 152 = 0
    16'b01000100_10011001 : OUT <= 0;  //68 / 153 = 0
    16'b01000100_10011010 : OUT <= 0;  //68 / 154 = 0
    16'b01000100_10011011 : OUT <= 0;  //68 / 155 = 0
    16'b01000100_10011100 : OUT <= 0;  //68 / 156 = 0
    16'b01000100_10011101 : OUT <= 0;  //68 / 157 = 0
    16'b01000100_10011110 : OUT <= 0;  //68 / 158 = 0
    16'b01000100_10011111 : OUT <= 0;  //68 / 159 = 0
    16'b01000100_10100000 : OUT <= 0;  //68 / 160 = 0
    16'b01000100_10100001 : OUT <= 0;  //68 / 161 = 0
    16'b01000100_10100010 : OUT <= 0;  //68 / 162 = 0
    16'b01000100_10100011 : OUT <= 0;  //68 / 163 = 0
    16'b01000100_10100100 : OUT <= 0;  //68 / 164 = 0
    16'b01000100_10100101 : OUT <= 0;  //68 / 165 = 0
    16'b01000100_10100110 : OUT <= 0;  //68 / 166 = 0
    16'b01000100_10100111 : OUT <= 0;  //68 / 167 = 0
    16'b01000100_10101000 : OUT <= 0;  //68 / 168 = 0
    16'b01000100_10101001 : OUT <= 0;  //68 / 169 = 0
    16'b01000100_10101010 : OUT <= 0;  //68 / 170 = 0
    16'b01000100_10101011 : OUT <= 0;  //68 / 171 = 0
    16'b01000100_10101100 : OUT <= 0;  //68 / 172 = 0
    16'b01000100_10101101 : OUT <= 0;  //68 / 173 = 0
    16'b01000100_10101110 : OUT <= 0;  //68 / 174 = 0
    16'b01000100_10101111 : OUT <= 0;  //68 / 175 = 0
    16'b01000100_10110000 : OUT <= 0;  //68 / 176 = 0
    16'b01000100_10110001 : OUT <= 0;  //68 / 177 = 0
    16'b01000100_10110010 : OUT <= 0;  //68 / 178 = 0
    16'b01000100_10110011 : OUT <= 0;  //68 / 179 = 0
    16'b01000100_10110100 : OUT <= 0;  //68 / 180 = 0
    16'b01000100_10110101 : OUT <= 0;  //68 / 181 = 0
    16'b01000100_10110110 : OUT <= 0;  //68 / 182 = 0
    16'b01000100_10110111 : OUT <= 0;  //68 / 183 = 0
    16'b01000100_10111000 : OUT <= 0;  //68 / 184 = 0
    16'b01000100_10111001 : OUT <= 0;  //68 / 185 = 0
    16'b01000100_10111010 : OUT <= 0;  //68 / 186 = 0
    16'b01000100_10111011 : OUT <= 0;  //68 / 187 = 0
    16'b01000100_10111100 : OUT <= 0;  //68 / 188 = 0
    16'b01000100_10111101 : OUT <= 0;  //68 / 189 = 0
    16'b01000100_10111110 : OUT <= 0;  //68 / 190 = 0
    16'b01000100_10111111 : OUT <= 0;  //68 / 191 = 0
    16'b01000100_11000000 : OUT <= 0;  //68 / 192 = 0
    16'b01000100_11000001 : OUT <= 0;  //68 / 193 = 0
    16'b01000100_11000010 : OUT <= 0;  //68 / 194 = 0
    16'b01000100_11000011 : OUT <= 0;  //68 / 195 = 0
    16'b01000100_11000100 : OUT <= 0;  //68 / 196 = 0
    16'b01000100_11000101 : OUT <= 0;  //68 / 197 = 0
    16'b01000100_11000110 : OUT <= 0;  //68 / 198 = 0
    16'b01000100_11000111 : OUT <= 0;  //68 / 199 = 0
    16'b01000100_11001000 : OUT <= 0;  //68 / 200 = 0
    16'b01000100_11001001 : OUT <= 0;  //68 / 201 = 0
    16'b01000100_11001010 : OUT <= 0;  //68 / 202 = 0
    16'b01000100_11001011 : OUT <= 0;  //68 / 203 = 0
    16'b01000100_11001100 : OUT <= 0;  //68 / 204 = 0
    16'b01000100_11001101 : OUT <= 0;  //68 / 205 = 0
    16'b01000100_11001110 : OUT <= 0;  //68 / 206 = 0
    16'b01000100_11001111 : OUT <= 0;  //68 / 207 = 0
    16'b01000100_11010000 : OUT <= 0;  //68 / 208 = 0
    16'b01000100_11010001 : OUT <= 0;  //68 / 209 = 0
    16'b01000100_11010010 : OUT <= 0;  //68 / 210 = 0
    16'b01000100_11010011 : OUT <= 0;  //68 / 211 = 0
    16'b01000100_11010100 : OUT <= 0;  //68 / 212 = 0
    16'b01000100_11010101 : OUT <= 0;  //68 / 213 = 0
    16'b01000100_11010110 : OUT <= 0;  //68 / 214 = 0
    16'b01000100_11010111 : OUT <= 0;  //68 / 215 = 0
    16'b01000100_11011000 : OUT <= 0;  //68 / 216 = 0
    16'b01000100_11011001 : OUT <= 0;  //68 / 217 = 0
    16'b01000100_11011010 : OUT <= 0;  //68 / 218 = 0
    16'b01000100_11011011 : OUT <= 0;  //68 / 219 = 0
    16'b01000100_11011100 : OUT <= 0;  //68 / 220 = 0
    16'b01000100_11011101 : OUT <= 0;  //68 / 221 = 0
    16'b01000100_11011110 : OUT <= 0;  //68 / 222 = 0
    16'b01000100_11011111 : OUT <= 0;  //68 / 223 = 0
    16'b01000100_11100000 : OUT <= 0;  //68 / 224 = 0
    16'b01000100_11100001 : OUT <= 0;  //68 / 225 = 0
    16'b01000100_11100010 : OUT <= 0;  //68 / 226 = 0
    16'b01000100_11100011 : OUT <= 0;  //68 / 227 = 0
    16'b01000100_11100100 : OUT <= 0;  //68 / 228 = 0
    16'b01000100_11100101 : OUT <= 0;  //68 / 229 = 0
    16'b01000100_11100110 : OUT <= 0;  //68 / 230 = 0
    16'b01000100_11100111 : OUT <= 0;  //68 / 231 = 0
    16'b01000100_11101000 : OUT <= 0;  //68 / 232 = 0
    16'b01000100_11101001 : OUT <= 0;  //68 / 233 = 0
    16'b01000100_11101010 : OUT <= 0;  //68 / 234 = 0
    16'b01000100_11101011 : OUT <= 0;  //68 / 235 = 0
    16'b01000100_11101100 : OUT <= 0;  //68 / 236 = 0
    16'b01000100_11101101 : OUT <= 0;  //68 / 237 = 0
    16'b01000100_11101110 : OUT <= 0;  //68 / 238 = 0
    16'b01000100_11101111 : OUT <= 0;  //68 / 239 = 0
    16'b01000100_11110000 : OUT <= 0;  //68 / 240 = 0
    16'b01000100_11110001 : OUT <= 0;  //68 / 241 = 0
    16'b01000100_11110010 : OUT <= 0;  //68 / 242 = 0
    16'b01000100_11110011 : OUT <= 0;  //68 / 243 = 0
    16'b01000100_11110100 : OUT <= 0;  //68 / 244 = 0
    16'b01000100_11110101 : OUT <= 0;  //68 / 245 = 0
    16'b01000100_11110110 : OUT <= 0;  //68 / 246 = 0
    16'b01000100_11110111 : OUT <= 0;  //68 / 247 = 0
    16'b01000100_11111000 : OUT <= 0;  //68 / 248 = 0
    16'b01000100_11111001 : OUT <= 0;  //68 / 249 = 0
    16'b01000100_11111010 : OUT <= 0;  //68 / 250 = 0
    16'b01000100_11111011 : OUT <= 0;  //68 / 251 = 0
    16'b01000100_11111100 : OUT <= 0;  //68 / 252 = 0
    16'b01000100_11111101 : OUT <= 0;  //68 / 253 = 0
    16'b01000100_11111110 : OUT <= 0;  //68 / 254 = 0
    16'b01000100_11111111 : OUT <= 0;  //68 / 255 = 0
    16'b01000101_00000000 : OUT <= 0;  //69 / 0 = 0
    16'b01000101_00000001 : OUT <= 69;  //69 / 1 = 69
    16'b01000101_00000010 : OUT <= 34;  //69 / 2 = 34
    16'b01000101_00000011 : OUT <= 23;  //69 / 3 = 23
    16'b01000101_00000100 : OUT <= 17;  //69 / 4 = 17
    16'b01000101_00000101 : OUT <= 13;  //69 / 5 = 13
    16'b01000101_00000110 : OUT <= 11;  //69 / 6 = 11
    16'b01000101_00000111 : OUT <= 9;  //69 / 7 = 9
    16'b01000101_00001000 : OUT <= 8;  //69 / 8 = 8
    16'b01000101_00001001 : OUT <= 7;  //69 / 9 = 7
    16'b01000101_00001010 : OUT <= 6;  //69 / 10 = 6
    16'b01000101_00001011 : OUT <= 6;  //69 / 11 = 6
    16'b01000101_00001100 : OUT <= 5;  //69 / 12 = 5
    16'b01000101_00001101 : OUT <= 5;  //69 / 13 = 5
    16'b01000101_00001110 : OUT <= 4;  //69 / 14 = 4
    16'b01000101_00001111 : OUT <= 4;  //69 / 15 = 4
    16'b01000101_00010000 : OUT <= 4;  //69 / 16 = 4
    16'b01000101_00010001 : OUT <= 4;  //69 / 17 = 4
    16'b01000101_00010010 : OUT <= 3;  //69 / 18 = 3
    16'b01000101_00010011 : OUT <= 3;  //69 / 19 = 3
    16'b01000101_00010100 : OUT <= 3;  //69 / 20 = 3
    16'b01000101_00010101 : OUT <= 3;  //69 / 21 = 3
    16'b01000101_00010110 : OUT <= 3;  //69 / 22 = 3
    16'b01000101_00010111 : OUT <= 3;  //69 / 23 = 3
    16'b01000101_00011000 : OUT <= 2;  //69 / 24 = 2
    16'b01000101_00011001 : OUT <= 2;  //69 / 25 = 2
    16'b01000101_00011010 : OUT <= 2;  //69 / 26 = 2
    16'b01000101_00011011 : OUT <= 2;  //69 / 27 = 2
    16'b01000101_00011100 : OUT <= 2;  //69 / 28 = 2
    16'b01000101_00011101 : OUT <= 2;  //69 / 29 = 2
    16'b01000101_00011110 : OUT <= 2;  //69 / 30 = 2
    16'b01000101_00011111 : OUT <= 2;  //69 / 31 = 2
    16'b01000101_00100000 : OUT <= 2;  //69 / 32 = 2
    16'b01000101_00100001 : OUT <= 2;  //69 / 33 = 2
    16'b01000101_00100010 : OUT <= 2;  //69 / 34 = 2
    16'b01000101_00100011 : OUT <= 1;  //69 / 35 = 1
    16'b01000101_00100100 : OUT <= 1;  //69 / 36 = 1
    16'b01000101_00100101 : OUT <= 1;  //69 / 37 = 1
    16'b01000101_00100110 : OUT <= 1;  //69 / 38 = 1
    16'b01000101_00100111 : OUT <= 1;  //69 / 39 = 1
    16'b01000101_00101000 : OUT <= 1;  //69 / 40 = 1
    16'b01000101_00101001 : OUT <= 1;  //69 / 41 = 1
    16'b01000101_00101010 : OUT <= 1;  //69 / 42 = 1
    16'b01000101_00101011 : OUT <= 1;  //69 / 43 = 1
    16'b01000101_00101100 : OUT <= 1;  //69 / 44 = 1
    16'b01000101_00101101 : OUT <= 1;  //69 / 45 = 1
    16'b01000101_00101110 : OUT <= 1;  //69 / 46 = 1
    16'b01000101_00101111 : OUT <= 1;  //69 / 47 = 1
    16'b01000101_00110000 : OUT <= 1;  //69 / 48 = 1
    16'b01000101_00110001 : OUT <= 1;  //69 / 49 = 1
    16'b01000101_00110010 : OUT <= 1;  //69 / 50 = 1
    16'b01000101_00110011 : OUT <= 1;  //69 / 51 = 1
    16'b01000101_00110100 : OUT <= 1;  //69 / 52 = 1
    16'b01000101_00110101 : OUT <= 1;  //69 / 53 = 1
    16'b01000101_00110110 : OUT <= 1;  //69 / 54 = 1
    16'b01000101_00110111 : OUT <= 1;  //69 / 55 = 1
    16'b01000101_00111000 : OUT <= 1;  //69 / 56 = 1
    16'b01000101_00111001 : OUT <= 1;  //69 / 57 = 1
    16'b01000101_00111010 : OUT <= 1;  //69 / 58 = 1
    16'b01000101_00111011 : OUT <= 1;  //69 / 59 = 1
    16'b01000101_00111100 : OUT <= 1;  //69 / 60 = 1
    16'b01000101_00111101 : OUT <= 1;  //69 / 61 = 1
    16'b01000101_00111110 : OUT <= 1;  //69 / 62 = 1
    16'b01000101_00111111 : OUT <= 1;  //69 / 63 = 1
    16'b01000101_01000000 : OUT <= 1;  //69 / 64 = 1
    16'b01000101_01000001 : OUT <= 1;  //69 / 65 = 1
    16'b01000101_01000010 : OUT <= 1;  //69 / 66 = 1
    16'b01000101_01000011 : OUT <= 1;  //69 / 67 = 1
    16'b01000101_01000100 : OUT <= 1;  //69 / 68 = 1
    16'b01000101_01000101 : OUT <= 1;  //69 / 69 = 1
    16'b01000101_01000110 : OUT <= 0;  //69 / 70 = 0
    16'b01000101_01000111 : OUT <= 0;  //69 / 71 = 0
    16'b01000101_01001000 : OUT <= 0;  //69 / 72 = 0
    16'b01000101_01001001 : OUT <= 0;  //69 / 73 = 0
    16'b01000101_01001010 : OUT <= 0;  //69 / 74 = 0
    16'b01000101_01001011 : OUT <= 0;  //69 / 75 = 0
    16'b01000101_01001100 : OUT <= 0;  //69 / 76 = 0
    16'b01000101_01001101 : OUT <= 0;  //69 / 77 = 0
    16'b01000101_01001110 : OUT <= 0;  //69 / 78 = 0
    16'b01000101_01001111 : OUT <= 0;  //69 / 79 = 0
    16'b01000101_01010000 : OUT <= 0;  //69 / 80 = 0
    16'b01000101_01010001 : OUT <= 0;  //69 / 81 = 0
    16'b01000101_01010010 : OUT <= 0;  //69 / 82 = 0
    16'b01000101_01010011 : OUT <= 0;  //69 / 83 = 0
    16'b01000101_01010100 : OUT <= 0;  //69 / 84 = 0
    16'b01000101_01010101 : OUT <= 0;  //69 / 85 = 0
    16'b01000101_01010110 : OUT <= 0;  //69 / 86 = 0
    16'b01000101_01010111 : OUT <= 0;  //69 / 87 = 0
    16'b01000101_01011000 : OUT <= 0;  //69 / 88 = 0
    16'b01000101_01011001 : OUT <= 0;  //69 / 89 = 0
    16'b01000101_01011010 : OUT <= 0;  //69 / 90 = 0
    16'b01000101_01011011 : OUT <= 0;  //69 / 91 = 0
    16'b01000101_01011100 : OUT <= 0;  //69 / 92 = 0
    16'b01000101_01011101 : OUT <= 0;  //69 / 93 = 0
    16'b01000101_01011110 : OUT <= 0;  //69 / 94 = 0
    16'b01000101_01011111 : OUT <= 0;  //69 / 95 = 0
    16'b01000101_01100000 : OUT <= 0;  //69 / 96 = 0
    16'b01000101_01100001 : OUT <= 0;  //69 / 97 = 0
    16'b01000101_01100010 : OUT <= 0;  //69 / 98 = 0
    16'b01000101_01100011 : OUT <= 0;  //69 / 99 = 0
    16'b01000101_01100100 : OUT <= 0;  //69 / 100 = 0
    16'b01000101_01100101 : OUT <= 0;  //69 / 101 = 0
    16'b01000101_01100110 : OUT <= 0;  //69 / 102 = 0
    16'b01000101_01100111 : OUT <= 0;  //69 / 103 = 0
    16'b01000101_01101000 : OUT <= 0;  //69 / 104 = 0
    16'b01000101_01101001 : OUT <= 0;  //69 / 105 = 0
    16'b01000101_01101010 : OUT <= 0;  //69 / 106 = 0
    16'b01000101_01101011 : OUT <= 0;  //69 / 107 = 0
    16'b01000101_01101100 : OUT <= 0;  //69 / 108 = 0
    16'b01000101_01101101 : OUT <= 0;  //69 / 109 = 0
    16'b01000101_01101110 : OUT <= 0;  //69 / 110 = 0
    16'b01000101_01101111 : OUT <= 0;  //69 / 111 = 0
    16'b01000101_01110000 : OUT <= 0;  //69 / 112 = 0
    16'b01000101_01110001 : OUT <= 0;  //69 / 113 = 0
    16'b01000101_01110010 : OUT <= 0;  //69 / 114 = 0
    16'b01000101_01110011 : OUT <= 0;  //69 / 115 = 0
    16'b01000101_01110100 : OUT <= 0;  //69 / 116 = 0
    16'b01000101_01110101 : OUT <= 0;  //69 / 117 = 0
    16'b01000101_01110110 : OUT <= 0;  //69 / 118 = 0
    16'b01000101_01110111 : OUT <= 0;  //69 / 119 = 0
    16'b01000101_01111000 : OUT <= 0;  //69 / 120 = 0
    16'b01000101_01111001 : OUT <= 0;  //69 / 121 = 0
    16'b01000101_01111010 : OUT <= 0;  //69 / 122 = 0
    16'b01000101_01111011 : OUT <= 0;  //69 / 123 = 0
    16'b01000101_01111100 : OUT <= 0;  //69 / 124 = 0
    16'b01000101_01111101 : OUT <= 0;  //69 / 125 = 0
    16'b01000101_01111110 : OUT <= 0;  //69 / 126 = 0
    16'b01000101_01111111 : OUT <= 0;  //69 / 127 = 0
    16'b01000101_10000000 : OUT <= 0;  //69 / 128 = 0
    16'b01000101_10000001 : OUT <= 0;  //69 / 129 = 0
    16'b01000101_10000010 : OUT <= 0;  //69 / 130 = 0
    16'b01000101_10000011 : OUT <= 0;  //69 / 131 = 0
    16'b01000101_10000100 : OUT <= 0;  //69 / 132 = 0
    16'b01000101_10000101 : OUT <= 0;  //69 / 133 = 0
    16'b01000101_10000110 : OUT <= 0;  //69 / 134 = 0
    16'b01000101_10000111 : OUT <= 0;  //69 / 135 = 0
    16'b01000101_10001000 : OUT <= 0;  //69 / 136 = 0
    16'b01000101_10001001 : OUT <= 0;  //69 / 137 = 0
    16'b01000101_10001010 : OUT <= 0;  //69 / 138 = 0
    16'b01000101_10001011 : OUT <= 0;  //69 / 139 = 0
    16'b01000101_10001100 : OUT <= 0;  //69 / 140 = 0
    16'b01000101_10001101 : OUT <= 0;  //69 / 141 = 0
    16'b01000101_10001110 : OUT <= 0;  //69 / 142 = 0
    16'b01000101_10001111 : OUT <= 0;  //69 / 143 = 0
    16'b01000101_10010000 : OUT <= 0;  //69 / 144 = 0
    16'b01000101_10010001 : OUT <= 0;  //69 / 145 = 0
    16'b01000101_10010010 : OUT <= 0;  //69 / 146 = 0
    16'b01000101_10010011 : OUT <= 0;  //69 / 147 = 0
    16'b01000101_10010100 : OUT <= 0;  //69 / 148 = 0
    16'b01000101_10010101 : OUT <= 0;  //69 / 149 = 0
    16'b01000101_10010110 : OUT <= 0;  //69 / 150 = 0
    16'b01000101_10010111 : OUT <= 0;  //69 / 151 = 0
    16'b01000101_10011000 : OUT <= 0;  //69 / 152 = 0
    16'b01000101_10011001 : OUT <= 0;  //69 / 153 = 0
    16'b01000101_10011010 : OUT <= 0;  //69 / 154 = 0
    16'b01000101_10011011 : OUT <= 0;  //69 / 155 = 0
    16'b01000101_10011100 : OUT <= 0;  //69 / 156 = 0
    16'b01000101_10011101 : OUT <= 0;  //69 / 157 = 0
    16'b01000101_10011110 : OUT <= 0;  //69 / 158 = 0
    16'b01000101_10011111 : OUT <= 0;  //69 / 159 = 0
    16'b01000101_10100000 : OUT <= 0;  //69 / 160 = 0
    16'b01000101_10100001 : OUT <= 0;  //69 / 161 = 0
    16'b01000101_10100010 : OUT <= 0;  //69 / 162 = 0
    16'b01000101_10100011 : OUT <= 0;  //69 / 163 = 0
    16'b01000101_10100100 : OUT <= 0;  //69 / 164 = 0
    16'b01000101_10100101 : OUT <= 0;  //69 / 165 = 0
    16'b01000101_10100110 : OUT <= 0;  //69 / 166 = 0
    16'b01000101_10100111 : OUT <= 0;  //69 / 167 = 0
    16'b01000101_10101000 : OUT <= 0;  //69 / 168 = 0
    16'b01000101_10101001 : OUT <= 0;  //69 / 169 = 0
    16'b01000101_10101010 : OUT <= 0;  //69 / 170 = 0
    16'b01000101_10101011 : OUT <= 0;  //69 / 171 = 0
    16'b01000101_10101100 : OUT <= 0;  //69 / 172 = 0
    16'b01000101_10101101 : OUT <= 0;  //69 / 173 = 0
    16'b01000101_10101110 : OUT <= 0;  //69 / 174 = 0
    16'b01000101_10101111 : OUT <= 0;  //69 / 175 = 0
    16'b01000101_10110000 : OUT <= 0;  //69 / 176 = 0
    16'b01000101_10110001 : OUT <= 0;  //69 / 177 = 0
    16'b01000101_10110010 : OUT <= 0;  //69 / 178 = 0
    16'b01000101_10110011 : OUT <= 0;  //69 / 179 = 0
    16'b01000101_10110100 : OUT <= 0;  //69 / 180 = 0
    16'b01000101_10110101 : OUT <= 0;  //69 / 181 = 0
    16'b01000101_10110110 : OUT <= 0;  //69 / 182 = 0
    16'b01000101_10110111 : OUT <= 0;  //69 / 183 = 0
    16'b01000101_10111000 : OUT <= 0;  //69 / 184 = 0
    16'b01000101_10111001 : OUT <= 0;  //69 / 185 = 0
    16'b01000101_10111010 : OUT <= 0;  //69 / 186 = 0
    16'b01000101_10111011 : OUT <= 0;  //69 / 187 = 0
    16'b01000101_10111100 : OUT <= 0;  //69 / 188 = 0
    16'b01000101_10111101 : OUT <= 0;  //69 / 189 = 0
    16'b01000101_10111110 : OUT <= 0;  //69 / 190 = 0
    16'b01000101_10111111 : OUT <= 0;  //69 / 191 = 0
    16'b01000101_11000000 : OUT <= 0;  //69 / 192 = 0
    16'b01000101_11000001 : OUT <= 0;  //69 / 193 = 0
    16'b01000101_11000010 : OUT <= 0;  //69 / 194 = 0
    16'b01000101_11000011 : OUT <= 0;  //69 / 195 = 0
    16'b01000101_11000100 : OUT <= 0;  //69 / 196 = 0
    16'b01000101_11000101 : OUT <= 0;  //69 / 197 = 0
    16'b01000101_11000110 : OUT <= 0;  //69 / 198 = 0
    16'b01000101_11000111 : OUT <= 0;  //69 / 199 = 0
    16'b01000101_11001000 : OUT <= 0;  //69 / 200 = 0
    16'b01000101_11001001 : OUT <= 0;  //69 / 201 = 0
    16'b01000101_11001010 : OUT <= 0;  //69 / 202 = 0
    16'b01000101_11001011 : OUT <= 0;  //69 / 203 = 0
    16'b01000101_11001100 : OUT <= 0;  //69 / 204 = 0
    16'b01000101_11001101 : OUT <= 0;  //69 / 205 = 0
    16'b01000101_11001110 : OUT <= 0;  //69 / 206 = 0
    16'b01000101_11001111 : OUT <= 0;  //69 / 207 = 0
    16'b01000101_11010000 : OUT <= 0;  //69 / 208 = 0
    16'b01000101_11010001 : OUT <= 0;  //69 / 209 = 0
    16'b01000101_11010010 : OUT <= 0;  //69 / 210 = 0
    16'b01000101_11010011 : OUT <= 0;  //69 / 211 = 0
    16'b01000101_11010100 : OUT <= 0;  //69 / 212 = 0
    16'b01000101_11010101 : OUT <= 0;  //69 / 213 = 0
    16'b01000101_11010110 : OUT <= 0;  //69 / 214 = 0
    16'b01000101_11010111 : OUT <= 0;  //69 / 215 = 0
    16'b01000101_11011000 : OUT <= 0;  //69 / 216 = 0
    16'b01000101_11011001 : OUT <= 0;  //69 / 217 = 0
    16'b01000101_11011010 : OUT <= 0;  //69 / 218 = 0
    16'b01000101_11011011 : OUT <= 0;  //69 / 219 = 0
    16'b01000101_11011100 : OUT <= 0;  //69 / 220 = 0
    16'b01000101_11011101 : OUT <= 0;  //69 / 221 = 0
    16'b01000101_11011110 : OUT <= 0;  //69 / 222 = 0
    16'b01000101_11011111 : OUT <= 0;  //69 / 223 = 0
    16'b01000101_11100000 : OUT <= 0;  //69 / 224 = 0
    16'b01000101_11100001 : OUT <= 0;  //69 / 225 = 0
    16'b01000101_11100010 : OUT <= 0;  //69 / 226 = 0
    16'b01000101_11100011 : OUT <= 0;  //69 / 227 = 0
    16'b01000101_11100100 : OUT <= 0;  //69 / 228 = 0
    16'b01000101_11100101 : OUT <= 0;  //69 / 229 = 0
    16'b01000101_11100110 : OUT <= 0;  //69 / 230 = 0
    16'b01000101_11100111 : OUT <= 0;  //69 / 231 = 0
    16'b01000101_11101000 : OUT <= 0;  //69 / 232 = 0
    16'b01000101_11101001 : OUT <= 0;  //69 / 233 = 0
    16'b01000101_11101010 : OUT <= 0;  //69 / 234 = 0
    16'b01000101_11101011 : OUT <= 0;  //69 / 235 = 0
    16'b01000101_11101100 : OUT <= 0;  //69 / 236 = 0
    16'b01000101_11101101 : OUT <= 0;  //69 / 237 = 0
    16'b01000101_11101110 : OUT <= 0;  //69 / 238 = 0
    16'b01000101_11101111 : OUT <= 0;  //69 / 239 = 0
    16'b01000101_11110000 : OUT <= 0;  //69 / 240 = 0
    16'b01000101_11110001 : OUT <= 0;  //69 / 241 = 0
    16'b01000101_11110010 : OUT <= 0;  //69 / 242 = 0
    16'b01000101_11110011 : OUT <= 0;  //69 / 243 = 0
    16'b01000101_11110100 : OUT <= 0;  //69 / 244 = 0
    16'b01000101_11110101 : OUT <= 0;  //69 / 245 = 0
    16'b01000101_11110110 : OUT <= 0;  //69 / 246 = 0
    16'b01000101_11110111 : OUT <= 0;  //69 / 247 = 0
    16'b01000101_11111000 : OUT <= 0;  //69 / 248 = 0
    16'b01000101_11111001 : OUT <= 0;  //69 / 249 = 0
    16'b01000101_11111010 : OUT <= 0;  //69 / 250 = 0
    16'b01000101_11111011 : OUT <= 0;  //69 / 251 = 0
    16'b01000101_11111100 : OUT <= 0;  //69 / 252 = 0
    16'b01000101_11111101 : OUT <= 0;  //69 / 253 = 0
    16'b01000101_11111110 : OUT <= 0;  //69 / 254 = 0
    16'b01000101_11111111 : OUT <= 0;  //69 / 255 = 0
    16'b01000110_00000000 : OUT <= 0;  //70 / 0 = 0
    16'b01000110_00000001 : OUT <= 70;  //70 / 1 = 70
    16'b01000110_00000010 : OUT <= 35;  //70 / 2 = 35
    16'b01000110_00000011 : OUT <= 23;  //70 / 3 = 23
    16'b01000110_00000100 : OUT <= 17;  //70 / 4 = 17
    16'b01000110_00000101 : OUT <= 14;  //70 / 5 = 14
    16'b01000110_00000110 : OUT <= 11;  //70 / 6 = 11
    16'b01000110_00000111 : OUT <= 10;  //70 / 7 = 10
    16'b01000110_00001000 : OUT <= 8;  //70 / 8 = 8
    16'b01000110_00001001 : OUT <= 7;  //70 / 9 = 7
    16'b01000110_00001010 : OUT <= 7;  //70 / 10 = 7
    16'b01000110_00001011 : OUT <= 6;  //70 / 11 = 6
    16'b01000110_00001100 : OUT <= 5;  //70 / 12 = 5
    16'b01000110_00001101 : OUT <= 5;  //70 / 13 = 5
    16'b01000110_00001110 : OUT <= 5;  //70 / 14 = 5
    16'b01000110_00001111 : OUT <= 4;  //70 / 15 = 4
    16'b01000110_00010000 : OUT <= 4;  //70 / 16 = 4
    16'b01000110_00010001 : OUT <= 4;  //70 / 17 = 4
    16'b01000110_00010010 : OUT <= 3;  //70 / 18 = 3
    16'b01000110_00010011 : OUT <= 3;  //70 / 19 = 3
    16'b01000110_00010100 : OUT <= 3;  //70 / 20 = 3
    16'b01000110_00010101 : OUT <= 3;  //70 / 21 = 3
    16'b01000110_00010110 : OUT <= 3;  //70 / 22 = 3
    16'b01000110_00010111 : OUT <= 3;  //70 / 23 = 3
    16'b01000110_00011000 : OUT <= 2;  //70 / 24 = 2
    16'b01000110_00011001 : OUT <= 2;  //70 / 25 = 2
    16'b01000110_00011010 : OUT <= 2;  //70 / 26 = 2
    16'b01000110_00011011 : OUT <= 2;  //70 / 27 = 2
    16'b01000110_00011100 : OUT <= 2;  //70 / 28 = 2
    16'b01000110_00011101 : OUT <= 2;  //70 / 29 = 2
    16'b01000110_00011110 : OUT <= 2;  //70 / 30 = 2
    16'b01000110_00011111 : OUT <= 2;  //70 / 31 = 2
    16'b01000110_00100000 : OUT <= 2;  //70 / 32 = 2
    16'b01000110_00100001 : OUT <= 2;  //70 / 33 = 2
    16'b01000110_00100010 : OUT <= 2;  //70 / 34 = 2
    16'b01000110_00100011 : OUT <= 2;  //70 / 35 = 2
    16'b01000110_00100100 : OUT <= 1;  //70 / 36 = 1
    16'b01000110_00100101 : OUT <= 1;  //70 / 37 = 1
    16'b01000110_00100110 : OUT <= 1;  //70 / 38 = 1
    16'b01000110_00100111 : OUT <= 1;  //70 / 39 = 1
    16'b01000110_00101000 : OUT <= 1;  //70 / 40 = 1
    16'b01000110_00101001 : OUT <= 1;  //70 / 41 = 1
    16'b01000110_00101010 : OUT <= 1;  //70 / 42 = 1
    16'b01000110_00101011 : OUT <= 1;  //70 / 43 = 1
    16'b01000110_00101100 : OUT <= 1;  //70 / 44 = 1
    16'b01000110_00101101 : OUT <= 1;  //70 / 45 = 1
    16'b01000110_00101110 : OUT <= 1;  //70 / 46 = 1
    16'b01000110_00101111 : OUT <= 1;  //70 / 47 = 1
    16'b01000110_00110000 : OUT <= 1;  //70 / 48 = 1
    16'b01000110_00110001 : OUT <= 1;  //70 / 49 = 1
    16'b01000110_00110010 : OUT <= 1;  //70 / 50 = 1
    16'b01000110_00110011 : OUT <= 1;  //70 / 51 = 1
    16'b01000110_00110100 : OUT <= 1;  //70 / 52 = 1
    16'b01000110_00110101 : OUT <= 1;  //70 / 53 = 1
    16'b01000110_00110110 : OUT <= 1;  //70 / 54 = 1
    16'b01000110_00110111 : OUT <= 1;  //70 / 55 = 1
    16'b01000110_00111000 : OUT <= 1;  //70 / 56 = 1
    16'b01000110_00111001 : OUT <= 1;  //70 / 57 = 1
    16'b01000110_00111010 : OUT <= 1;  //70 / 58 = 1
    16'b01000110_00111011 : OUT <= 1;  //70 / 59 = 1
    16'b01000110_00111100 : OUT <= 1;  //70 / 60 = 1
    16'b01000110_00111101 : OUT <= 1;  //70 / 61 = 1
    16'b01000110_00111110 : OUT <= 1;  //70 / 62 = 1
    16'b01000110_00111111 : OUT <= 1;  //70 / 63 = 1
    16'b01000110_01000000 : OUT <= 1;  //70 / 64 = 1
    16'b01000110_01000001 : OUT <= 1;  //70 / 65 = 1
    16'b01000110_01000010 : OUT <= 1;  //70 / 66 = 1
    16'b01000110_01000011 : OUT <= 1;  //70 / 67 = 1
    16'b01000110_01000100 : OUT <= 1;  //70 / 68 = 1
    16'b01000110_01000101 : OUT <= 1;  //70 / 69 = 1
    16'b01000110_01000110 : OUT <= 1;  //70 / 70 = 1
    16'b01000110_01000111 : OUT <= 0;  //70 / 71 = 0
    16'b01000110_01001000 : OUT <= 0;  //70 / 72 = 0
    16'b01000110_01001001 : OUT <= 0;  //70 / 73 = 0
    16'b01000110_01001010 : OUT <= 0;  //70 / 74 = 0
    16'b01000110_01001011 : OUT <= 0;  //70 / 75 = 0
    16'b01000110_01001100 : OUT <= 0;  //70 / 76 = 0
    16'b01000110_01001101 : OUT <= 0;  //70 / 77 = 0
    16'b01000110_01001110 : OUT <= 0;  //70 / 78 = 0
    16'b01000110_01001111 : OUT <= 0;  //70 / 79 = 0
    16'b01000110_01010000 : OUT <= 0;  //70 / 80 = 0
    16'b01000110_01010001 : OUT <= 0;  //70 / 81 = 0
    16'b01000110_01010010 : OUT <= 0;  //70 / 82 = 0
    16'b01000110_01010011 : OUT <= 0;  //70 / 83 = 0
    16'b01000110_01010100 : OUT <= 0;  //70 / 84 = 0
    16'b01000110_01010101 : OUT <= 0;  //70 / 85 = 0
    16'b01000110_01010110 : OUT <= 0;  //70 / 86 = 0
    16'b01000110_01010111 : OUT <= 0;  //70 / 87 = 0
    16'b01000110_01011000 : OUT <= 0;  //70 / 88 = 0
    16'b01000110_01011001 : OUT <= 0;  //70 / 89 = 0
    16'b01000110_01011010 : OUT <= 0;  //70 / 90 = 0
    16'b01000110_01011011 : OUT <= 0;  //70 / 91 = 0
    16'b01000110_01011100 : OUT <= 0;  //70 / 92 = 0
    16'b01000110_01011101 : OUT <= 0;  //70 / 93 = 0
    16'b01000110_01011110 : OUT <= 0;  //70 / 94 = 0
    16'b01000110_01011111 : OUT <= 0;  //70 / 95 = 0
    16'b01000110_01100000 : OUT <= 0;  //70 / 96 = 0
    16'b01000110_01100001 : OUT <= 0;  //70 / 97 = 0
    16'b01000110_01100010 : OUT <= 0;  //70 / 98 = 0
    16'b01000110_01100011 : OUT <= 0;  //70 / 99 = 0
    16'b01000110_01100100 : OUT <= 0;  //70 / 100 = 0
    16'b01000110_01100101 : OUT <= 0;  //70 / 101 = 0
    16'b01000110_01100110 : OUT <= 0;  //70 / 102 = 0
    16'b01000110_01100111 : OUT <= 0;  //70 / 103 = 0
    16'b01000110_01101000 : OUT <= 0;  //70 / 104 = 0
    16'b01000110_01101001 : OUT <= 0;  //70 / 105 = 0
    16'b01000110_01101010 : OUT <= 0;  //70 / 106 = 0
    16'b01000110_01101011 : OUT <= 0;  //70 / 107 = 0
    16'b01000110_01101100 : OUT <= 0;  //70 / 108 = 0
    16'b01000110_01101101 : OUT <= 0;  //70 / 109 = 0
    16'b01000110_01101110 : OUT <= 0;  //70 / 110 = 0
    16'b01000110_01101111 : OUT <= 0;  //70 / 111 = 0
    16'b01000110_01110000 : OUT <= 0;  //70 / 112 = 0
    16'b01000110_01110001 : OUT <= 0;  //70 / 113 = 0
    16'b01000110_01110010 : OUT <= 0;  //70 / 114 = 0
    16'b01000110_01110011 : OUT <= 0;  //70 / 115 = 0
    16'b01000110_01110100 : OUT <= 0;  //70 / 116 = 0
    16'b01000110_01110101 : OUT <= 0;  //70 / 117 = 0
    16'b01000110_01110110 : OUT <= 0;  //70 / 118 = 0
    16'b01000110_01110111 : OUT <= 0;  //70 / 119 = 0
    16'b01000110_01111000 : OUT <= 0;  //70 / 120 = 0
    16'b01000110_01111001 : OUT <= 0;  //70 / 121 = 0
    16'b01000110_01111010 : OUT <= 0;  //70 / 122 = 0
    16'b01000110_01111011 : OUT <= 0;  //70 / 123 = 0
    16'b01000110_01111100 : OUT <= 0;  //70 / 124 = 0
    16'b01000110_01111101 : OUT <= 0;  //70 / 125 = 0
    16'b01000110_01111110 : OUT <= 0;  //70 / 126 = 0
    16'b01000110_01111111 : OUT <= 0;  //70 / 127 = 0
    16'b01000110_10000000 : OUT <= 0;  //70 / 128 = 0
    16'b01000110_10000001 : OUT <= 0;  //70 / 129 = 0
    16'b01000110_10000010 : OUT <= 0;  //70 / 130 = 0
    16'b01000110_10000011 : OUT <= 0;  //70 / 131 = 0
    16'b01000110_10000100 : OUT <= 0;  //70 / 132 = 0
    16'b01000110_10000101 : OUT <= 0;  //70 / 133 = 0
    16'b01000110_10000110 : OUT <= 0;  //70 / 134 = 0
    16'b01000110_10000111 : OUT <= 0;  //70 / 135 = 0
    16'b01000110_10001000 : OUT <= 0;  //70 / 136 = 0
    16'b01000110_10001001 : OUT <= 0;  //70 / 137 = 0
    16'b01000110_10001010 : OUT <= 0;  //70 / 138 = 0
    16'b01000110_10001011 : OUT <= 0;  //70 / 139 = 0
    16'b01000110_10001100 : OUT <= 0;  //70 / 140 = 0
    16'b01000110_10001101 : OUT <= 0;  //70 / 141 = 0
    16'b01000110_10001110 : OUT <= 0;  //70 / 142 = 0
    16'b01000110_10001111 : OUT <= 0;  //70 / 143 = 0
    16'b01000110_10010000 : OUT <= 0;  //70 / 144 = 0
    16'b01000110_10010001 : OUT <= 0;  //70 / 145 = 0
    16'b01000110_10010010 : OUT <= 0;  //70 / 146 = 0
    16'b01000110_10010011 : OUT <= 0;  //70 / 147 = 0
    16'b01000110_10010100 : OUT <= 0;  //70 / 148 = 0
    16'b01000110_10010101 : OUT <= 0;  //70 / 149 = 0
    16'b01000110_10010110 : OUT <= 0;  //70 / 150 = 0
    16'b01000110_10010111 : OUT <= 0;  //70 / 151 = 0
    16'b01000110_10011000 : OUT <= 0;  //70 / 152 = 0
    16'b01000110_10011001 : OUT <= 0;  //70 / 153 = 0
    16'b01000110_10011010 : OUT <= 0;  //70 / 154 = 0
    16'b01000110_10011011 : OUT <= 0;  //70 / 155 = 0
    16'b01000110_10011100 : OUT <= 0;  //70 / 156 = 0
    16'b01000110_10011101 : OUT <= 0;  //70 / 157 = 0
    16'b01000110_10011110 : OUT <= 0;  //70 / 158 = 0
    16'b01000110_10011111 : OUT <= 0;  //70 / 159 = 0
    16'b01000110_10100000 : OUT <= 0;  //70 / 160 = 0
    16'b01000110_10100001 : OUT <= 0;  //70 / 161 = 0
    16'b01000110_10100010 : OUT <= 0;  //70 / 162 = 0
    16'b01000110_10100011 : OUT <= 0;  //70 / 163 = 0
    16'b01000110_10100100 : OUT <= 0;  //70 / 164 = 0
    16'b01000110_10100101 : OUT <= 0;  //70 / 165 = 0
    16'b01000110_10100110 : OUT <= 0;  //70 / 166 = 0
    16'b01000110_10100111 : OUT <= 0;  //70 / 167 = 0
    16'b01000110_10101000 : OUT <= 0;  //70 / 168 = 0
    16'b01000110_10101001 : OUT <= 0;  //70 / 169 = 0
    16'b01000110_10101010 : OUT <= 0;  //70 / 170 = 0
    16'b01000110_10101011 : OUT <= 0;  //70 / 171 = 0
    16'b01000110_10101100 : OUT <= 0;  //70 / 172 = 0
    16'b01000110_10101101 : OUT <= 0;  //70 / 173 = 0
    16'b01000110_10101110 : OUT <= 0;  //70 / 174 = 0
    16'b01000110_10101111 : OUT <= 0;  //70 / 175 = 0
    16'b01000110_10110000 : OUT <= 0;  //70 / 176 = 0
    16'b01000110_10110001 : OUT <= 0;  //70 / 177 = 0
    16'b01000110_10110010 : OUT <= 0;  //70 / 178 = 0
    16'b01000110_10110011 : OUT <= 0;  //70 / 179 = 0
    16'b01000110_10110100 : OUT <= 0;  //70 / 180 = 0
    16'b01000110_10110101 : OUT <= 0;  //70 / 181 = 0
    16'b01000110_10110110 : OUT <= 0;  //70 / 182 = 0
    16'b01000110_10110111 : OUT <= 0;  //70 / 183 = 0
    16'b01000110_10111000 : OUT <= 0;  //70 / 184 = 0
    16'b01000110_10111001 : OUT <= 0;  //70 / 185 = 0
    16'b01000110_10111010 : OUT <= 0;  //70 / 186 = 0
    16'b01000110_10111011 : OUT <= 0;  //70 / 187 = 0
    16'b01000110_10111100 : OUT <= 0;  //70 / 188 = 0
    16'b01000110_10111101 : OUT <= 0;  //70 / 189 = 0
    16'b01000110_10111110 : OUT <= 0;  //70 / 190 = 0
    16'b01000110_10111111 : OUT <= 0;  //70 / 191 = 0
    16'b01000110_11000000 : OUT <= 0;  //70 / 192 = 0
    16'b01000110_11000001 : OUT <= 0;  //70 / 193 = 0
    16'b01000110_11000010 : OUT <= 0;  //70 / 194 = 0
    16'b01000110_11000011 : OUT <= 0;  //70 / 195 = 0
    16'b01000110_11000100 : OUT <= 0;  //70 / 196 = 0
    16'b01000110_11000101 : OUT <= 0;  //70 / 197 = 0
    16'b01000110_11000110 : OUT <= 0;  //70 / 198 = 0
    16'b01000110_11000111 : OUT <= 0;  //70 / 199 = 0
    16'b01000110_11001000 : OUT <= 0;  //70 / 200 = 0
    16'b01000110_11001001 : OUT <= 0;  //70 / 201 = 0
    16'b01000110_11001010 : OUT <= 0;  //70 / 202 = 0
    16'b01000110_11001011 : OUT <= 0;  //70 / 203 = 0
    16'b01000110_11001100 : OUT <= 0;  //70 / 204 = 0
    16'b01000110_11001101 : OUT <= 0;  //70 / 205 = 0
    16'b01000110_11001110 : OUT <= 0;  //70 / 206 = 0
    16'b01000110_11001111 : OUT <= 0;  //70 / 207 = 0
    16'b01000110_11010000 : OUT <= 0;  //70 / 208 = 0
    16'b01000110_11010001 : OUT <= 0;  //70 / 209 = 0
    16'b01000110_11010010 : OUT <= 0;  //70 / 210 = 0
    16'b01000110_11010011 : OUT <= 0;  //70 / 211 = 0
    16'b01000110_11010100 : OUT <= 0;  //70 / 212 = 0
    16'b01000110_11010101 : OUT <= 0;  //70 / 213 = 0
    16'b01000110_11010110 : OUT <= 0;  //70 / 214 = 0
    16'b01000110_11010111 : OUT <= 0;  //70 / 215 = 0
    16'b01000110_11011000 : OUT <= 0;  //70 / 216 = 0
    16'b01000110_11011001 : OUT <= 0;  //70 / 217 = 0
    16'b01000110_11011010 : OUT <= 0;  //70 / 218 = 0
    16'b01000110_11011011 : OUT <= 0;  //70 / 219 = 0
    16'b01000110_11011100 : OUT <= 0;  //70 / 220 = 0
    16'b01000110_11011101 : OUT <= 0;  //70 / 221 = 0
    16'b01000110_11011110 : OUT <= 0;  //70 / 222 = 0
    16'b01000110_11011111 : OUT <= 0;  //70 / 223 = 0
    16'b01000110_11100000 : OUT <= 0;  //70 / 224 = 0
    16'b01000110_11100001 : OUT <= 0;  //70 / 225 = 0
    16'b01000110_11100010 : OUT <= 0;  //70 / 226 = 0
    16'b01000110_11100011 : OUT <= 0;  //70 / 227 = 0
    16'b01000110_11100100 : OUT <= 0;  //70 / 228 = 0
    16'b01000110_11100101 : OUT <= 0;  //70 / 229 = 0
    16'b01000110_11100110 : OUT <= 0;  //70 / 230 = 0
    16'b01000110_11100111 : OUT <= 0;  //70 / 231 = 0
    16'b01000110_11101000 : OUT <= 0;  //70 / 232 = 0
    16'b01000110_11101001 : OUT <= 0;  //70 / 233 = 0
    16'b01000110_11101010 : OUT <= 0;  //70 / 234 = 0
    16'b01000110_11101011 : OUT <= 0;  //70 / 235 = 0
    16'b01000110_11101100 : OUT <= 0;  //70 / 236 = 0
    16'b01000110_11101101 : OUT <= 0;  //70 / 237 = 0
    16'b01000110_11101110 : OUT <= 0;  //70 / 238 = 0
    16'b01000110_11101111 : OUT <= 0;  //70 / 239 = 0
    16'b01000110_11110000 : OUT <= 0;  //70 / 240 = 0
    16'b01000110_11110001 : OUT <= 0;  //70 / 241 = 0
    16'b01000110_11110010 : OUT <= 0;  //70 / 242 = 0
    16'b01000110_11110011 : OUT <= 0;  //70 / 243 = 0
    16'b01000110_11110100 : OUT <= 0;  //70 / 244 = 0
    16'b01000110_11110101 : OUT <= 0;  //70 / 245 = 0
    16'b01000110_11110110 : OUT <= 0;  //70 / 246 = 0
    16'b01000110_11110111 : OUT <= 0;  //70 / 247 = 0
    16'b01000110_11111000 : OUT <= 0;  //70 / 248 = 0
    16'b01000110_11111001 : OUT <= 0;  //70 / 249 = 0
    16'b01000110_11111010 : OUT <= 0;  //70 / 250 = 0
    16'b01000110_11111011 : OUT <= 0;  //70 / 251 = 0
    16'b01000110_11111100 : OUT <= 0;  //70 / 252 = 0
    16'b01000110_11111101 : OUT <= 0;  //70 / 253 = 0
    16'b01000110_11111110 : OUT <= 0;  //70 / 254 = 0
    16'b01000110_11111111 : OUT <= 0;  //70 / 255 = 0
    16'b01000111_00000000 : OUT <= 0;  //71 / 0 = 0
    16'b01000111_00000001 : OUT <= 71;  //71 / 1 = 71
    16'b01000111_00000010 : OUT <= 35;  //71 / 2 = 35
    16'b01000111_00000011 : OUT <= 23;  //71 / 3 = 23
    16'b01000111_00000100 : OUT <= 17;  //71 / 4 = 17
    16'b01000111_00000101 : OUT <= 14;  //71 / 5 = 14
    16'b01000111_00000110 : OUT <= 11;  //71 / 6 = 11
    16'b01000111_00000111 : OUT <= 10;  //71 / 7 = 10
    16'b01000111_00001000 : OUT <= 8;  //71 / 8 = 8
    16'b01000111_00001001 : OUT <= 7;  //71 / 9 = 7
    16'b01000111_00001010 : OUT <= 7;  //71 / 10 = 7
    16'b01000111_00001011 : OUT <= 6;  //71 / 11 = 6
    16'b01000111_00001100 : OUT <= 5;  //71 / 12 = 5
    16'b01000111_00001101 : OUT <= 5;  //71 / 13 = 5
    16'b01000111_00001110 : OUT <= 5;  //71 / 14 = 5
    16'b01000111_00001111 : OUT <= 4;  //71 / 15 = 4
    16'b01000111_00010000 : OUT <= 4;  //71 / 16 = 4
    16'b01000111_00010001 : OUT <= 4;  //71 / 17 = 4
    16'b01000111_00010010 : OUT <= 3;  //71 / 18 = 3
    16'b01000111_00010011 : OUT <= 3;  //71 / 19 = 3
    16'b01000111_00010100 : OUT <= 3;  //71 / 20 = 3
    16'b01000111_00010101 : OUT <= 3;  //71 / 21 = 3
    16'b01000111_00010110 : OUT <= 3;  //71 / 22 = 3
    16'b01000111_00010111 : OUT <= 3;  //71 / 23 = 3
    16'b01000111_00011000 : OUT <= 2;  //71 / 24 = 2
    16'b01000111_00011001 : OUT <= 2;  //71 / 25 = 2
    16'b01000111_00011010 : OUT <= 2;  //71 / 26 = 2
    16'b01000111_00011011 : OUT <= 2;  //71 / 27 = 2
    16'b01000111_00011100 : OUT <= 2;  //71 / 28 = 2
    16'b01000111_00011101 : OUT <= 2;  //71 / 29 = 2
    16'b01000111_00011110 : OUT <= 2;  //71 / 30 = 2
    16'b01000111_00011111 : OUT <= 2;  //71 / 31 = 2
    16'b01000111_00100000 : OUT <= 2;  //71 / 32 = 2
    16'b01000111_00100001 : OUT <= 2;  //71 / 33 = 2
    16'b01000111_00100010 : OUT <= 2;  //71 / 34 = 2
    16'b01000111_00100011 : OUT <= 2;  //71 / 35 = 2
    16'b01000111_00100100 : OUT <= 1;  //71 / 36 = 1
    16'b01000111_00100101 : OUT <= 1;  //71 / 37 = 1
    16'b01000111_00100110 : OUT <= 1;  //71 / 38 = 1
    16'b01000111_00100111 : OUT <= 1;  //71 / 39 = 1
    16'b01000111_00101000 : OUT <= 1;  //71 / 40 = 1
    16'b01000111_00101001 : OUT <= 1;  //71 / 41 = 1
    16'b01000111_00101010 : OUT <= 1;  //71 / 42 = 1
    16'b01000111_00101011 : OUT <= 1;  //71 / 43 = 1
    16'b01000111_00101100 : OUT <= 1;  //71 / 44 = 1
    16'b01000111_00101101 : OUT <= 1;  //71 / 45 = 1
    16'b01000111_00101110 : OUT <= 1;  //71 / 46 = 1
    16'b01000111_00101111 : OUT <= 1;  //71 / 47 = 1
    16'b01000111_00110000 : OUT <= 1;  //71 / 48 = 1
    16'b01000111_00110001 : OUT <= 1;  //71 / 49 = 1
    16'b01000111_00110010 : OUT <= 1;  //71 / 50 = 1
    16'b01000111_00110011 : OUT <= 1;  //71 / 51 = 1
    16'b01000111_00110100 : OUT <= 1;  //71 / 52 = 1
    16'b01000111_00110101 : OUT <= 1;  //71 / 53 = 1
    16'b01000111_00110110 : OUT <= 1;  //71 / 54 = 1
    16'b01000111_00110111 : OUT <= 1;  //71 / 55 = 1
    16'b01000111_00111000 : OUT <= 1;  //71 / 56 = 1
    16'b01000111_00111001 : OUT <= 1;  //71 / 57 = 1
    16'b01000111_00111010 : OUT <= 1;  //71 / 58 = 1
    16'b01000111_00111011 : OUT <= 1;  //71 / 59 = 1
    16'b01000111_00111100 : OUT <= 1;  //71 / 60 = 1
    16'b01000111_00111101 : OUT <= 1;  //71 / 61 = 1
    16'b01000111_00111110 : OUT <= 1;  //71 / 62 = 1
    16'b01000111_00111111 : OUT <= 1;  //71 / 63 = 1
    16'b01000111_01000000 : OUT <= 1;  //71 / 64 = 1
    16'b01000111_01000001 : OUT <= 1;  //71 / 65 = 1
    16'b01000111_01000010 : OUT <= 1;  //71 / 66 = 1
    16'b01000111_01000011 : OUT <= 1;  //71 / 67 = 1
    16'b01000111_01000100 : OUT <= 1;  //71 / 68 = 1
    16'b01000111_01000101 : OUT <= 1;  //71 / 69 = 1
    16'b01000111_01000110 : OUT <= 1;  //71 / 70 = 1
    16'b01000111_01000111 : OUT <= 1;  //71 / 71 = 1
    16'b01000111_01001000 : OUT <= 0;  //71 / 72 = 0
    16'b01000111_01001001 : OUT <= 0;  //71 / 73 = 0
    16'b01000111_01001010 : OUT <= 0;  //71 / 74 = 0
    16'b01000111_01001011 : OUT <= 0;  //71 / 75 = 0
    16'b01000111_01001100 : OUT <= 0;  //71 / 76 = 0
    16'b01000111_01001101 : OUT <= 0;  //71 / 77 = 0
    16'b01000111_01001110 : OUT <= 0;  //71 / 78 = 0
    16'b01000111_01001111 : OUT <= 0;  //71 / 79 = 0
    16'b01000111_01010000 : OUT <= 0;  //71 / 80 = 0
    16'b01000111_01010001 : OUT <= 0;  //71 / 81 = 0
    16'b01000111_01010010 : OUT <= 0;  //71 / 82 = 0
    16'b01000111_01010011 : OUT <= 0;  //71 / 83 = 0
    16'b01000111_01010100 : OUT <= 0;  //71 / 84 = 0
    16'b01000111_01010101 : OUT <= 0;  //71 / 85 = 0
    16'b01000111_01010110 : OUT <= 0;  //71 / 86 = 0
    16'b01000111_01010111 : OUT <= 0;  //71 / 87 = 0
    16'b01000111_01011000 : OUT <= 0;  //71 / 88 = 0
    16'b01000111_01011001 : OUT <= 0;  //71 / 89 = 0
    16'b01000111_01011010 : OUT <= 0;  //71 / 90 = 0
    16'b01000111_01011011 : OUT <= 0;  //71 / 91 = 0
    16'b01000111_01011100 : OUT <= 0;  //71 / 92 = 0
    16'b01000111_01011101 : OUT <= 0;  //71 / 93 = 0
    16'b01000111_01011110 : OUT <= 0;  //71 / 94 = 0
    16'b01000111_01011111 : OUT <= 0;  //71 / 95 = 0
    16'b01000111_01100000 : OUT <= 0;  //71 / 96 = 0
    16'b01000111_01100001 : OUT <= 0;  //71 / 97 = 0
    16'b01000111_01100010 : OUT <= 0;  //71 / 98 = 0
    16'b01000111_01100011 : OUT <= 0;  //71 / 99 = 0
    16'b01000111_01100100 : OUT <= 0;  //71 / 100 = 0
    16'b01000111_01100101 : OUT <= 0;  //71 / 101 = 0
    16'b01000111_01100110 : OUT <= 0;  //71 / 102 = 0
    16'b01000111_01100111 : OUT <= 0;  //71 / 103 = 0
    16'b01000111_01101000 : OUT <= 0;  //71 / 104 = 0
    16'b01000111_01101001 : OUT <= 0;  //71 / 105 = 0
    16'b01000111_01101010 : OUT <= 0;  //71 / 106 = 0
    16'b01000111_01101011 : OUT <= 0;  //71 / 107 = 0
    16'b01000111_01101100 : OUT <= 0;  //71 / 108 = 0
    16'b01000111_01101101 : OUT <= 0;  //71 / 109 = 0
    16'b01000111_01101110 : OUT <= 0;  //71 / 110 = 0
    16'b01000111_01101111 : OUT <= 0;  //71 / 111 = 0
    16'b01000111_01110000 : OUT <= 0;  //71 / 112 = 0
    16'b01000111_01110001 : OUT <= 0;  //71 / 113 = 0
    16'b01000111_01110010 : OUT <= 0;  //71 / 114 = 0
    16'b01000111_01110011 : OUT <= 0;  //71 / 115 = 0
    16'b01000111_01110100 : OUT <= 0;  //71 / 116 = 0
    16'b01000111_01110101 : OUT <= 0;  //71 / 117 = 0
    16'b01000111_01110110 : OUT <= 0;  //71 / 118 = 0
    16'b01000111_01110111 : OUT <= 0;  //71 / 119 = 0
    16'b01000111_01111000 : OUT <= 0;  //71 / 120 = 0
    16'b01000111_01111001 : OUT <= 0;  //71 / 121 = 0
    16'b01000111_01111010 : OUT <= 0;  //71 / 122 = 0
    16'b01000111_01111011 : OUT <= 0;  //71 / 123 = 0
    16'b01000111_01111100 : OUT <= 0;  //71 / 124 = 0
    16'b01000111_01111101 : OUT <= 0;  //71 / 125 = 0
    16'b01000111_01111110 : OUT <= 0;  //71 / 126 = 0
    16'b01000111_01111111 : OUT <= 0;  //71 / 127 = 0
    16'b01000111_10000000 : OUT <= 0;  //71 / 128 = 0
    16'b01000111_10000001 : OUT <= 0;  //71 / 129 = 0
    16'b01000111_10000010 : OUT <= 0;  //71 / 130 = 0
    16'b01000111_10000011 : OUT <= 0;  //71 / 131 = 0
    16'b01000111_10000100 : OUT <= 0;  //71 / 132 = 0
    16'b01000111_10000101 : OUT <= 0;  //71 / 133 = 0
    16'b01000111_10000110 : OUT <= 0;  //71 / 134 = 0
    16'b01000111_10000111 : OUT <= 0;  //71 / 135 = 0
    16'b01000111_10001000 : OUT <= 0;  //71 / 136 = 0
    16'b01000111_10001001 : OUT <= 0;  //71 / 137 = 0
    16'b01000111_10001010 : OUT <= 0;  //71 / 138 = 0
    16'b01000111_10001011 : OUT <= 0;  //71 / 139 = 0
    16'b01000111_10001100 : OUT <= 0;  //71 / 140 = 0
    16'b01000111_10001101 : OUT <= 0;  //71 / 141 = 0
    16'b01000111_10001110 : OUT <= 0;  //71 / 142 = 0
    16'b01000111_10001111 : OUT <= 0;  //71 / 143 = 0
    16'b01000111_10010000 : OUT <= 0;  //71 / 144 = 0
    16'b01000111_10010001 : OUT <= 0;  //71 / 145 = 0
    16'b01000111_10010010 : OUT <= 0;  //71 / 146 = 0
    16'b01000111_10010011 : OUT <= 0;  //71 / 147 = 0
    16'b01000111_10010100 : OUT <= 0;  //71 / 148 = 0
    16'b01000111_10010101 : OUT <= 0;  //71 / 149 = 0
    16'b01000111_10010110 : OUT <= 0;  //71 / 150 = 0
    16'b01000111_10010111 : OUT <= 0;  //71 / 151 = 0
    16'b01000111_10011000 : OUT <= 0;  //71 / 152 = 0
    16'b01000111_10011001 : OUT <= 0;  //71 / 153 = 0
    16'b01000111_10011010 : OUT <= 0;  //71 / 154 = 0
    16'b01000111_10011011 : OUT <= 0;  //71 / 155 = 0
    16'b01000111_10011100 : OUT <= 0;  //71 / 156 = 0
    16'b01000111_10011101 : OUT <= 0;  //71 / 157 = 0
    16'b01000111_10011110 : OUT <= 0;  //71 / 158 = 0
    16'b01000111_10011111 : OUT <= 0;  //71 / 159 = 0
    16'b01000111_10100000 : OUT <= 0;  //71 / 160 = 0
    16'b01000111_10100001 : OUT <= 0;  //71 / 161 = 0
    16'b01000111_10100010 : OUT <= 0;  //71 / 162 = 0
    16'b01000111_10100011 : OUT <= 0;  //71 / 163 = 0
    16'b01000111_10100100 : OUT <= 0;  //71 / 164 = 0
    16'b01000111_10100101 : OUT <= 0;  //71 / 165 = 0
    16'b01000111_10100110 : OUT <= 0;  //71 / 166 = 0
    16'b01000111_10100111 : OUT <= 0;  //71 / 167 = 0
    16'b01000111_10101000 : OUT <= 0;  //71 / 168 = 0
    16'b01000111_10101001 : OUT <= 0;  //71 / 169 = 0
    16'b01000111_10101010 : OUT <= 0;  //71 / 170 = 0
    16'b01000111_10101011 : OUT <= 0;  //71 / 171 = 0
    16'b01000111_10101100 : OUT <= 0;  //71 / 172 = 0
    16'b01000111_10101101 : OUT <= 0;  //71 / 173 = 0
    16'b01000111_10101110 : OUT <= 0;  //71 / 174 = 0
    16'b01000111_10101111 : OUT <= 0;  //71 / 175 = 0
    16'b01000111_10110000 : OUT <= 0;  //71 / 176 = 0
    16'b01000111_10110001 : OUT <= 0;  //71 / 177 = 0
    16'b01000111_10110010 : OUT <= 0;  //71 / 178 = 0
    16'b01000111_10110011 : OUT <= 0;  //71 / 179 = 0
    16'b01000111_10110100 : OUT <= 0;  //71 / 180 = 0
    16'b01000111_10110101 : OUT <= 0;  //71 / 181 = 0
    16'b01000111_10110110 : OUT <= 0;  //71 / 182 = 0
    16'b01000111_10110111 : OUT <= 0;  //71 / 183 = 0
    16'b01000111_10111000 : OUT <= 0;  //71 / 184 = 0
    16'b01000111_10111001 : OUT <= 0;  //71 / 185 = 0
    16'b01000111_10111010 : OUT <= 0;  //71 / 186 = 0
    16'b01000111_10111011 : OUT <= 0;  //71 / 187 = 0
    16'b01000111_10111100 : OUT <= 0;  //71 / 188 = 0
    16'b01000111_10111101 : OUT <= 0;  //71 / 189 = 0
    16'b01000111_10111110 : OUT <= 0;  //71 / 190 = 0
    16'b01000111_10111111 : OUT <= 0;  //71 / 191 = 0
    16'b01000111_11000000 : OUT <= 0;  //71 / 192 = 0
    16'b01000111_11000001 : OUT <= 0;  //71 / 193 = 0
    16'b01000111_11000010 : OUT <= 0;  //71 / 194 = 0
    16'b01000111_11000011 : OUT <= 0;  //71 / 195 = 0
    16'b01000111_11000100 : OUT <= 0;  //71 / 196 = 0
    16'b01000111_11000101 : OUT <= 0;  //71 / 197 = 0
    16'b01000111_11000110 : OUT <= 0;  //71 / 198 = 0
    16'b01000111_11000111 : OUT <= 0;  //71 / 199 = 0
    16'b01000111_11001000 : OUT <= 0;  //71 / 200 = 0
    16'b01000111_11001001 : OUT <= 0;  //71 / 201 = 0
    16'b01000111_11001010 : OUT <= 0;  //71 / 202 = 0
    16'b01000111_11001011 : OUT <= 0;  //71 / 203 = 0
    16'b01000111_11001100 : OUT <= 0;  //71 / 204 = 0
    16'b01000111_11001101 : OUT <= 0;  //71 / 205 = 0
    16'b01000111_11001110 : OUT <= 0;  //71 / 206 = 0
    16'b01000111_11001111 : OUT <= 0;  //71 / 207 = 0
    16'b01000111_11010000 : OUT <= 0;  //71 / 208 = 0
    16'b01000111_11010001 : OUT <= 0;  //71 / 209 = 0
    16'b01000111_11010010 : OUT <= 0;  //71 / 210 = 0
    16'b01000111_11010011 : OUT <= 0;  //71 / 211 = 0
    16'b01000111_11010100 : OUT <= 0;  //71 / 212 = 0
    16'b01000111_11010101 : OUT <= 0;  //71 / 213 = 0
    16'b01000111_11010110 : OUT <= 0;  //71 / 214 = 0
    16'b01000111_11010111 : OUT <= 0;  //71 / 215 = 0
    16'b01000111_11011000 : OUT <= 0;  //71 / 216 = 0
    16'b01000111_11011001 : OUT <= 0;  //71 / 217 = 0
    16'b01000111_11011010 : OUT <= 0;  //71 / 218 = 0
    16'b01000111_11011011 : OUT <= 0;  //71 / 219 = 0
    16'b01000111_11011100 : OUT <= 0;  //71 / 220 = 0
    16'b01000111_11011101 : OUT <= 0;  //71 / 221 = 0
    16'b01000111_11011110 : OUT <= 0;  //71 / 222 = 0
    16'b01000111_11011111 : OUT <= 0;  //71 / 223 = 0
    16'b01000111_11100000 : OUT <= 0;  //71 / 224 = 0
    16'b01000111_11100001 : OUT <= 0;  //71 / 225 = 0
    16'b01000111_11100010 : OUT <= 0;  //71 / 226 = 0
    16'b01000111_11100011 : OUT <= 0;  //71 / 227 = 0
    16'b01000111_11100100 : OUT <= 0;  //71 / 228 = 0
    16'b01000111_11100101 : OUT <= 0;  //71 / 229 = 0
    16'b01000111_11100110 : OUT <= 0;  //71 / 230 = 0
    16'b01000111_11100111 : OUT <= 0;  //71 / 231 = 0
    16'b01000111_11101000 : OUT <= 0;  //71 / 232 = 0
    16'b01000111_11101001 : OUT <= 0;  //71 / 233 = 0
    16'b01000111_11101010 : OUT <= 0;  //71 / 234 = 0
    16'b01000111_11101011 : OUT <= 0;  //71 / 235 = 0
    16'b01000111_11101100 : OUT <= 0;  //71 / 236 = 0
    16'b01000111_11101101 : OUT <= 0;  //71 / 237 = 0
    16'b01000111_11101110 : OUT <= 0;  //71 / 238 = 0
    16'b01000111_11101111 : OUT <= 0;  //71 / 239 = 0
    16'b01000111_11110000 : OUT <= 0;  //71 / 240 = 0
    16'b01000111_11110001 : OUT <= 0;  //71 / 241 = 0
    16'b01000111_11110010 : OUT <= 0;  //71 / 242 = 0
    16'b01000111_11110011 : OUT <= 0;  //71 / 243 = 0
    16'b01000111_11110100 : OUT <= 0;  //71 / 244 = 0
    16'b01000111_11110101 : OUT <= 0;  //71 / 245 = 0
    16'b01000111_11110110 : OUT <= 0;  //71 / 246 = 0
    16'b01000111_11110111 : OUT <= 0;  //71 / 247 = 0
    16'b01000111_11111000 : OUT <= 0;  //71 / 248 = 0
    16'b01000111_11111001 : OUT <= 0;  //71 / 249 = 0
    16'b01000111_11111010 : OUT <= 0;  //71 / 250 = 0
    16'b01000111_11111011 : OUT <= 0;  //71 / 251 = 0
    16'b01000111_11111100 : OUT <= 0;  //71 / 252 = 0
    16'b01000111_11111101 : OUT <= 0;  //71 / 253 = 0
    16'b01000111_11111110 : OUT <= 0;  //71 / 254 = 0
    16'b01000111_11111111 : OUT <= 0;  //71 / 255 = 0
    16'b01001000_00000000 : OUT <= 0;  //72 / 0 = 0
    16'b01001000_00000001 : OUT <= 72;  //72 / 1 = 72
    16'b01001000_00000010 : OUT <= 36;  //72 / 2 = 36
    16'b01001000_00000011 : OUT <= 24;  //72 / 3 = 24
    16'b01001000_00000100 : OUT <= 18;  //72 / 4 = 18
    16'b01001000_00000101 : OUT <= 14;  //72 / 5 = 14
    16'b01001000_00000110 : OUT <= 12;  //72 / 6 = 12
    16'b01001000_00000111 : OUT <= 10;  //72 / 7 = 10
    16'b01001000_00001000 : OUT <= 9;  //72 / 8 = 9
    16'b01001000_00001001 : OUT <= 8;  //72 / 9 = 8
    16'b01001000_00001010 : OUT <= 7;  //72 / 10 = 7
    16'b01001000_00001011 : OUT <= 6;  //72 / 11 = 6
    16'b01001000_00001100 : OUT <= 6;  //72 / 12 = 6
    16'b01001000_00001101 : OUT <= 5;  //72 / 13 = 5
    16'b01001000_00001110 : OUT <= 5;  //72 / 14 = 5
    16'b01001000_00001111 : OUT <= 4;  //72 / 15 = 4
    16'b01001000_00010000 : OUT <= 4;  //72 / 16 = 4
    16'b01001000_00010001 : OUT <= 4;  //72 / 17 = 4
    16'b01001000_00010010 : OUT <= 4;  //72 / 18 = 4
    16'b01001000_00010011 : OUT <= 3;  //72 / 19 = 3
    16'b01001000_00010100 : OUT <= 3;  //72 / 20 = 3
    16'b01001000_00010101 : OUT <= 3;  //72 / 21 = 3
    16'b01001000_00010110 : OUT <= 3;  //72 / 22 = 3
    16'b01001000_00010111 : OUT <= 3;  //72 / 23 = 3
    16'b01001000_00011000 : OUT <= 3;  //72 / 24 = 3
    16'b01001000_00011001 : OUT <= 2;  //72 / 25 = 2
    16'b01001000_00011010 : OUT <= 2;  //72 / 26 = 2
    16'b01001000_00011011 : OUT <= 2;  //72 / 27 = 2
    16'b01001000_00011100 : OUT <= 2;  //72 / 28 = 2
    16'b01001000_00011101 : OUT <= 2;  //72 / 29 = 2
    16'b01001000_00011110 : OUT <= 2;  //72 / 30 = 2
    16'b01001000_00011111 : OUT <= 2;  //72 / 31 = 2
    16'b01001000_00100000 : OUT <= 2;  //72 / 32 = 2
    16'b01001000_00100001 : OUT <= 2;  //72 / 33 = 2
    16'b01001000_00100010 : OUT <= 2;  //72 / 34 = 2
    16'b01001000_00100011 : OUT <= 2;  //72 / 35 = 2
    16'b01001000_00100100 : OUT <= 2;  //72 / 36 = 2
    16'b01001000_00100101 : OUT <= 1;  //72 / 37 = 1
    16'b01001000_00100110 : OUT <= 1;  //72 / 38 = 1
    16'b01001000_00100111 : OUT <= 1;  //72 / 39 = 1
    16'b01001000_00101000 : OUT <= 1;  //72 / 40 = 1
    16'b01001000_00101001 : OUT <= 1;  //72 / 41 = 1
    16'b01001000_00101010 : OUT <= 1;  //72 / 42 = 1
    16'b01001000_00101011 : OUT <= 1;  //72 / 43 = 1
    16'b01001000_00101100 : OUT <= 1;  //72 / 44 = 1
    16'b01001000_00101101 : OUT <= 1;  //72 / 45 = 1
    16'b01001000_00101110 : OUT <= 1;  //72 / 46 = 1
    16'b01001000_00101111 : OUT <= 1;  //72 / 47 = 1
    16'b01001000_00110000 : OUT <= 1;  //72 / 48 = 1
    16'b01001000_00110001 : OUT <= 1;  //72 / 49 = 1
    16'b01001000_00110010 : OUT <= 1;  //72 / 50 = 1
    16'b01001000_00110011 : OUT <= 1;  //72 / 51 = 1
    16'b01001000_00110100 : OUT <= 1;  //72 / 52 = 1
    16'b01001000_00110101 : OUT <= 1;  //72 / 53 = 1
    16'b01001000_00110110 : OUT <= 1;  //72 / 54 = 1
    16'b01001000_00110111 : OUT <= 1;  //72 / 55 = 1
    16'b01001000_00111000 : OUT <= 1;  //72 / 56 = 1
    16'b01001000_00111001 : OUT <= 1;  //72 / 57 = 1
    16'b01001000_00111010 : OUT <= 1;  //72 / 58 = 1
    16'b01001000_00111011 : OUT <= 1;  //72 / 59 = 1
    16'b01001000_00111100 : OUT <= 1;  //72 / 60 = 1
    16'b01001000_00111101 : OUT <= 1;  //72 / 61 = 1
    16'b01001000_00111110 : OUT <= 1;  //72 / 62 = 1
    16'b01001000_00111111 : OUT <= 1;  //72 / 63 = 1
    16'b01001000_01000000 : OUT <= 1;  //72 / 64 = 1
    16'b01001000_01000001 : OUT <= 1;  //72 / 65 = 1
    16'b01001000_01000010 : OUT <= 1;  //72 / 66 = 1
    16'b01001000_01000011 : OUT <= 1;  //72 / 67 = 1
    16'b01001000_01000100 : OUT <= 1;  //72 / 68 = 1
    16'b01001000_01000101 : OUT <= 1;  //72 / 69 = 1
    16'b01001000_01000110 : OUT <= 1;  //72 / 70 = 1
    16'b01001000_01000111 : OUT <= 1;  //72 / 71 = 1
    16'b01001000_01001000 : OUT <= 1;  //72 / 72 = 1
    16'b01001000_01001001 : OUT <= 0;  //72 / 73 = 0
    16'b01001000_01001010 : OUT <= 0;  //72 / 74 = 0
    16'b01001000_01001011 : OUT <= 0;  //72 / 75 = 0
    16'b01001000_01001100 : OUT <= 0;  //72 / 76 = 0
    16'b01001000_01001101 : OUT <= 0;  //72 / 77 = 0
    16'b01001000_01001110 : OUT <= 0;  //72 / 78 = 0
    16'b01001000_01001111 : OUT <= 0;  //72 / 79 = 0
    16'b01001000_01010000 : OUT <= 0;  //72 / 80 = 0
    16'b01001000_01010001 : OUT <= 0;  //72 / 81 = 0
    16'b01001000_01010010 : OUT <= 0;  //72 / 82 = 0
    16'b01001000_01010011 : OUT <= 0;  //72 / 83 = 0
    16'b01001000_01010100 : OUT <= 0;  //72 / 84 = 0
    16'b01001000_01010101 : OUT <= 0;  //72 / 85 = 0
    16'b01001000_01010110 : OUT <= 0;  //72 / 86 = 0
    16'b01001000_01010111 : OUT <= 0;  //72 / 87 = 0
    16'b01001000_01011000 : OUT <= 0;  //72 / 88 = 0
    16'b01001000_01011001 : OUT <= 0;  //72 / 89 = 0
    16'b01001000_01011010 : OUT <= 0;  //72 / 90 = 0
    16'b01001000_01011011 : OUT <= 0;  //72 / 91 = 0
    16'b01001000_01011100 : OUT <= 0;  //72 / 92 = 0
    16'b01001000_01011101 : OUT <= 0;  //72 / 93 = 0
    16'b01001000_01011110 : OUT <= 0;  //72 / 94 = 0
    16'b01001000_01011111 : OUT <= 0;  //72 / 95 = 0
    16'b01001000_01100000 : OUT <= 0;  //72 / 96 = 0
    16'b01001000_01100001 : OUT <= 0;  //72 / 97 = 0
    16'b01001000_01100010 : OUT <= 0;  //72 / 98 = 0
    16'b01001000_01100011 : OUT <= 0;  //72 / 99 = 0
    16'b01001000_01100100 : OUT <= 0;  //72 / 100 = 0
    16'b01001000_01100101 : OUT <= 0;  //72 / 101 = 0
    16'b01001000_01100110 : OUT <= 0;  //72 / 102 = 0
    16'b01001000_01100111 : OUT <= 0;  //72 / 103 = 0
    16'b01001000_01101000 : OUT <= 0;  //72 / 104 = 0
    16'b01001000_01101001 : OUT <= 0;  //72 / 105 = 0
    16'b01001000_01101010 : OUT <= 0;  //72 / 106 = 0
    16'b01001000_01101011 : OUT <= 0;  //72 / 107 = 0
    16'b01001000_01101100 : OUT <= 0;  //72 / 108 = 0
    16'b01001000_01101101 : OUT <= 0;  //72 / 109 = 0
    16'b01001000_01101110 : OUT <= 0;  //72 / 110 = 0
    16'b01001000_01101111 : OUT <= 0;  //72 / 111 = 0
    16'b01001000_01110000 : OUT <= 0;  //72 / 112 = 0
    16'b01001000_01110001 : OUT <= 0;  //72 / 113 = 0
    16'b01001000_01110010 : OUT <= 0;  //72 / 114 = 0
    16'b01001000_01110011 : OUT <= 0;  //72 / 115 = 0
    16'b01001000_01110100 : OUT <= 0;  //72 / 116 = 0
    16'b01001000_01110101 : OUT <= 0;  //72 / 117 = 0
    16'b01001000_01110110 : OUT <= 0;  //72 / 118 = 0
    16'b01001000_01110111 : OUT <= 0;  //72 / 119 = 0
    16'b01001000_01111000 : OUT <= 0;  //72 / 120 = 0
    16'b01001000_01111001 : OUT <= 0;  //72 / 121 = 0
    16'b01001000_01111010 : OUT <= 0;  //72 / 122 = 0
    16'b01001000_01111011 : OUT <= 0;  //72 / 123 = 0
    16'b01001000_01111100 : OUT <= 0;  //72 / 124 = 0
    16'b01001000_01111101 : OUT <= 0;  //72 / 125 = 0
    16'b01001000_01111110 : OUT <= 0;  //72 / 126 = 0
    16'b01001000_01111111 : OUT <= 0;  //72 / 127 = 0
    16'b01001000_10000000 : OUT <= 0;  //72 / 128 = 0
    16'b01001000_10000001 : OUT <= 0;  //72 / 129 = 0
    16'b01001000_10000010 : OUT <= 0;  //72 / 130 = 0
    16'b01001000_10000011 : OUT <= 0;  //72 / 131 = 0
    16'b01001000_10000100 : OUT <= 0;  //72 / 132 = 0
    16'b01001000_10000101 : OUT <= 0;  //72 / 133 = 0
    16'b01001000_10000110 : OUT <= 0;  //72 / 134 = 0
    16'b01001000_10000111 : OUT <= 0;  //72 / 135 = 0
    16'b01001000_10001000 : OUT <= 0;  //72 / 136 = 0
    16'b01001000_10001001 : OUT <= 0;  //72 / 137 = 0
    16'b01001000_10001010 : OUT <= 0;  //72 / 138 = 0
    16'b01001000_10001011 : OUT <= 0;  //72 / 139 = 0
    16'b01001000_10001100 : OUT <= 0;  //72 / 140 = 0
    16'b01001000_10001101 : OUT <= 0;  //72 / 141 = 0
    16'b01001000_10001110 : OUT <= 0;  //72 / 142 = 0
    16'b01001000_10001111 : OUT <= 0;  //72 / 143 = 0
    16'b01001000_10010000 : OUT <= 0;  //72 / 144 = 0
    16'b01001000_10010001 : OUT <= 0;  //72 / 145 = 0
    16'b01001000_10010010 : OUT <= 0;  //72 / 146 = 0
    16'b01001000_10010011 : OUT <= 0;  //72 / 147 = 0
    16'b01001000_10010100 : OUT <= 0;  //72 / 148 = 0
    16'b01001000_10010101 : OUT <= 0;  //72 / 149 = 0
    16'b01001000_10010110 : OUT <= 0;  //72 / 150 = 0
    16'b01001000_10010111 : OUT <= 0;  //72 / 151 = 0
    16'b01001000_10011000 : OUT <= 0;  //72 / 152 = 0
    16'b01001000_10011001 : OUT <= 0;  //72 / 153 = 0
    16'b01001000_10011010 : OUT <= 0;  //72 / 154 = 0
    16'b01001000_10011011 : OUT <= 0;  //72 / 155 = 0
    16'b01001000_10011100 : OUT <= 0;  //72 / 156 = 0
    16'b01001000_10011101 : OUT <= 0;  //72 / 157 = 0
    16'b01001000_10011110 : OUT <= 0;  //72 / 158 = 0
    16'b01001000_10011111 : OUT <= 0;  //72 / 159 = 0
    16'b01001000_10100000 : OUT <= 0;  //72 / 160 = 0
    16'b01001000_10100001 : OUT <= 0;  //72 / 161 = 0
    16'b01001000_10100010 : OUT <= 0;  //72 / 162 = 0
    16'b01001000_10100011 : OUT <= 0;  //72 / 163 = 0
    16'b01001000_10100100 : OUT <= 0;  //72 / 164 = 0
    16'b01001000_10100101 : OUT <= 0;  //72 / 165 = 0
    16'b01001000_10100110 : OUT <= 0;  //72 / 166 = 0
    16'b01001000_10100111 : OUT <= 0;  //72 / 167 = 0
    16'b01001000_10101000 : OUT <= 0;  //72 / 168 = 0
    16'b01001000_10101001 : OUT <= 0;  //72 / 169 = 0
    16'b01001000_10101010 : OUT <= 0;  //72 / 170 = 0
    16'b01001000_10101011 : OUT <= 0;  //72 / 171 = 0
    16'b01001000_10101100 : OUT <= 0;  //72 / 172 = 0
    16'b01001000_10101101 : OUT <= 0;  //72 / 173 = 0
    16'b01001000_10101110 : OUT <= 0;  //72 / 174 = 0
    16'b01001000_10101111 : OUT <= 0;  //72 / 175 = 0
    16'b01001000_10110000 : OUT <= 0;  //72 / 176 = 0
    16'b01001000_10110001 : OUT <= 0;  //72 / 177 = 0
    16'b01001000_10110010 : OUT <= 0;  //72 / 178 = 0
    16'b01001000_10110011 : OUT <= 0;  //72 / 179 = 0
    16'b01001000_10110100 : OUT <= 0;  //72 / 180 = 0
    16'b01001000_10110101 : OUT <= 0;  //72 / 181 = 0
    16'b01001000_10110110 : OUT <= 0;  //72 / 182 = 0
    16'b01001000_10110111 : OUT <= 0;  //72 / 183 = 0
    16'b01001000_10111000 : OUT <= 0;  //72 / 184 = 0
    16'b01001000_10111001 : OUT <= 0;  //72 / 185 = 0
    16'b01001000_10111010 : OUT <= 0;  //72 / 186 = 0
    16'b01001000_10111011 : OUT <= 0;  //72 / 187 = 0
    16'b01001000_10111100 : OUT <= 0;  //72 / 188 = 0
    16'b01001000_10111101 : OUT <= 0;  //72 / 189 = 0
    16'b01001000_10111110 : OUT <= 0;  //72 / 190 = 0
    16'b01001000_10111111 : OUT <= 0;  //72 / 191 = 0
    16'b01001000_11000000 : OUT <= 0;  //72 / 192 = 0
    16'b01001000_11000001 : OUT <= 0;  //72 / 193 = 0
    16'b01001000_11000010 : OUT <= 0;  //72 / 194 = 0
    16'b01001000_11000011 : OUT <= 0;  //72 / 195 = 0
    16'b01001000_11000100 : OUT <= 0;  //72 / 196 = 0
    16'b01001000_11000101 : OUT <= 0;  //72 / 197 = 0
    16'b01001000_11000110 : OUT <= 0;  //72 / 198 = 0
    16'b01001000_11000111 : OUT <= 0;  //72 / 199 = 0
    16'b01001000_11001000 : OUT <= 0;  //72 / 200 = 0
    16'b01001000_11001001 : OUT <= 0;  //72 / 201 = 0
    16'b01001000_11001010 : OUT <= 0;  //72 / 202 = 0
    16'b01001000_11001011 : OUT <= 0;  //72 / 203 = 0
    16'b01001000_11001100 : OUT <= 0;  //72 / 204 = 0
    16'b01001000_11001101 : OUT <= 0;  //72 / 205 = 0
    16'b01001000_11001110 : OUT <= 0;  //72 / 206 = 0
    16'b01001000_11001111 : OUT <= 0;  //72 / 207 = 0
    16'b01001000_11010000 : OUT <= 0;  //72 / 208 = 0
    16'b01001000_11010001 : OUT <= 0;  //72 / 209 = 0
    16'b01001000_11010010 : OUT <= 0;  //72 / 210 = 0
    16'b01001000_11010011 : OUT <= 0;  //72 / 211 = 0
    16'b01001000_11010100 : OUT <= 0;  //72 / 212 = 0
    16'b01001000_11010101 : OUT <= 0;  //72 / 213 = 0
    16'b01001000_11010110 : OUT <= 0;  //72 / 214 = 0
    16'b01001000_11010111 : OUT <= 0;  //72 / 215 = 0
    16'b01001000_11011000 : OUT <= 0;  //72 / 216 = 0
    16'b01001000_11011001 : OUT <= 0;  //72 / 217 = 0
    16'b01001000_11011010 : OUT <= 0;  //72 / 218 = 0
    16'b01001000_11011011 : OUT <= 0;  //72 / 219 = 0
    16'b01001000_11011100 : OUT <= 0;  //72 / 220 = 0
    16'b01001000_11011101 : OUT <= 0;  //72 / 221 = 0
    16'b01001000_11011110 : OUT <= 0;  //72 / 222 = 0
    16'b01001000_11011111 : OUT <= 0;  //72 / 223 = 0
    16'b01001000_11100000 : OUT <= 0;  //72 / 224 = 0
    16'b01001000_11100001 : OUT <= 0;  //72 / 225 = 0
    16'b01001000_11100010 : OUT <= 0;  //72 / 226 = 0
    16'b01001000_11100011 : OUT <= 0;  //72 / 227 = 0
    16'b01001000_11100100 : OUT <= 0;  //72 / 228 = 0
    16'b01001000_11100101 : OUT <= 0;  //72 / 229 = 0
    16'b01001000_11100110 : OUT <= 0;  //72 / 230 = 0
    16'b01001000_11100111 : OUT <= 0;  //72 / 231 = 0
    16'b01001000_11101000 : OUT <= 0;  //72 / 232 = 0
    16'b01001000_11101001 : OUT <= 0;  //72 / 233 = 0
    16'b01001000_11101010 : OUT <= 0;  //72 / 234 = 0
    16'b01001000_11101011 : OUT <= 0;  //72 / 235 = 0
    16'b01001000_11101100 : OUT <= 0;  //72 / 236 = 0
    16'b01001000_11101101 : OUT <= 0;  //72 / 237 = 0
    16'b01001000_11101110 : OUT <= 0;  //72 / 238 = 0
    16'b01001000_11101111 : OUT <= 0;  //72 / 239 = 0
    16'b01001000_11110000 : OUT <= 0;  //72 / 240 = 0
    16'b01001000_11110001 : OUT <= 0;  //72 / 241 = 0
    16'b01001000_11110010 : OUT <= 0;  //72 / 242 = 0
    16'b01001000_11110011 : OUT <= 0;  //72 / 243 = 0
    16'b01001000_11110100 : OUT <= 0;  //72 / 244 = 0
    16'b01001000_11110101 : OUT <= 0;  //72 / 245 = 0
    16'b01001000_11110110 : OUT <= 0;  //72 / 246 = 0
    16'b01001000_11110111 : OUT <= 0;  //72 / 247 = 0
    16'b01001000_11111000 : OUT <= 0;  //72 / 248 = 0
    16'b01001000_11111001 : OUT <= 0;  //72 / 249 = 0
    16'b01001000_11111010 : OUT <= 0;  //72 / 250 = 0
    16'b01001000_11111011 : OUT <= 0;  //72 / 251 = 0
    16'b01001000_11111100 : OUT <= 0;  //72 / 252 = 0
    16'b01001000_11111101 : OUT <= 0;  //72 / 253 = 0
    16'b01001000_11111110 : OUT <= 0;  //72 / 254 = 0
    16'b01001000_11111111 : OUT <= 0;  //72 / 255 = 0
    16'b01001001_00000000 : OUT <= 0;  //73 / 0 = 0
    16'b01001001_00000001 : OUT <= 73;  //73 / 1 = 73
    16'b01001001_00000010 : OUT <= 36;  //73 / 2 = 36
    16'b01001001_00000011 : OUT <= 24;  //73 / 3 = 24
    16'b01001001_00000100 : OUT <= 18;  //73 / 4 = 18
    16'b01001001_00000101 : OUT <= 14;  //73 / 5 = 14
    16'b01001001_00000110 : OUT <= 12;  //73 / 6 = 12
    16'b01001001_00000111 : OUT <= 10;  //73 / 7 = 10
    16'b01001001_00001000 : OUT <= 9;  //73 / 8 = 9
    16'b01001001_00001001 : OUT <= 8;  //73 / 9 = 8
    16'b01001001_00001010 : OUT <= 7;  //73 / 10 = 7
    16'b01001001_00001011 : OUT <= 6;  //73 / 11 = 6
    16'b01001001_00001100 : OUT <= 6;  //73 / 12 = 6
    16'b01001001_00001101 : OUT <= 5;  //73 / 13 = 5
    16'b01001001_00001110 : OUT <= 5;  //73 / 14 = 5
    16'b01001001_00001111 : OUT <= 4;  //73 / 15 = 4
    16'b01001001_00010000 : OUT <= 4;  //73 / 16 = 4
    16'b01001001_00010001 : OUT <= 4;  //73 / 17 = 4
    16'b01001001_00010010 : OUT <= 4;  //73 / 18 = 4
    16'b01001001_00010011 : OUT <= 3;  //73 / 19 = 3
    16'b01001001_00010100 : OUT <= 3;  //73 / 20 = 3
    16'b01001001_00010101 : OUT <= 3;  //73 / 21 = 3
    16'b01001001_00010110 : OUT <= 3;  //73 / 22 = 3
    16'b01001001_00010111 : OUT <= 3;  //73 / 23 = 3
    16'b01001001_00011000 : OUT <= 3;  //73 / 24 = 3
    16'b01001001_00011001 : OUT <= 2;  //73 / 25 = 2
    16'b01001001_00011010 : OUT <= 2;  //73 / 26 = 2
    16'b01001001_00011011 : OUT <= 2;  //73 / 27 = 2
    16'b01001001_00011100 : OUT <= 2;  //73 / 28 = 2
    16'b01001001_00011101 : OUT <= 2;  //73 / 29 = 2
    16'b01001001_00011110 : OUT <= 2;  //73 / 30 = 2
    16'b01001001_00011111 : OUT <= 2;  //73 / 31 = 2
    16'b01001001_00100000 : OUT <= 2;  //73 / 32 = 2
    16'b01001001_00100001 : OUT <= 2;  //73 / 33 = 2
    16'b01001001_00100010 : OUT <= 2;  //73 / 34 = 2
    16'b01001001_00100011 : OUT <= 2;  //73 / 35 = 2
    16'b01001001_00100100 : OUT <= 2;  //73 / 36 = 2
    16'b01001001_00100101 : OUT <= 1;  //73 / 37 = 1
    16'b01001001_00100110 : OUT <= 1;  //73 / 38 = 1
    16'b01001001_00100111 : OUT <= 1;  //73 / 39 = 1
    16'b01001001_00101000 : OUT <= 1;  //73 / 40 = 1
    16'b01001001_00101001 : OUT <= 1;  //73 / 41 = 1
    16'b01001001_00101010 : OUT <= 1;  //73 / 42 = 1
    16'b01001001_00101011 : OUT <= 1;  //73 / 43 = 1
    16'b01001001_00101100 : OUT <= 1;  //73 / 44 = 1
    16'b01001001_00101101 : OUT <= 1;  //73 / 45 = 1
    16'b01001001_00101110 : OUT <= 1;  //73 / 46 = 1
    16'b01001001_00101111 : OUT <= 1;  //73 / 47 = 1
    16'b01001001_00110000 : OUT <= 1;  //73 / 48 = 1
    16'b01001001_00110001 : OUT <= 1;  //73 / 49 = 1
    16'b01001001_00110010 : OUT <= 1;  //73 / 50 = 1
    16'b01001001_00110011 : OUT <= 1;  //73 / 51 = 1
    16'b01001001_00110100 : OUT <= 1;  //73 / 52 = 1
    16'b01001001_00110101 : OUT <= 1;  //73 / 53 = 1
    16'b01001001_00110110 : OUT <= 1;  //73 / 54 = 1
    16'b01001001_00110111 : OUT <= 1;  //73 / 55 = 1
    16'b01001001_00111000 : OUT <= 1;  //73 / 56 = 1
    16'b01001001_00111001 : OUT <= 1;  //73 / 57 = 1
    16'b01001001_00111010 : OUT <= 1;  //73 / 58 = 1
    16'b01001001_00111011 : OUT <= 1;  //73 / 59 = 1
    16'b01001001_00111100 : OUT <= 1;  //73 / 60 = 1
    16'b01001001_00111101 : OUT <= 1;  //73 / 61 = 1
    16'b01001001_00111110 : OUT <= 1;  //73 / 62 = 1
    16'b01001001_00111111 : OUT <= 1;  //73 / 63 = 1
    16'b01001001_01000000 : OUT <= 1;  //73 / 64 = 1
    16'b01001001_01000001 : OUT <= 1;  //73 / 65 = 1
    16'b01001001_01000010 : OUT <= 1;  //73 / 66 = 1
    16'b01001001_01000011 : OUT <= 1;  //73 / 67 = 1
    16'b01001001_01000100 : OUT <= 1;  //73 / 68 = 1
    16'b01001001_01000101 : OUT <= 1;  //73 / 69 = 1
    16'b01001001_01000110 : OUT <= 1;  //73 / 70 = 1
    16'b01001001_01000111 : OUT <= 1;  //73 / 71 = 1
    16'b01001001_01001000 : OUT <= 1;  //73 / 72 = 1
    16'b01001001_01001001 : OUT <= 1;  //73 / 73 = 1
    16'b01001001_01001010 : OUT <= 0;  //73 / 74 = 0
    16'b01001001_01001011 : OUT <= 0;  //73 / 75 = 0
    16'b01001001_01001100 : OUT <= 0;  //73 / 76 = 0
    16'b01001001_01001101 : OUT <= 0;  //73 / 77 = 0
    16'b01001001_01001110 : OUT <= 0;  //73 / 78 = 0
    16'b01001001_01001111 : OUT <= 0;  //73 / 79 = 0
    16'b01001001_01010000 : OUT <= 0;  //73 / 80 = 0
    16'b01001001_01010001 : OUT <= 0;  //73 / 81 = 0
    16'b01001001_01010010 : OUT <= 0;  //73 / 82 = 0
    16'b01001001_01010011 : OUT <= 0;  //73 / 83 = 0
    16'b01001001_01010100 : OUT <= 0;  //73 / 84 = 0
    16'b01001001_01010101 : OUT <= 0;  //73 / 85 = 0
    16'b01001001_01010110 : OUT <= 0;  //73 / 86 = 0
    16'b01001001_01010111 : OUT <= 0;  //73 / 87 = 0
    16'b01001001_01011000 : OUT <= 0;  //73 / 88 = 0
    16'b01001001_01011001 : OUT <= 0;  //73 / 89 = 0
    16'b01001001_01011010 : OUT <= 0;  //73 / 90 = 0
    16'b01001001_01011011 : OUT <= 0;  //73 / 91 = 0
    16'b01001001_01011100 : OUT <= 0;  //73 / 92 = 0
    16'b01001001_01011101 : OUT <= 0;  //73 / 93 = 0
    16'b01001001_01011110 : OUT <= 0;  //73 / 94 = 0
    16'b01001001_01011111 : OUT <= 0;  //73 / 95 = 0
    16'b01001001_01100000 : OUT <= 0;  //73 / 96 = 0
    16'b01001001_01100001 : OUT <= 0;  //73 / 97 = 0
    16'b01001001_01100010 : OUT <= 0;  //73 / 98 = 0
    16'b01001001_01100011 : OUT <= 0;  //73 / 99 = 0
    16'b01001001_01100100 : OUT <= 0;  //73 / 100 = 0
    16'b01001001_01100101 : OUT <= 0;  //73 / 101 = 0
    16'b01001001_01100110 : OUT <= 0;  //73 / 102 = 0
    16'b01001001_01100111 : OUT <= 0;  //73 / 103 = 0
    16'b01001001_01101000 : OUT <= 0;  //73 / 104 = 0
    16'b01001001_01101001 : OUT <= 0;  //73 / 105 = 0
    16'b01001001_01101010 : OUT <= 0;  //73 / 106 = 0
    16'b01001001_01101011 : OUT <= 0;  //73 / 107 = 0
    16'b01001001_01101100 : OUT <= 0;  //73 / 108 = 0
    16'b01001001_01101101 : OUT <= 0;  //73 / 109 = 0
    16'b01001001_01101110 : OUT <= 0;  //73 / 110 = 0
    16'b01001001_01101111 : OUT <= 0;  //73 / 111 = 0
    16'b01001001_01110000 : OUT <= 0;  //73 / 112 = 0
    16'b01001001_01110001 : OUT <= 0;  //73 / 113 = 0
    16'b01001001_01110010 : OUT <= 0;  //73 / 114 = 0
    16'b01001001_01110011 : OUT <= 0;  //73 / 115 = 0
    16'b01001001_01110100 : OUT <= 0;  //73 / 116 = 0
    16'b01001001_01110101 : OUT <= 0;  //73 / 117 = 0
    16'b01001001_01110110 : OUT <= 0;  //73 / 118 = 0
    16'b01001001_01110111 : OUT <= 0;  //73 / 119 = 0
    16'b01001001_01111000 : OUT <= 0;  //73 / 120 = 0
    16'b01001001_01111001 : OUT <= 0;  //73 / 121 = 0
    16'b01001001_01111010 : OUT <= 0;  //73 / 122 = 0
    16'b01001001_01111011 : OUT <= 0;  //73 / 123 = 0
    16'b01001001_01111100 : OUT <= 0;  //73 / 124 = 0
    16'b01001001_01111101 : OUT <= 0;  //73 / 125 = 0
    16'b01001001_01111110 : OUT <= 0;  //73 / 126 = 0
    16'b01001001_01111111 : OUT <= 0;  //73 / 127 = 0
    16'b01001001_10000000 : OUT <= 0;  //73 / 128 = 0
    16'b01001001_10000001 : OUT <= 0;  //73 / 129 = 0
    16'b01001001_10000010 : OUT <= 0;  //73 / 130 = 0
    16'b01001001_10000011 : OUT <= 0;  //73 / 131 = 0
    16'b01001001_10000100 : OUT <= 0;  //73 / 132 = 0
    16'b01001001_10000101 : OUT <= 0;  //73 / 133 = 0
    16'b01001001_10000110 : OUT <= 0;  //73 / 134 = 0
    16'b01001001_10000111 : OUT <= 0;  //73 / 135 = 0
    16'b01001001_10001000 : OUT <= 0;  //73 / 136 = 0
    16'b01001001_10001001 : OUT <= 0;  //73 / 137 = 0
    16'b01001001_10001010 : OUT <= 0;  //73 / 138 = 0
    16'b01001001_10001011 : OUT <= 0;  //73 / 139 = 0
    16'b01001001_10001100 : OUT <= 0;  //73 / 140 = 0
    16'b01001001_10001101 : OUT <= 0;  //73 / 141 = 0
    16'b01001001_10001110 : OUT <= 0;  //73 / 142 = 0
    16'b01001001_10001111 : OUT <= 0;  //73 / 143 = 0
    16'b01001001_10010000 : OUT <= 0;  //73 / 144 = 0
    16'b01001001_10010001 : OUT <= 0;  //73 / 145 = 0
    16'b01001001_10010010 : OUT <= 0;  //73 / 146 = 0
    16'b01001001_10010011 : OUT <= 0;  //73 / 147 = 0
    16'b01001001_10010100 : OUT <= 0;  //73 / 148 = 0
    16'b01001001_10010101 : OUT <= 0;  //73 / 149 = 0
    16'b01001001_10010110 : OUT <= 0;  //73 / 150 = 0
    16'b01001001_10010111 : OUT <= 0;  //73 / 151 = 0
    16'b01001001_10011000 : OUT <= 0;  //73 / 152 = 0
    16'b01001001_10011001 : OUT <= 0;  //73 / 153 = 0
    16'b01001001_10011010 : OUT <= 0;  //73 / 154 = 0
    16'b01001001_10011011 : OUT <= 0;  //73 / 155 = 0
    16'b01001001_10011100 : OUT <= 0;  //73 / 156 = 0
    16'b01001001_10011101 : OUT <= 0;  //73 / 157 = 0
    16'b01001001_10011110 : OUT <= 0;  //73 / 158 = 0
    16'b01001001_10011111 : OUT <= 0;  //73 / 159 = 0
    16'b01001001_10100000 : OUT <= 0;  //73 / 160 = 0
    16'b01001001_10100001 : OUT <= 0;  //73 / 161 = 0
    16'b01001001_10100010 : OUT <= 0;  //73 / 162 = 0
    16'b01001001_10100011 : OUT <= 0;  //73 / 163 = 0
    16'b01001001_10100100 : OUT <= 0;  //73 / 164 = 0
    16'b01001001_10100101 : OUT <= 0;  //73 / 165 = 0
    16'b01001001_10100110 : OUT <= 0;  //73 / 166 = 0
    16'b01001001_10100111 : OUT <= 0;  //73 / 167 = 0
    16'b01001001_10101000 : OUT <= 0;  //73 / 168 = 0
    16'b01001001_10101001 : OUT <= 0;  //73 / 169 = 0
    16'b01001001_10101010 : OUT <= 0;  //73 / 170 = 0
    16'b01001001_10101011 : OUT <= 0;  //73 / 171 = 0
    16'b01001001_10101100 : OUT <= 0;  //73 / 172 = 0
    16'b01001001_10101101 : OUT <= 0;  //73 / 173 = 0
    16'b01001001_10101110 : OUT <= 0;  //73 / 174 = 0
    16'b01001001_10101111 : OUT <= 0;  //73 / 175 = 0
    16'b01001001_10110000 : OUT <= 0;  //73 / 176 = 0
    16'b01001001_10110001 : OUT <= 0;  //73 / 177 = 0
    16'b01001001_10110010 : OUT <= 0;  //73 / 178 = 0
    16'b01001001_10110011 : OUT <= 0;  //73 / 179 = 0
    16'b01001001_10110100 : OUT <= 0;  //73 / 180 = 0
    16'b01001001_10110101 : OUT <= 0;  //73 / 181 = 0
    16'b01001001_10110110 : OUT <= 0;  //73 / 182 = 0
    16'b01001001_10110111 : OUT <= 0;  //73 / 183 = 0
    16'b01001001_10111000 : OUT <= 0;  //73 / 184 = 0
    16'b01001001_10111001 : OUT <= 0;  //73 / 185 = 0
    16'b01001001_10111010 : OUT <= 0;  //73 / 186 = 0
    16'b01001001_10111011 : OUT <= 0;  //73 / 187 = 0
    16'b01001001_10111100 : OUT <= 0;  //73 / 188 = 0
    16'b01001001_10111101 : OUT <= 0;  //73 / 189 = 0
    16'b01001001_10111110 : OUT <= 0;  //73 / 190 = 0
    16'b01001001_10111111 : OUT <= 0;  //73 / 191 = 0
    16'b01001001_11000000 : OUT <= 0;  //73 / 192 = 0
    16'b01001001_11000001 : OUT <= 0;  //73 / 193 = 0
    16'b01001001_11000010 : OUT <= 0;  //73 / 194 = 0
    16'b01001001_11000011 : OUT <= 0;  //73 / 195 = 0
    16'b01001001_11000100 : OUT <= 0;  //73 / 196 = 0
    16'b01001001_11000101 : OUT <= 0;  //73 / 197 = 0
    16'b01001001_11000110 : OUT <= 0;  //73 / 198 = 0
    16'b01001001_11000111 : OUT <= 0;  //73 / 199 = 0
    16'b01001001_11001000 : OUT <= 0;  //73 / 200 = 0
    16'b01001001_11001001 : OUT <= 0;  //73 / 201 = 0
    16'b01001001_11001010 : OUT <= 0;  //73 / 202 = 0
    16'b01001001_11001011 : OUT <= 0;  //73 / 203 = 0
    16'b01001001_11001100 : OUT <= 0;  //73 / 204 = 0
    16'b01001001_11001101 : OUT <= 0;  //73 / 205 = 0
    16'b01001001_11001110 : OUT <= 0;  //73 / 206 = 0
    16'b01001001_11001111 : OUT <= 0;  //73 / 207 = 0
    16'b01001001_11010000 : OUT <= 0;  //73 / 208 = 0
    16'b01001001_11010001 : OUT <= 0;  //73 / 209 = 0
    16'b01001001_11010010 : OUT <= 0;  //73 / 210 = 0
    16'b01001001_11010011 : OUT <= 0;  //73 / 211 = 0
    16'b01001001_11010100 : OUT <= 0;  //73 / 212 = 0
    16'b01001001_11010101 : OUT <= 0;  //73 / 213 = 0
    16'b01001001_11010110 : OUT <= 0;  //73 / 214 = 0
    16'b01001001_11010111 : OUT <= 0;  //73 / 215 = 0
    16'b01001001_11011000 : OUT <= 0;  //73 / 216 = 0
    16'b01001001_11011001 : OUT <= 0;  //73 / 217 = 0
    16'b01001001_11011010 : OUT <= 0;  //73 / 218 = 0
    16'b01001001_11011011 : OUT <= 0;  //73 / 219 = 0
    16'b01001001_11011100 : OUT <= 0;  //73 / 220 = 0
    16'b01001001_11011101 : OUT <= 0;  //73 / 221 = 0
    16'b01001001_11011110 : OUT <= 0;  //73 / 222 = 0
    16'b01001001_11011111 : OUT <= 0;  //73 / 223 = 0
    16'b01001001_11100000 : OUT <= 0;  //73 / 224 = 0
    16'b01001001_11100001 : OUT <= 0;  //73 / 225 = 0
    16'b01001001_11100010 : OUT <= 0;  //73 / 226 = 0
    16'b01001001_11100011 : OUT <= 0;  //73 / 227 = 0
    16'b01001001_11100100 : OUT <= 0;  //73 / 228 = 0
    16'b01001001_11100101 : OUT <= 0;  //73 / 229 = 0
    16'b01001001_11100110 : OUT <= 0;  //73 / 230 = 0
    16'b01001001_11100111 : OUT <= 0;  //73 / 231 = 0
    16'b01001001_11101000 : OUT <= 0;  //73 / 232 = 0
    16'b01001001_11101001 : OUT <= 0;  //73 / 233 = 0
    16'b01001001_11101010 : OUT <= 0;  //73 / 234 = 0
    16'b01001001_11101011 : OUT <= 0;  //73 / 235 = 0
    16'b01001001_11101100 : OUT <= 0;  //73 / 236 = 0
    16'b01001001_11101101 : OUT <= 0;  //73 / 237 = 0
    16'b01001001_11101110 : OUT <= 0;  //73 / 238 = 0
    16'b01001001_11101111 : OUT <= 0;  //73 / 239 = 0
    16'b01001001_11110000 : OUT <= 0;  //73 / 240 = 0
    16'b01001001_11110001 : OUT <= 0;  //73 / 241 = 0
    16'b01001001_11110010 : OUT <= 0;  //73 / 242 = 0
    16'b01001001_11110011 : OUT <= 0;  //73 / 243 = 0
    16'b01001001_11110100 : OUT <= 0;  //73 / 244 = 0
    16'b01001001_11110101 : OUT <= 0;  //73 / 245 = 0
    16'b01001001_11110110 : OUT <= 0;  //73 / 246 = 0
    16'b01001001_11110111 : OUT <= 0;  //73 / 247 = 0
    16'b01001001_11111000 : OUT <= 0;  //73 / 248 = 0
    16'b01001001_11111001 : OUT <= 0;  //73 / 249 = 0
    16'b01001001_11111010 : OUT <= 0;  //73 / 250 = 0
    16'b01001001_11111011 : OUT <= 0;  //73 / 251 = 0
    16'b01001001_11111100 : OUT <= 0;  //73 / 252 = 0
    16'b01001001_11111101 : OUT <= 0;  //73 / 253 = 0
    16'b01001001_11111110 : OUT <= 0;  //73 / 254 = 0
    16'b01001001_11111111 : OUT <= 0;  //73 / 255 = 0
    16'b01001010_00000000 : OUT <= 0;  //74 / 0 = 0
    16'b01001010_00000001 : OUT <= 74;  //74 / 1 = 74
    16'b01001010_00000010 : OUT <= 37;  //74 / 2 = 37
    16'b01001010_00000011 : OUT <= 24;  //74 / 3 = 24
    16'b01001010_00000100 : OUT <= 18;  //74 / 4 = 18
    16'b01001010_00000101 : OUT <= 14;  //74 / 5 = 14
    16'b01001010_00000110 : OUT <= 12;  //74 / 6 = 12
    16'b01001010_00000111 : OUT <= 10;  //74 / 7 = 10
    16'b01001010_00001000 : OUT <= 9;  //74 / 8 = 9
    16'b01001010_00001001 : OUT <= 8;  //74 / 9 = 8
    16'b01001010_00001010 : OUT <= 7;  //74 / 10 = 7
    16'b01001010_00001011 : OUT <= 6;  //74 / 11 = 6
    16'b01001010_00001100 : OUT <= 6;  //74 / 12 = 6
    16'b01001010_00001101 : OUT <= 5;  //74 / 13 = 5
    16'b01001010_00001110 : OUT <= 5;  //74 / 14 = 5
    16'b01001010_00001111 : OUT <= 4;  //74 / 15 = 4
    16'b01001010_00010000 : OUT <= 4;  //74 / 16 = 4
    16'b01001010_00010001 : OUT <= 4;  //74 / 17 = 4
    16'b01001010_00010010 : OUT <= 4;  //74 / 18 = 4
    16'b01001010_00010011 : OUT <= 3;  //74 / 19 = 3
    16'b01001010_00010100 : OUT <= 3;  //74 / 20 = 3
    16'b01001010_00010101 : OUT <= 3;  //74 / 21 = 3
    16'b01001010_00010110 : OUT <= 3;  //74 / 22 = 3
    16'b01001010_00010111 : OUT <= 3;  //74 / 23 = 3
    16'b01001010_00011000 : OUT <= 3;  //74 / 24 = 3
    16'b01001010_00011001 : OUT <= 2;  //74 / 25 = 2
    16'b01001010_00011010 : OUT <= 2;  //74 / 26 = 2
    16'b01001010_00011011 : OUT <= 2;  //74 / 27 = 2
    16'b01001010_00011100 : OUT <= 2;  //74 / 28 = 2
    16'b01001010_00011101 : OUT <= 2;  //74 / 29 = 2
    16'b01001010_00011110 : OUT <= 2;  //74 / 30 = 2
    16'b01001010_00011111 : OUT <= 2;  //74 / 31 = 2
    16'b01001010_00100000 : OUT <= 2;  //74 / 32 = 2
    16'b01001010_00100001 : OUT <= 2;  //74 / 33 = 2
    16'b01001010_00100010 : OUT <= 2;  //74 / 34 = 2
    16'b01001010_00100011 : OUT <= 2;  //74 / 35 = 2
    16'b01001010_00100100 : OUT <= 2;  //74 / 36 = 2
    16'b01001010_00100101 : OUT <= 2;  //74 / 37 = 2
    16'b01001010_00100110 : OUT <= 1;  //74 / 38 = 1
    16'b01001010_00100111 : OUT <= 1;  //74 / 39 = 1
    16'b01001010_00101000 : OUT <= 1;  //74 / 40 = 1
    16'b01001010_00101001 : OUT <= 1;  //74 / 41 = 1
    16'b01001010_00101010 : OUT <= 1;  //74 / 42 = 1
    16'b01001010_00101011 : OUT <= 1;  //74 / 43 = 1
    16'b01001010_00101100 : OUT <= 1;  //74 / 44 = 1
    16'b01001010_00101101 : OUT <= 1;  //74 / 45 = 1
    16'b01001010_00101110 : OUT <= 1;  //74 / 46 = 1
    16'b01001010_00101111 : OUT <= 1;  //74 / 47 = 1
    16'b01001010_00110000 : OUT <= 1;  //74 / 48 = 1
    16'b01001010_00110001 : OUT <= 1;  //74 / 49 = 1
    16'b01001010_00110010 : OUT <= 1;  //74 / 50 = 1
    16'b01001010_00110011 : OUT <= 1;  //74 / 51 = 1
    16'b01001010_00110100 : OUT <= 1;  //74 / 52 = 1
    16'b01001010_00110101 : OUT <= 1;  //74 / 53 = 1
    16'b01001010_00110110 : OUT <= 1;  //74 / 54 = 1
    16'b01001010_00110111 : OUT <= 1;  //74 / 55 = 1
    16'b01001010_00111000 : OUT <= 1;  //74 / 56 = 1
    16'b01001010_00111001 : OUT <= 1;  //74 / 57 = 1
    16'b01001010_00111010 : OUT <= 1;  //74 / 58 = 1
    16'b01001010_00111011 : OUT <= 1;  //74 / 59 = 1
    16'b01001010_00111100 : OUT <= 1;  //74 / 60 = 1
    16'b01001010_00111101 : OUT <= 1;  //74 / 61 = 1
    16'b01001010_00111110 : OUT <= 1;  //74 / 62 = 1
    16'b01001010_00111111 : OUT <= 1;  //74 / 63 = 1
    16'b01001010_01000000 : OUT <= 1;  //74 / 64 = 1
    16'b01001010_01000001 : OUT <= 1;  //74 / 65 = 1
    16'b01001010_01000010 : OUT <= 1;  //74 / 66 = 1
    16'b01001010_01000011 : OUT <= 1;  //74 / 67 = 1
    16'b01001010_01000100 : OUT <= 1;  //74 / 68 = 1
    16'b01001010_01000101 : OUT <= 1;  //74 / 69 = 1
    16'b01001010_01000110 : OUT <= 1;  //74 / 70 = 1
    16'b01001010_01000111 : OUT <= 1;  //74 / 71 = 1
    16'b01001010_01001000 : OUT <= 1;  //74 / 72 = 1
    16'b01001010_01001001 : OUT <= 1;  //74 / 73 = 1
    16'b01001010_01001010 : OUT <= 1;  //74 / 74 = 1
    16'b01001010_01001011 : OUT <= 0;  //74 / 75 = 0
    16'b01001010_01001100 : OUT <= 0;  //74 / 76 = 0
    16'b01001010_01001101 : OUT <= 0;  //74 / 77 = 0
    16'b01001010_01001110 : OUT <= 0;  //74 / 78 = 0
    16'b01001010_01001111 : OUT <= 0;  //74 / 79 = 0
    16'b01001010_01010000 : OUT <= 0;  //74 / 80 = 0
    16'b01001010_01010001 : OUT <= 0;  //74 / 81 = 0
    16'b01001010_01010010 : OUT <= 0;  //74 / 82 = 0
    16'b01001010_01010011 : OUT <= 0;  //74 / 83 = 0
    16'b01001010_01010100 : OUT <= 0;  //74 / 84 = 0
    16'b01001010_01010101 : OUT <= 0;  //74 / 85 = 0
    16'b01001010_01010110 : OUT <= 0;  //74 / 86 = 0
    16'b01001010_01010111 : OUT <= 0;  //74 / 87 = 0
    16'b01001010_01011000 : OUT <= 0;  //74 / 88 = 0
    16'b01001010_01011001 : OUT <= 0;  //74 / 89 = 0
    16'b01001010_01011010 : OUT <= 0;  //74 / 90 = 0
    16'b01001010_01011011 : OUT <= 0;  //74 / 91 = 0
    16'b01001010_01011100 : OUT <= 0;  //74 / 92 = 0
    16'b01001010_01011101 : OUT <= 0;  //74 / 93 = 0
    16'b01001010_01011110 : OUT <= 0;  //74 / 94 = 0
    16'b01001010_01011111 : OUT <= 0;  //74 / 95 = 0
    16'b01001010_01100000 : OUT <= 0;  //74 / 96 = 0
    16'b01001010_01100001 : OUT <= 0;  //74 / 97 = 0
    16'b01001010_01100010 : OUT <= 0;  //74 / 98 = 0
    16'b01001010_01100011 : OUT <= 0;  //74 / 99 = 0
    16'b01001010_01100100 : OUT <= 0;  //74 / 100 = 0
    16'b01001010_01100101 : OUT <= 0;  //74 / 101 = 0
    16'b01001010_01100110 : OUT <= 0;  //74 / 102 = 0
    16'b01001010_01100111 : OUT <= 0;  //74 / 103 = 0
    16'b01001010_01101000 : OUT <= 0;  //74 / 104 = 0
    16'b01001010_01101001 : OUT <= 0;  //74 / 105 = 0
    16'b01001010_01101010 : OUT <= 0;  //74 / 106 = 0
    16'b01001010_01101011 : OUT <= 0;  //74 / 107 = 0
    16'b01001010_01101100 : OUT <= 0;  //74 / 108 = 0
    16'b01001010_01101101 : OUT <= 0;  //74 / 109 = 0
    16'b01001010_01101110 : OUT <= 0;  //74 / 110 = 0
    16'b01001010_01101111 : OUT <= 0;  //74 / 111 = 0
    16'b01001010_01110000 : OUT <= 0;  //74 / 112 = 0
    16'b01001010_01110001 : OUT <= 0;  //74 / 113 = 0
    16'b01001010_01110010 : OUT <= 0;  //74 / 114 = 0
    16'b01001010_01110011 : OUT <= 0;  //74 / 115 = 0
    16'b01001010_01110100 : OUT <= 0;  //74 / 116 = 0
    16'b01001010_01110101 : OUT <= 0;  //74 / 117 = 0
    16'b01001010_01110110 : OUT <= 0;  //74 / 118 = 0
    16'b01001010_01110111 : OUT <= 0;  //74 / 119 = 0
    16'b01001010_01111000 : OUT <= 0;  //74 / 120 = 0
    16'b01001010_01111001 : OUT <= 0;  //74 / 121 = 0
    16'b01001010_01111010 : OUT <= 0;  //74 / 122 = 0
    16'b01001010_01111011 : OUT <= 0;  //74 / 123 = 0
    16'b01001010_01111100 : OUT <= 0;  //74 / 124 = 0
    16'b01001010_01111101 : OUT <= 0;  //74 / 125 = 0
    16'b01001010_01111110 : OUT <= 0;  //74 / 126 = 0
    16'b01001010_01111111 : OUT <= 0;  //74 / 127 = 0
    16'b01001010_10000000 : OUT <= 0;  //74 / 128 = 0
    16'b01001010_10000001 : OUT <= 0;  //74 / 129 = 0
    16'b01001010_10000010 : OUT <= 0;  //74 / 130 = 0
    16'b01001010_10000011 : OUT <= 0;  //74 / 131 = 0
    16'b01001010_10000100 : OUT <= 0;  //74 / 132 = 0
    16'b01001010_10000101 : OUT <= 0;  //74 / 133 = 0
    16'b01001010_10000110 : OUT <= 0;  //74 / 134 = 0
    16'b01001010_10000111 : OUT <= 0;  //74 / 135 = 0
    16'b01001010_10001000 : OUT <= 0;  //74 / 136 = 0
    16'b01001010_10001001 : OUT <= 0;  //74 / 137 = 0
    16'b01001010_10001010 : OUT <= 0;  //74 / 138 = 0
    16'b01001010_10001011 : OUT <= 0;  //74 / 139 = 0
    16'b01001010_10001100 : OUT <= 0;  //74 / 140 = 0
    16'b01001010_10001101 : OUT <= 0;  //74 / 141 = 0
    16'b01001010_10001110 : OUT <= 0;  //74 / 142 = 0
    16'b01001010_10001111 : OUT <= 0;  //74 / 143 = 0
    16'b01001010_10010000 : OUT <= 0;  //74 / 144 = 0
    16'b01001010_10010001 : OUT <= 0;  //74 / 145 = 0
    16'b01001010_10010010 : OUT <= 0;  //74 / 146 = 0
    16'b01001010_10010011 : OUT <= 0;  //74 / 147 = 0
    16'b01001010_10010100 : OUT <= 0;  //74 / 148 = 0
    16'b01001010_10010101 : OUT <= 0;  //74 / 149 = 0
    16'b01001010_10010110 : OUT <= 0;  //74 / 150 = 0
    16'b01001010_10010111 : OUT <= 0;  //74 / 151 = 0
    16'b01001010_10011000 : OUT <= 0;  //74 / 152 = 0
    16'b01001010_10011001 : OUT <= 0;  //74 / 153 = 0
    16'b01001010_10011010 : OUT <= 0;  //74 / 154 = 0
    16'b01001010_10011011 : OUT <= 0;  //74 / 155 = 0
    16'b01001010_10011100 : OUT <= 0;  //74 / 156 = 0
    16'b01001010_10011101 : OUT <= 0;  //74 / 157 = 0
    16'b01001010_10011110 : OUT <= 0;  //74 / 158 = 0
    16'b01001010_10011111 : OUT <= 0;  //74 / 159 = 0
    16'b01001010_10100000 : OUT <= 0;  //74 / 160 = 0
    16'b01001010_10100001 : OUT <= 0;  //74 / 161 = 0
    16'b01001010_10100010 : OUT <= 0;  //74 / 162 = 0
    16'b01001010_10100011 : OUT <= 0;  //74 / 163 = 0
    16'b01001010_10100100 : OUT <= 0;  //74 / 164 = 0
    16'b01001010_10100101 : OUT <= 0;  //74 / 165 = 0
    16'b01001010_10100110 : OUT <= 0;  //74 / 166 = 0
    16'b01001010_10100111 : OUT <= 0;  //74 / 167 = 0
    16'b01001010_10101000 : OUT <= 0;  //74 / 168 = 0
    16'b01001010_10101001 : OUT <= 0;  //74 / 169 = 0
    16'b01001010_10101010 : OUT <= 0;  //74 / 170 = 0
    16'b01001010_10101011 : OUT <= 0;  //74 / 171 = 0
    16'b01001010_10101100 : OUT <= 0;  //74 / 172 = 0
    16'b01001010_10101101 : OUT <= 0;  //74 / 173 = 0
    16'b01001010_10101110 : OUT <= 0;  //74 / 174 = 0
    16'b01001010_10101111 : OUT <= 0;  //74 / 175 = 0
    16'b01001010_10110000 : OUT <= 0;  //74 / 176 = 0
    16'b01001010_10110001 : OUT <= 0;  //74 / 177 = 0
    16'b01001010_10110010 : OUT <= 0;  //74 / 178 = 0
    16'b01001010_10110011 : OUT <= 0;  //74 / 179 = 0
    16'b01001010_10110100 : OUT <= 0;  //74 / 180 = 0
    16'b01001010_10110101 : OUT <= 0;  //74 / 181 = 0
    16'b01001010_10110110 : OUT <= 0;  //74 / 182 = 0
    16'b01001010_10110111 : OUT <= 0;  //74 / 183 = 0
    16'b01001010_10111000 : OUT <= 0;  //74 / 184 = 0
    16'b01001010_10111001 : OUT <= 0;  //74 / 185 = 0
    16'b01001010_10111010 : OUT <= 0;  //74 / 186 = 0
    16'b01001010_10111011 : OUT <= 0;  //74 / 187 = 0
    16'b01001010_10111100 : OUT <= 0;  //74 / 188 = 0
    16'b01001010_10111101 : OUT <= 0;  //74 / 189 = 0
    16'b01001010_10111110 : OUT <= 0;  //74 / 190 = 0
    16'b01001010_10111111 : OUT <= 0;  //74 / 191 = 0
    16'b01001010_11000000 : OUT <= 0;  //74 / 192 = 0
    16'b01001010_11000001 : OUT <= 0;  //74 / 193 = 0
    16'b01001010_11000010 : OUT <= 0;  //74 / 194 = 0
    16'b01001010_11000011 : OUT <= 0;  //74 / 195 = 0
    16'b01001010_11000100 : OUT <= 0;  //74 / 196 = 0
    16'b01001010_11000101 : OUT <= 0;  //74 / 197 = 0
    16'b01001010_11000110 : OUT <= 0;  //74 / 198 = 0
    16'b01001010_11000111 : OUT <= 0;  //74 / 199 = 0
    16'b01001010_11001000 : OUT <= 0;  //74 / 200 = 0
    16'b01001010_11001001 : OUT <= 0;  //74 / 201 = 0
    16'b01001010_11001010 : OUT <= 0;  //74 / 202 = 0
    16'b01001010_11001011 : OUT <= 0;  //74 / 203 = 0
    16'b01001010_11001100 : OUT <= 0;  //74 / 204 = 0
    16'b01001010_11001101 : OUT <= 0;  //74 / 205 = 0
    16'b01001010_11001110 : OUT <= 0;  //74 / 206 = 0
    16'b01001010_11001111 : OUT <= 0;  //74 / 207 = 0
    16'b01001010_11010000 : OUT <= 0;  //74 / 208 = 0
    16'b01001010_11010001 : OUT <= 0;  //74 / 209 = 0
    16'b01001010_11010010 : OUT <= 0;  //74 / 210 = 0
    16'b01001010_11010011 : OUT <= 0;  //74 / 211 = 0
    16'b01001010_11010100 : OUT <= 0;  //74 / 212 = 0
    16'b01001010_11010101 : OUT <= 0;  //74 / 213 = 0
    16'b01001010_11010110 : OUT <= 0;  //74 / 214 = 0
    16'b01001010_11010111 : OUT <= 0;  //74 / 215 = 0
    16'b01001010_11011000 : OUT <= 0;  //74 / 216 = 0
    16'b01001010_11011001 : OUT <= 0;  //74 / 217 = 0
    16'b01001010_11011010 : OUT <= 0;  //74 / 218 = 0
    16'b01001010_11011011 : OUT <= 0;  //74 / 219 = 0
    16'b01001010_11011100 : OUT <= 0;  //74 / 220 = 0
    16'b01001010_11011101 : OUT <= 0;  //74 / 221 = 0
    16'b01001010_11011110 : OUT <= 0;  //74 / 222 = 0
    16'b01001010_11011111 : OUT <= 0;  //74 / 223 = 0
    16'b01001010_11100000 : OUT <= 0;  //74 / 224 = 0
    16'b01001010_11100001 : OUT <= 0;  //74 / 225 = 0
    16'b01001010_11100010 : OUT <= 0;  //74 / 226 = 0
    16'b01001010_11100011 : OUT <= 0;  //74 / 227 = 0
    16'b01001010_11100100 : OUT <= 0;  //74 / 228 = 0
    16'b01001010_11100101 : OUT <= 0;  //74 / 229 = 0
    16'b01001010_11100110 : OUT <= 0;  //74 / 230 = 0
    16'b01001010_11100111 : OUT <= 0;  //74 / 231 = 0
    16'b01001010_11101000 : OUT <= 0;  //74 / 232 = 0
    16'b01001010_11101001 : OUT <= 0;  //74 / 233 = 0
    16'b01001010_11101010 : OUT <= 0;  //74 / 234 = 0
    16'b01001010_11101011 : OUT <= 0;  //74 / 235 = 0
    16'b01001010_11101100 : OUT <= 0;  //74 / 236 = 0
    16'b01001010_11101101 : OUT <= 0;  //74 / 237 = 0
    16'b01001010_11101110 : OUT <= 0;  //74 / 238 = 0
    16'b01001010_11101111 : OUT <= 0;  //74 / 239 = 0
    16'b01001010_11110000 : OUT <= 0;  //74 / 240 = 0
    16'b01001010_11110001 : OUT <= 0;  //74 / 241 = 0
    16'b01001010_11110010 : OUT <= 0;  //74 / 242 = 0
    16'b01001010_11110011 : OUT <= 0;  //74 / 243 = 0
    16'b01001010_11110100 : OUT <= 0;  //74 / 244 = 0
    16'b01001010_11110101 : OUT <= 0;  //74 / 245 = 0
    16'b01001010_11110110 : OUT <= 0;  //74 / 246 = 0
    16'b01001010_11110111 : OUT <= 0;  //74 / 247 = 0
    16'b01001010_11111000 : OUT <= 0;  //74 / 248 = 0
    16'b01001010_11111001 : OUT <= 0;  //74 / 249 = 0
    16'b01001010_11111010 : OUT <= 0;  //74 / 250 = 0
    16'b01001010_11111011 : OUT <= 0;  //74 / 251 = 0
    16'b01001010_11111100 : OUT <= 0;  //74 / 252 = 0
    16'b01001010_11111101 : OUT <= 0;  //74 / 253 = 0
    16'b01001010_11111110 : OUT <= 0;  //74 / 254 = 0
    16'b01001010_11111111 : OUT <= 0;  //74 / 255 = 0
    16'b01001011_00000000 : OUT <= 0;  //75 / 0 = 0
    16'b01001011_00000001 : OUT <= 75;  //75 / 1 = 75
    16'b01001011_00000010 : OUT <= 37;  //75 / 2 = 37
    16'b01001011_00000011 : OUT <= 25;  //75 / 3 = 25
    16'b01001011_00000100 : OUT <= 18;  //75 / 4 = 18
    16'b01001011_00000101 : OUT <= 15;  //75 / 5 = 15
    16'b01001011_00000110 : OUT <= 12;  //75 / 6 = 12
    16'b01001011_00000111 : OUT <= 10;  //75 / 7 = 10
    16'b01001011_00001000 : OUT <= 9;  //75 / 8 = 9
    16'b01001011_00001001 : OUT <= 8;  //75 / 9 = 8
    16'b01001011_00001010 : OUT <= 7;  //75 / 10 = 7
    16'b01001011_00001011 : OUT <= 6;  //75 / 11 = 6
    16'b01001011_00001100 : OUT <= 6;  //75 / 12 = 6
    16'b01001011_00001101 : OUT <= 5;  //75 / 13 = 5
    16'b01001011_00001110 : OUT <= 5;  //75 / 14 = 5
    16'b01001011_00001111 : OUT <= 5;  //75 / 15 = 5
    16'b01001011_00010000 : OUT <= 4;  //75 / 16 = 4
    16'b01001011_00010001 : OUT <= 4;  //75 / 17 = 4
    16'b01001011_00010010 : OUT <= 4;  //75 / 18 = 4
    16'b01001011_00010011 : OUT <= 3;  //75 / 19 = 3
    16'b01001011_00010100 : OUT <= 3;  //75 / 20 = 3
    16'b01001011_00010101 : OUT <= 3;  //75 / 21 = 3
    16'b01001011_00010110 : OUT <= 3;  //75 / 22 = 3
    16'b01001011_00010111 : OUT <= 3;  //75 / 23 = 3
    16'b01001011_00011000 : OUT <= 3;  //75 / 24 = 3
    16'b01001011_00011001 : OUT <= 3;  //75 / 25 = 3
    16'b01001011_00011010 : OUT <= 2;  //75 / 26 = 2
    16'b01001011_00011011 : OUT <= 2;  //75 / 27 = 2
    16'b01001011_00011100 : OUT <= 2;  //75 / 28 = 2
    16'b01001011_00011101 : OUT <= 2;  //75 / 29 = 2
    16'b01001011_00011110 : OUT <= 2;  //75 / 30 = 2
    16'b01001011_00011111 : OUT <= 2;  //75 / 31 = 2
    16'b01001011_00100000 : OUT <= 2;  //75 / 32 = 2
    16'b01001011_00100001 : OUT <= 2;  //75 / 33 = 2
    16'b01001011_00100010 : OUT <= 2;  //75 / 34 = 2
    16'b01001011_00100011 : OUT <= 2;  //75 / 35 = 2
    16'b01001011_00100100 : OUT <= 2;  //75 / 36 = 2
    16'b01001011_00100101 : OUT <= 2;  //75 / 37 = 2
    16'b01001011_00100110 : OUT <= 1;  //75 / 38 = 1
    16'b01001011_00100111 : OUT <= 1;  //75 / 39 = 1
    16'b01001011_00101000 : OUT <= 1;  //75 / 40 = 1
    16'b01001011_00101001 : OUT <= 1;  //75 / 41 = 1
    16'b01001011_00101010 : OUT <= 1;  //75 / 42 = 1
    16'b01001011_00101011 : OUT <= 1;  //75 / 43 = 1
    16'b01001011_00101100 : OUT <= 1;  //75 / 44 = 1
    16'b01001011_00101101 : OUT <= 1;  //75 / 45 = 1
    16'b01001011_00101110 : OUT <= 1;  //75 / 46 = 1
    16'b01001011_00101111 : OUT <= 1;  //75 / 47 = 1
    16'b01001011_00110000 : OUT <= 1;  //75 / 48 = 1
    16'b01001011_00110001 : OUT <= 1;  //75 / 49 = 1
    16'b01001011_00110010 : OUT <= 1;  //75 / 50 = 1
    16'b01001011_00110011 : OUT <= 1;  //75 / 51 = 1
    16'b01001011_00110100 : OUT <= 1;  //75 / 52 = 1
    16'b01001011_00110101 : OUT <= 1;  //75 / 53 = 1
    16'b01001011_00110110 : OUT <= 1;  //75 / 54 = 1
    16'b01001011_00110111 : OUT <= 1;  //75 / 55 = 1
    16'b01001011_00111000 : OUT <= 1;  //75 / 56 = 1
    16'b01001011_00111001 : OUT <= 1;  //75 / 57 = 1
    16'b01001011_00111010 : OUT <= 1;  //75 / 58 = 1
    16'b01001011_00111011 : OUT <= 1;  //75 / 59 = 1
    16'b01001011_00111100 : OUT <= 1;  //75 / 60 = 1
    16'b01001011_00111101 : OUT <= 1;  //75 / 61 = 1
    16'b01001011_00111110 : OUT <= 1;  //75 / 62 = 1
    16'b01001011_00111111 : OUT <= 1;  //75 / 63 = 1
    16'b01001011_01000000 : OUT <= 1;  //75 / 64 = 1
    16'b01001011_01000001 : OUT <= 1;  //75 / 65 = 1
    16'b01001011_01000010 : OUT <= 1;  //75 / 66 = 1
    16'b01001011_01000011 : OUT <= 1;  //75 / 67 = 1
    16'b01001011_01000100 : OUT <= 1;  //75 / 68 = 1
    16'b01001011_01000101 : OUT <= 1;  //75 / 69 = 1
    16'b01001011_01000110 : OUT <= 1;  //75 / 70 = 1
    16'b01001011_01000111 : OUT <= 1;  //75 / 71 = 1
    16'b01001011_01001000 : OUT <= 1;  //75 / 72 = 1
    16'b01001011_01001001 : OUT <= 1;  //75 / 73 = 1
    16'b01001011_01001010 : OUT <= 1;  //75 / 74 = 1
    16'b01001011_01001011 : OUT <= 1;  //75 / 75 = 1
    16'b01001011_01001100 : OUT <= 0;  //75 / 76 = 0
    16'b01001011_01001101 : OUT <= 0;  //75 / 77 = 0
    16'b01001011_01001110 : OUT <= 0;  //75 / 78 = 0
    16'b01001011_01001111 : OUT <= 0;  //75 / 79 = 0
    16'b01001011_01010000 : OUT <= 0;  //75 / 80 = 0
    16'b01001011_01010001 : OUT <= 0;  //75 / 81 = 0
    16'b01001011_01010010 : OUT <= 0;  //75 / 82 = 0
    16'b01001011_01010011 : OUT <= 0;  //75 / 83 = 0
    16'b01001011_01010100 : OUT <= 0;  //75 / 84 = 0
    16'b01001011_01010101 : OUT <= 0;  //75 / 85 = 0
    16'b01001011_01010110 : OUT <= 0;  //75 / 86 = 0
    16'b01001011_01010111 : OUT <= 0;  //75 / 87 = 0
    16'b01001011_01011000 : OUT <= 0;  //75 / 88 = 0
    16'b01001011_01011001 : OUT <= 0;  //75 / 89 = 0
    16'b01001011_01011010 : OUT <= 0;  //75 / 90 = 0
    16'b01001011_01011011 : OUT <= 0;  //75 / 91 = 0
    16'b01001011_01011100 : OUT <= 0;  //75 / 92 = 0
    16'b01001011_01011101 : OUT <= 0;  //75 / 93 = 0
    16'b01001011_01011110 : OUT <= 0;  //75 / 94 = 0
    16'b01001011_01011111 : OUT <= 0;  //75 / 95 = 0
    16'b01001011_01100000 : OUT <= 0;  //75 / 96 = 0
    16'b01001011_01100001 : OUT <= 0;  //75 / 97 = 0
    16'b01001011_01100010 : OUT <= 0;  //75 / 98 = 0
    16'b01001011_01100011 : OUT <= 0;  //75 / 99 = 0
    16'b01001011_01100100 : OUT <= 0;  //75 / 100 = 0
    16'b01001011_01100101 : OUT <= 0;  //75 / 101 = 0
    16'b01001011_01100110 : OUT <= 0;  //75 / 102 = 0
    16'b01001011_01100111 : OUT <= 0;  //75 / 103 = 0
    16'b01001011_01101000 : OUT <= 0;  //75 / 104 = 0
    16'b01001011_01101001 : OUT <= 0;  //75 / 105 = 0
    16'b01001011_01101010 : OUT <= 0;  //75 / 106 = 0
    16'b01001011_01101011 : OUT <= 0;  //75 / 107 = 0
    16'b01001011_01101100 : OUT <= 0;  //75 / 108 = 0
    16'b01001011_01101101 : OUT <= 0;  //75 / 109 = 0
    16'b01001011_01101110 : OUT <= 0;  //75 / 110 = 0
    16'b01001011_01101111 : OUT <= 0;  //75 / 111 = 0
    16'b01001011_01110000 : OUT <= 0;  //75 / 112 = 0
    16'b01001011_01110001 : OUT <= 0;  //75 / 113 = 0
    16'b01001011_01110010 : OUT <= 0;  //75 / 114 = 0
    16'b01001011_01110011 : OUT <= 0;  //75 / 115 = 0
    16'b01001011_01110100 : OUT <= 0;  //75 / 116 = 0
    16'b01001011_01110101 : OUT <= 0;  //75 / 117 = 0
    16'b01001011_01110110 : OUT <= 0;  //75 / 118 = 0
    16'b01001011_01110111 : OUT <= 0;  //75 / 119 = 0
    16'b01001011_01111000 : OUT <= 0;  //75 / 120 = 0
    16'b01001011_01111001 : OUT <= 0;  //75 / 121 = 0
    16'b01001011_01111010 : OUT <= 0;  //75 / 122 = 0
    16'b01001011_01111011 : OUT <= 0;  //75 / 123 = 0
    16'b01001011_01111100 : OUT <= 0;  //75 / 124 = 0
    16'b01001011_01111101 : OUT <= 0;  //75 / 125 = 0
    16'b01001011_01111110 : OUT <= 0;  //75 / 126 = 0
    16'b01001011_01111111 : OUT <= 0;  //75 / 127 = 0
    16'b01001011_10000000 : OUT <= 0;  //75 / 128 = 0
    16'b01001011_10000001 : OUT <= 0;  //75 / 129 = 0
    16'b01001011_10000010 : OUT <= 0;  //75 / 130 = 0
    16'b01001011_10000011 : OUT <= 0;  //75 / 131 = 0
    16'b01001011_10000100 : OUT <= 0;  //75 / 132 = 0
    16'b01001011_10000101 : OUT <= 0;  //75 / 133 = 0
    16'b01001011_10000110 : OUT <= 0;  //75 / 134 = 0
    16'b01001011_10000111 : OUT <= 0;  //75 / 135 = 0
    16'b01001011_10001000 : OUT <= 0;  //75 / 136 = 0
    16'b01001011_10001001 : OUT <= 0;  //75 / 137 = 0
    16'b01001011_10001010 : OUT <= 0;  //75 / 138 = 0
    16'b01001011_10001011 : OUT <= 0;  //75 / 139 = 0
    16'b01001011_10001100 : OUT <= 0;  //75 / 140 = 0
    16'b01001011_10001101 : OUT <= 0;  //75 / 141 = 0
    16'b01001011_10001110 : OUT <= 0;  //75 / 142 = 0
    16'b01001011_10001111 : OUT <= 0;  //75 / 143 = 0
    16'b01001011_10010000 : OUT <= 0;  //75 / 144 = 0
    16'b01001011_10010001 : OUT <= 0;  //75 / 145 = 0
    16'b01001011_10010010 : OUT <= 0;  //75 / 146 = 0
    16'b01001011_10010011 : OUT <= 0;  //75 / 147 = 0
    16'b01001011_10010100 : OUT <= 0;  //75 / 148 = 0
    16'b01001011_10010101 : OUT <= 0;  //75 / 149 = 0
    16'b01001011_10010110 : OUT <= 0;  //75 / 150 = 0
    16'b01001011_10010111 : OUT <= 0;  //75 / 151 = 0
    16'b01001011_10011000 : OUT <= 0;  //75 / 152 = 0
    16'b01001011_10011001 : OUT <= 0;  //75 / 153 = 0
    16'b01001011_10011010 : OUT <= 0;  //75 / 154 = 0
    16'b01001011_10011011 : OUT <= 0;  //75 / 155 = 0
    16'b01001011_10011100 : OUT <= 0;  //75 / 156 = 0
    16'b01001011_10011101 : OUT <= 0;  //75 / 157 = 0
    16'b01001011_10011110 : OUT <= 0;  //75 / 158 = 0
    16'b01001011_10011111 : OUT <= 0;  //75 / 159 = 0
    16'b01001011_10100000 : OUT <= 0;  //75 / 160 = 0
    16'b01001011_10100001 : OUT <= 0;  //75 / 161 = 0
    16'b01001011_10100010 : OUT <= 0;  //75 / 162 = 0
    16'b01001011_10100011 : OUT <= 0;  //75 / 163 = 0
    16'b01001011_10100100 : OUT <= 0;  //75 / 164 = 0
    16'b01001011_10100101 : OUT <= 0;  //75 / 165 = 0
    16'b01001011_10100110 : OUT <= 0;  //75 / 166 = 0
    16'b01001011_10100111 : OUT <= 0;  //75 / 167 = 0
    16'b01001011_10101000 : OUT <= 0;  //75 / 168 = 0
    16'b01001011_10101001 : OUT <= 0;  //75 / 169 = 0
    16'b01001011_10101010 : OUT <= 0;  //75 / 170 = 0
    16'b01001011_10101011 : OUT <= 0;  //75 / 171 = 0
    16'b01001011_10101100 : OUT <= 0;  //75 / 172 = 0
    16'b01001011_10101101 : OUT <= 0;  //75 / 173 = 0
    16'b01001011_10101110 : OUT <= 0;  //75 / 174 = 0
    16'b01001011_10101111 : OUT <= 0;  //75 / 175 = 0
    16'b01001011_10110000 : OUT <= 0;  //75 / 176 = 0
    16'b01001011_10110001 : OUT <= 0;  //75 / 177 = 0
    16'b01001011_10110010 : OUT <= 0;  //75 / 178 = 0
    16'b01001011_10110011 : OUT <= 0;  //75 / 179 = 0
    16'b01001011_10110100 : OUT <= 0;  //75 / 180 = 0
    16'b01001011_10110101 : OUT <= 0;  //75 / 181 = 0
    16'b01001011_10110110 : OUT <= 0;  //75 / 182 = 0
    16'b01001011_10110111 : OUT <= 0;  //75 / 183 = 0
    16'b01001011_10111000 : OUT <= 0;  //75 / 184 = 0
    16'b01001011_10111001 : OUT <= 0;  //75 / 185 = 0
    16'b01001011_10111010 : OUT <= 0;  //75 / 186 = 0
    16'b01001011_10111011 : OUT <= 0;  //75 / 187 = 0
    16'b01001011_10111100 : OUT <= 0;  //75 / 188 = 0
    16'b01001011_10111101 : OUT <= 0;  //75 / 189 = 0
    16'b01001011_10111110 : OUT <= 0;  //75 / 190 = 0
    16'b01001011_10111111 : OUT <= 0;  //75 / 191 = 0
    16'b01001011_11000000 : OUT <= 0;  //75 / 192 = 0
    16'b01001011_11000001 : OUT <= 0;  //75 / 193 = 0
    16'b01001011_11000010 : OUT <= 0;  //75 / 194 = 0
    16'b01001011_11000011 : OUT <= 0;  //75 / 195 = 0
    16'b01001011_11000100 : OUT <= 0;  //75 / 196 = 0
    16'b01001011_11000101 : OUT <= 0;  //75 / 197 = 0
    16'b01001011_11000110 : OUT <= 0;  //75 / 198 = 0
    16'b01001011_11000111 : OUT <= 0;  //75 / 199 = 0
    16'b01001011_11001000 : OUT <= 0;  //75 / 200 = 0
    16'b01001011_11001001 : OUT <= 0;  //75 / 201 = 0
    16'b01001011_11001010 : OUT <= 0;  //75 / 202 = 0
    16'b01001011_11001011 : OUT <= 0;  //75 / 203 = 0
    16'b01001011_11001100 : OUT <= 0;  //75 / 204 = 0
    16'b01001011_11001101 : OUT <= 0;  //75 / 205 = 0
    16'b01001011_11001110 : OUT <= 0;  //75 / 206 = 0
    16'b01001011_11001111 : OUT <= 0;  //75 / 207 = 0
    16'b01001011_11010000 : OUT <= 0;  //75 / 208 = 0
    16'b01001011_11010001 : OUT <= 0;  //75 / 209 = 0
    16'b01001011_11010010 : OUT <= 0;  //75 / 210 = 0
    16'b01001011_11010011 : OUT <= 0;  //75 / 211 = 0
    16'b01001011_11010100 : OUT <= 0;  //75 / 212 = 0
    16'b01001011_11010101 : OUT <= 0;  //75 / 213 = 0
    16'b01001011_11010110 : OUT <= 0;  //75 / 214 = 0
    16'b01001011_11010111 : OUT <= 0;  //75 / 215 = 0
    16'b01001011_11011000 : OUT <= 0;  //75 / 216 = 0
    16'b01001011_11011001 : OUT <= 0;  //75 / 217 = 0
    16'b01001011_11011010 : OUT <= 0;  //75 / 218 = 0
    16'b01001011_11011011 : OUT <= 0;  //75 / 219 = 0
    16'b01001011_11011100 : OUT <= 0;  //75 / 220 = 0
    16'b01001011_11011101 : OUT <= 0;  //75 / 221 = 0
    16'b01001011_11011110 : OUT <= 0;  //75 / 222 = 0
    16'b01001011_11011111 : OUT <= 0;  //75 / 223 = 0
    16'b01001011_11100000 : OUT <= 0;  //75 / 224 = 0
    16'b01001011_11100001 : OUT <= 0;  //75 / 225 = 0
    16'b01001011_11100010 : OUT <= 0;  //75 / 226 = 0
    16'b01001011_11100011 : OUT <= 0;  //75 / 227 = 0
    16'b01001011_11100100 : OUT <= 0;  //75 / 228 = 0
    16'b01001011_11100101 : OUT <= 0;  //75 / 229 = 0
    16'b01001011_11100110 : OUT <= 0;  //75 / 230 = 0
    16'b01001011_11100111 : OUT <= 0;  //75 / 231 = 0
    16'b01001011_11101000 : OUT <= 0;  //75 / 232 = 0
    16'b01001011_11101001 : OUT <= 0;  //75 / 233 = 0
    16'b01001011_11101010 : OUT <= 0;  //75 / 234 = 0
    16'b01001011_11101011 : OUT <= 0;  //75 / 235 = 0
    16'b01001011_11101100 : OUT <= 0;  //75 / 236 = 0
    16'b01001011_11101101 : OUT <= 0;  //75 / 237 = 0
    16'b01001011_11101110 : OUT <= 0;  //75 / 238 = 0
    16'b01001011_11101111 : OUT <= 0;  //75 / 239 = 0
    16'b01001011_11110000 : OUT <= 0;  //75 / 240 = 0
    16'b01001011_11110001 : OUT <= 0;  //75 / 241 = 0
    16'b01001011_11110010 : OUT <= 0;  //75 / 242 = 0
    16'b01001011_11110011 : OUT <= 0;  //75 / 243 = 0
    16'b01001011_11110100 : OUT <= 0;  //75 / 244 = 0
    16'b01001011_11110101 : OUT <= 0;  //75 / 245 = 0
    16'b01001011_11110110 : OUT <= 0;  //75 / 246 = 0
    16'b01001011_11110111 : OUT <= 0;  //75 / 247 = 0
    16'b01001011_11111000 : OUT <= 0;  //75 / 248 = 0
    16'b01001011_11111001 : OUT <= 0;  //75 / 249 = 0
    16'b01001011_11111010 : OUT <= 0;  //75 / 250 = 0
    16'b01001011_11111011 : OUT <= 0;  //75 / 251 = 0
    16'b01001011_11111100 : OUT <= 0;  //75 / 252 = 0
    16'b01001011_11111101 : OUT <= 0;  //75 / 253 = 0
    16'b01001011_11111110 : OUT <= 0;  //75 / 254 = 0
    16'b01001011_11111111 : OUT <= 0;  //75 / 255 = 0
    16'b01001100_00000000 : OUT <= 0;  //76 / 0 = 0
    16'b01001100_00000001 : OUT <= 76;  //76 / 1 = 76
    16'b01001100_00000010 : OUT <= 38;  //76 / 2 = 38
    16'b01001100_00000011 : OUT <= 25;  //76 / 3 = 25
    16'b01001100_00000100 : OUT <= 19;  //76 / 4 = 19
    16'b01001100_00000101 : OUT <= 15;  //76 / 5 = 15
    16'b01001100_00000110 : OUT <= 12;  //76 / 6 = 12
    16'b01001100_00000111 : OUT <= 10;  //76 / 7 = 10
    16'b01001100_00001000 : OUT <= 9;  //76 / 8 = 9
    16'b01001100_00001001 : OUT <= 8;  //76 / 9 = 8
    16'b01001100_00001010 : OUT <= 7;  //76 / 10 = 7
    16'b01001100_00001011 : OUT <= 6;  //76 / 11 = 6
    16'b01001100_00001100 : OUT <= 6;  //76 / 12 = 6
    16'b01001100_00001101 : OUT <= 5;  //76 / 13 = 5
    16'b01001100_00001110 : OUT <= 5;  //76 / 14 = 5
    16'b01001100_00001111 : OUT <= 5;  //76 / 15 = 5
    16'b01001100_00010000 : OUT <= 4;  //76 / 16 = 4
    16'b01001100_00010001 : OUT <= 4;  //76 / 17 = 4
    16'b01001100_00010010 : OUT <= 4;  //76 / 18 = 4
    16'b01001100_00010011 : OUT <= 4;  //76 / 19 = 4
    16'b01001100_00010100 : OUT <= 3;  //76 / 20 = 3
    16'b01001100_00010101 : OUT <= 3;  //76 / 21 = 3
    16'b01001100_00010110 : OUT <= 3;  //76 / 22 = 3
    16'b01001100_00010111 : OUT <= 3;  //76 / 23 = 3
    16'b01001100_00011000 : OUT <= 3;  //76 / 24 = 3
    16'b01001100_00011001 : OUT <= 3;  //76 / 25 = 3
    16'b01001100_00011010 : OUT <= 2;  //76 / 26 = 2
    16'b01001100_00011011 : OUT <= 2;  //76 / 27 = 2
    16'b01001100_00011100 : OUT <= 2;  //76 / 28 = 2
    16'b01001100_00011101 : OUT <= 2;  //76 / 29 = 2
    16'b01001100_00011110 : OUT <= 2;  //76 / 30 = 2
    16'b01001100_00011111 : OUT <= 2;  //76 / 31 = 2
    16'b01001100_00100000 : OUT <= 2;  //76 / 32 = 2
    16'b01001100_00100001 : OUT <= 2;  //76 / 33 = 2
    16'b01001100_00100010 : OUT <= 2;  //76 / 34 = 2
    16'b01001100_00100011 : OUT <= 2;  //76 / 35 = 2
    16'b01001100_00100100 : OUT <= 2;  //76 / 36 = 2
    16'b01001100_00100101 : OUT <= 2;  //76 / 37 = 2
    16'b01001100_00100110 : OUT <= 2;  //76 / 38 = 2
    16'b01001100_00100111 : OUT <= 1;  //76 / 39 = 1
    16'b01001100_00101000 : OUT <= 1;  //76 / 40 = 1
    16'b01001100_00101001 : OUT <= 1;  //76 / 41 = 1
    16'b01001100_00101010 : OUT <= 1;  //76 / 42 = 1
    16'b01001100_00101011 : OUT <= 1;  //76 / 43 = 1
    16'b01001100_00101100 : OUT <= 1;  //76 / 44 = 1
    16'b01001100_00101101 : OUT <= 1;  //76 / 45 = 1
    16'b01001100_00101110 : OUT <= 1;  //76 / 46 = 1
    16'b01001100_00101111 : OUT <= 1;  //76 / 47 = 1
    16'b01001100_00110000 : OUT <= 1;  //76 / 48 = 1
    16'b01001100_00110001 : OUT <= 1;  //76 / 49 = 1
    16'b01001100_00110010 : OUT <= 1;  //76 / 50 = 1
    16'b01001100_00110011 : OUT <= 1;  //76 / 51 = 1
    16'b01001100_00110100 : OUT <= 1;  //76 / 52 = 1
    16'b01001100_00110101 : OUT <= 1;  //76 / 53 = 1
    16'b01001100_00110110 : OUT <= 1;  //76 / 54 = 1
    16'b01001100_00110111 : OUT <= 1;  //76 / 55 = 1
    16'b01001100_00111000 : OUT <= 1;  //76 / 56 = 1
    16'b01001100_00111001 : OUT <= 1;  //76 / 57 = 1
    16'b01001100_00111010 : OUT <= 1;  //76 / 58 = 1
    16'b01001100_00111011 : OUT <= 1;  //76 / 59 = 1
    16'b01001100_00111100 : OUT <= 1;  //76 / 60 = 1
    16'b01001100_00111101 : OUT <= 1;  //76 / 61 = 1
    16'b01001100_00111110 : OUT <= 1;  //76 / 62 = 1
    16'b01001100_00111111 : OUT <= 1;  //76 / 63 = 1
    16'b01001100_01000000 : OUT <= 1;  //76 / 64 = 1
    16'b01001100_01000001 : OUT <= 1;  //76 / 65 = 1
    16'b01001100_01000010 : OUT <= 1;  //76 / 66 = 1
    16'b01001100_01000011 : OUT <= 1;  //76 / 67 = 1
    16'b01001100_01000100 : OUT <= 1;  //76 / 68 = 1
    16'b01001100_01000101 : OUT <= 1;  //76 / 69 = 1
    16'b01001100_01000110 : OUT <= 1;  //76 / 70 = 1
    16'b01001100_01000111 : OUT <= 1;  //76 / 71 = 1
    16'b01001100_01001000 : OUT <= 1;  //76 / 72 = 1
    16'b01001100_01001001 : OUT <= 1;  //76 / 73 = 1
    16'b01001100_01001010 : OUT <= 1;  //76 / 74 = 1
    16'b01001100_01001011 : OUT <= 1;  //76 / 75 = 1
    16'b01001100_01001100 : OUT <= 1;  //76 / 76 = 1
    16'b01001100_01001101 : OUT <= 0;  //76 / 77 = 0
    16'b01001100_01001110 : OUT <= 0;  //76 / 78 = 0
    16'b01001100_01001111 : OUT <= 0;  //76 / 79 = 0
    16'b01001100_01010000 : OUT <= 0;  //76 / 80 = 0
    16'b01001100_01010001 : OUT <= 0;  //76 / 81 = 0
    16'b01001100_01010010 : OUT <= 0;  //76 / 82 = 0
    16'b01001100_01010011 : OUT <= 0;  //76 / 83 = 0
    16'b01001100_01010100 : OUT <= 0;  //76 / 84 = 0
    16'b01001100_01010101 : OUT <= 0;  //76 / 85 = 0
    16'b01001100_01010110 : OUT <= 0;  //76 / 86 = 0
    16'b01001100_01010111 : OUT <= 0;  //76 / 87 = 0
    16'b01001100_01011000 : OUT <= 0;  //76 / 88 = 0
    16'b01001100_01011001 : OUT <= 0;  //76 / 89 = 0
    16'b01001100_01011010 : OUT <= 0;  //76 / 90 = 0
    16'b01001100_01011011 : OUT <= 0;  //76 / 91 = 0
    16'b01001100_01011100 : OUT <= 0;  //76 / 92 = 0
    16'b01001100_01011101 : OUT <= 0;  //76 / 93 = 0
    16'b01001100_01011110 : OUT <= 0;  //76 / 94 = 0
    16'b01001100_01011111 : OUT <= 0;  //76 / 95 = 0
    16'b01001100_01100000 : OUT <= 0;  //76 / 96 = 0
    16'b01001100_01100001 : OUT <= 0;  //76 / 97 = 0
    16'b01001100_01100010 : OUT <= 0;  //76 / 98 = 0
    16'b01001100_01100011 : OUT <= 0;  //76 / 99 = 0
    16'b01001100_01100100 : OUT <= 0;  //76 / 100 = 0
    16'b01001100_01100101 : OUT <= 0;  //76 / 101 = 0
    16'b01001100_01100110 : OUT <= 0;  //76 / 102 = 0
    16'b01001100_01100111 : OUT <= 0;  //76 / 103 = 0
    16'b01001100_01101000 : OUT <= 0;  //76 / 104 = 0
    16'b01001100_01101001 : OUT <= 0;  //76 / 105 = 0
    16'b01001100_01101010 : OUT <= 0;  //76 / 106 = 0
    16'b01001100_01101011 : OUT <= 0;  //76 / 107 = 0
    16'b01001100_01101100 : OUT <= 0;  //76 / 108 = 0
    16'b01001100_01101101 : OUT <= 0;  //76 / 109 = 0
    16'b01001100_01101110 : OUT <= 0;  //76 / 110 = 0
    16'b01001100_01101111 : OUT <= 0;  //76 / 111 = 0
    16'b01001100_01110000 : OUT <= 0;  //76 / 112 = 0
    16'b01001100_01110001 : OUT <= 0;  //76 / 113 = 0
    16'b01001100_01110010 : OUT <= 0;  //76 / 114 = 0
    16'b01001100_01110011 : OUT <= 0;  //76 / 115 = 0
    16'b01001100_01110100 : OUT <= 0;  //76 / 116 = 0
    16'b01001100_01110101 : OUT <= 0;  //76 / 117 = 0
    16'b01001100_01110110 : OUT <= 0;  //76 / 118 = 0
    16'b01001100_01110111 : OUT <= 0;  //76 / 119 = 0
    16'b01001100_01111000 : OUT <= 0;  //76 / 120 = 0
    16'b01001100_01111001 : OUT <= 0;  //76 / 121 = 0
    16'b01001100_01111010 : OUT <= 0;  //76 / 122 = 0
    16'b01001100_01111011 : OUT <= 0;  //76 / 123 = 0
    16'b01001100_01111100 : OUT <= 0;  //76 / 124 = 0
    16'b01001100_01111101 : OUT <= 0;  //76 / 125 = 0
    16'b01001100_01111110 : OUT <= 0;  //76 / 126 = 0
    16'b01001100_01111111 : OUT <= 0;  //76 / 127 = 0
    16'b01001100_10000000 : OUT <= 0;  //76 / 128 = 0
    16'b01001100_10000001 : OUT <= 0;  //76 / 129 = 0
    16'b01001100_10000010 : OUT <= 0;  //76 / 130 = 0
    16'b01001100_10000011 : OUT <= 0;  //76 / 131 = 0
    16'b01001100_10000100 : OUT <= 0;  //76 / 132 = 0
    16'b01001100_10000101 : OUT <= 0;  //76 / 133 = 0
    16'b01001100_10000110 : OUT <= 0;  //76 / 134 = 0
    16'b01001100_10000111 : OUT <= 0;  //76 / 135 = 0
    16'b01001100_10001000 : OUT <= 0;  //76 / 136 = 0
    16'b01001100_10001001 : OUT <= 0;  //76 / 137 = 0
    16'b01001100_10001010 : OUT <= 0;  //76 / 138 = 0
    16'b01001100_10001011 : OUT <= 0;  //76 / 139 = 0
    16'b01001100_10001100 : OUT <= 0;  //76 / 140 = 0
    16'b01001100_10001101 : OUT <= 0;  //76 / 141 = 0
    16'b01001100_10001110 : OUT <= 0;  //76 / 142 = 0
    16'b01001100_10001111 : OUT <= 0;  //76 / 143 = 0
    16'b01001100_10010000 : OUT <= 0;  //76 / 144 = 0
    16'b01001100_10010001 : OUT <= 0;  //76 / 145 = 0
    16'b01001100_10010010 : OUT <= 0;  //76 / 146 = 0
    16'b01001100_10010011 : OUT <= 0;  //76 / 147 = 0
    16'b01001100_10010100 : OUT <= 0;  //76 / 148 = 0
    16'b01001100_10010101 : OUT <= 0;  //76 / 149 = 0
    16'b01001100_10010110 : OUT <= 0;  //76 / 150 = 0
    16'b01001100_10010111 : OUT <= 0;  //76 / 151 = 0
    16'b01001100_10011000 : OUT <= 0;  //76 / 152 = 0
    16'b01001100_10011001 : OUT <= 0;  //76 / 153 = 0
    16'b01001100_10011010 : OUT <= 0;  //76 / 154 = 0
    16'b01001100_10011011 : OUT <= 0;  //76 / 155 = 0
    16'b01001100_10011100 : OUT <= 0;  //76 / 156 = 0
    16'b01001100_10011101 : OUT <= 0;  //76 / 157 = 0
    16'b01001100_10011110 : OUT <= 0;  //76 / 158 = 0
    16'b01001100_10011111 : OUT <= 0;  //76 / 159 = 0
    16'b01001100_10100000 : OUT <= 0;  //76 / 160 = 0
    16'b01001100_10100001 : OUT <= 0;  //76 / 161 = 0
    16'b01001100_10100010 : OUT <= 0;  //76 / 162 = 0
    16'b01001100_10100011 : OUT <= 0;  //76 / 163 = 0
    16'b01001100_10100100 : OUT <= 0;  //76 / 164 = 0
    16'b01001100_10100101 : OUT <= 0;  //76 / 165 = 0
    16'b01001100_10100110 : OUT <= 0;  //76 / 166 = 0
    16'b01001100_10100111 : OUT <= 0;  //76 / 167 = 0
    16'b01001100_10101000 : OUT <= 0;  //76 / 168 = 0
    16'b01001100_10101001 : OUT <= 0;  //76 / 169 = 0
    16'b01001100_10101010 : OUT <= 0;  //76 / 170 = 0
    16'b01001100_10101011 : OUT <= 0;  //76 / 171 = 0
    16'b01001100_10101100 : OUT <= 0;  //76 / 172 = 0
    16'b01001100_10101101 : OUT <= 0;  //76 / 173 = 0
    16'b01001100_10101110 : OUT <= 0;  //76 / 174 = 0
    16'b01001100_10101111 : OUT <= 0;  //76 / 175 = 0
    16'b01001100_10110000 : OUT <= 0;  //76 / 176 = 0
    16'b01001100_10110001 : OUT <= 0;  //76 / 177 = 0
    16'b01001100_10110010 : OUT <= 0;  //76 / 178 = 0
    16'b01001100_10110011 : OUT <= 0;  //76 / 179 = 0
    16'b01001100_10110100 : OUT <= 0;  //76 / 180 = 0
    16'b01001100_10110101 : OUT <= 0;  //76 / 181 = 0
    16'b01001100_10110110 : OUT <= 0;  //76 / 182 = 0
    16'b01001100_10110111 : OUT <= 0;  //76 / 183 = 0
    16'b01001100_10111000 : OUT <= 0;  //76 / 184 = 0
    16'b01001100_10111001 : OUT <= 0;  //76 / 185 = 0
    16'b01001100_10111010 : OUT <= 0;  //76 / 186 = 0
    16'b01001100_10111011 : OUT <= 0;  //76 / 187 = 0
    16'b01001100_10111100 : OUT <= 0;  //76 / 188 = 0
    16'b01001100_10111101 : OUT <= 0;  //76 / 189 = 0
    16'b01001100_10111110 : OUT <= 0;  //76 / 190 = 0
    16'b01001100_10111111 : OUT <= 0;  //76 / 191 = 0
    16'b01001100_11000000 : OUT <= 0;  //76 / 192 = 0
    16'b01001100_11000001 : OUT <= 0;  //76 / 193 = 0
    16'b01001100_11000010 : OUT <= 0;  //76 / 194 = 0
    16'b01001100_11000011 : OUT <= 0;  //76 / 195 = 0
    16'b01001100_11000100 : OUT <= 0;  //76 / 196 = 0
    16'b01001100_11000101 : OUT <= 0;  //76 / 197 = 0
    16'b01001100_11000110 : OUT <= 0;  //76 / 198 = 0
    16'b01001100_11000111 : OUT <= 0;  //76 / 199 = 0
    16'b01001100_11001000 : OUT <= 0;  //76 / 200 = 0
    16'b01001100_11001001 : OUT <= 0;  //76 / 201 = 0
    16'b01001100_11001010 : OUT <= 0;  //76 / 202 = 0
    16'b01001100_11001011 : OUT <= 0;  //76 / 203 = 0
    16'b01001100_11001100 : OUT <= 0;  //76 / 204 = 0
    16'b01001100_11001101 : OUT <= 0;  //76 / 205 = 0
    16'b01001100_11001110 : OUT <= 0;  //76 / 206 = 0
    16'b01001100_11001111 : OUT <= 0;  //76 / 207 = 0
    16'b01001100_11010000 : OUT <= 0;  //76 / 208 = 0
    16'b01001100_11010001 : OUT <= 0;  //76 / 209 = 0
    16'b01001100_11010010 : OUT <= 0;  //76 / 210 = 0
    16'b01001100_11010011 : OUT <= 0;  //76 / 211 = 0
    16'b01001100_11010100 : OUT <= 0;  //76 / 212 = 0
    16'b01001100_11010101 : OUT <= 0;  //76 / 213 = 0
    16'b01001100_11010110 : OUT <= 0;  //76 / 214 = 0
    16'b01001100_11010111 : OUT <= 0;  //76 / 215 = 0
    16'b01001100_11011000 : OUT <= 0;  //76 / 216 = 0
    16'b01001100_11011001 : OUT <= 0;  //76 / 217 = 0
    16'b01001100_11011010 : OUT <= 0;  //76 / 218 = 0
    16'b01001100_11011011 : OUT <= 0;  //76 / 219 = 0
    16'b01001100_11011100 : OUT <= 0;  //76 / 220 = 0
    16'b01001100_11011101 : OUT <= 0;  //76 / 221 = 0
    16'b01001100_11011110 : OUT <= 0;  //76 / 222 = 0
    16'b01001100_11011111 : OUT <= 0;  //76 / 223 = 0
    16'b01001100_11100000 : OUT <= 0;  //76 / 224 = 0
    16'b01001100_11100001 : OUT <= 0;  //76 / 225 = 0
    16'b01001100_11100010 : OUT <= 0;  //76 / 226 = 0
    16'b01001100_11100011 : OUT <= 0;  //76 / 227 = 0
    16'b01001100_11100100 : OUT <= 0;  //76 / 228 = 0
    16'b01001100_11100101 : OUT <= 0;  //76 / 229 = 0
    16'b01001100_11100110 : OUT <= 0;  //76 / 230 = 0
    16'b01001100_11100111 : OUT <= 0;  //76 / 231 = 0
    16'b01001100_11101000 : OUT <= 0;  //76 / 232 = 0
    16'b01001100_11101001 : OUT <= 0;  //76 / 233 = 0
    16'b01001100_11101010 : OUT <= 0;  //76 / 234 = 0
    16'b01001100_11101011 : OUT <= 0;  //76 / 235 = 0
    16'b01001100_11101100 : OUT <= 0;  //76 / 236 = 0
    16'b01001100_11101101 : OUT <= 0;  //76 / 237 = 0
    16'b01001100_11101110 : OUT <= 0;  //76 / 238 = 0
    16'b01001100_11101111 : OUT <= 0;  //76 / 239 = 0
    16'b01001100_11110000 : OUT <= 0;  //76 / 240 = 0
    16'b01001100_11110001 : OUT <= 0;  //76 / 241 = 0
    16'b01001100_11110010 : OUT <= 0;  //76 / 242 = 0
    16'b01001100_11110011 : OUT <= 0;  //76 / 243 = 0
    16'b01001100_11110100 : OUT <= 0;  //76 / 244 = 0
    16'b01001100_11110101 : OUT <= 0;  //76 / 245 = 0
    16'b01001100_11110110 : OUT <= 0;  //76 / 246 = 0
    16'b01001100_11110111 : OUT <= 0;  //76 / 247 = 0
    16'b01001100_11111000 : OUT <= 0;  //76 / 248 = 0
    16'b01001100_11111001 : OUT <= 0;  //76 / 249 = 0
    16'b01001100_11111010 : OUT <= 0;  //76 / 250 = 0
    16'b01001100_11111011 : OUT <= 0;  //76 / 251 = 0
    16'b01001100_11111100 : OUT <= 0;  //76 / 252 = 0
    16'b01001100_11111101 : OUT <= 0;  //76 / 253 = 0
    16'b01001100_11111110 : OUT <= 0;  //76 / 254 = 0
    16'b01001100_11111111 : OUT <= 0;  //76 / 255 = 0
    16'b01001101_00000000 : OUT <= 0;  //77 / 0 = 0
    16'b01001101_00000001 : OUT <= 77;  //77 / 1 = 77
    16'b01001101_00000010 : OUT <= 38;  //77 / 2 = 38
    16'b01001101_00000011 : OUT <= 25;  //77 / 3 = 25
    16'b01001101_00000100 : OUT <= 19;  //77 / 4 = 19
    16'b01001101_00000101 : OUT <= 15;  //77 / 5 = 15
    16'b01001101_00000110 : OUT <= 12;  //77 / 6 = 12
    16'b01001101_00000111 : OUT <= 11;  //77 / 7 = 11
    16'b01001101_00001000 : OUT <= 9;  //77 / 8 = 9
    16'b01001101_00001001 : OUT <= 8;  //77 / 9 = 8
    16'b01001101_00001010 : OUT <= 7;  //77 / 10 = 7
    16'b01001101_00001011 : OUT <= 7;  //77 / 11 = 7
    16'b01001101_00001100 : OUT <= 6;  //77 / 12 = 6
    16'b01001101_00001101 : OUT <= 5;  //77 / 13 = 5
    16'b01001101_00001110 : OUT <= 5;  //77 / 14 = 5
    16'b01001101_00001111 : OUT <= 5;  //77 / 15 = 5
    16'b01001101_00010000 : OUT <= 4;  //77 / 16 = 4
    16'b01001101_00010001 : OUT <= 4;  //77 / 17 = 4
    16'b01001101_00010010 : OUT <= 4;  //77 / 18 = 4
    16'b01001101_00010011 : OUT <= 4;  //77 / 19 = 4
    16'b01001101_00010100 : OUT <= 3;  //77 / 20 = 3
    16'b01001101_00010101 : OUT <= 3;  //77 / 21 = 3
    16'b01001101_00010110 : OUT <= 3;  //77 / 22 = 3
    16'b01001101_00010111 : OUT <= 3;  //77 / 23 = 3
    16'b01001101_00011000 : OUT <= 3;  //77 / 24 = 3
    16'b01001101_00011001 : OUT <= 3;  //77 / 25 = 3
    16'b01001101_00011010 : OUT <= 2;  //77 / 26 = 2
    16'b01001101_00011011 : OUT <= 2;  //77 / 27 = 2
    16'b01001101_00011100 : OUT <= 2;  //77 / 28 = 2
    16'b01001101_00011101 : OUT <= 2;  //77 / 29 = 2
    16'b01001101_00011110 : OUT <= 2;  //77 / 30 = 2
    16'b01001101_00011111 : OUT <= 2;  //77 / 31 = 2
    16'b01001101_00100000 : OUT <= 2;  //77 / 32 = 2
    16'b01001101_00100001 : OUT <= 2;  //77 / 33 = 2
    16'b01001101_00100010 : OUT <= 2;  //77 / 34 = 2
    16'b01001101_00100011 : OUT <= 2;  //77 / 35 = 2
    16'b01001101_00100100 : OUT <= 2;  //77 / 36 = 2
    16'b01001101_00100101 : OUT <= 2;  //77 / 37 = 2
    16'b01001101_00100110 : OUT <= 2;  //77 / 38 = 2
    16'b01001101_00100111 : OUT <= 1;  //77 / 39 = 1
    16'b01001101_00101000 : OUT <= 1;  //77 / 40 = 1
    16'b01001101_00101001 : OUT <= 1;  //77 / 41 = 1
    16'b01001101_00101010 : OUT <= 1;  //77 / 42 = 1
    16'b01001101_00101011 : OUT <= 1;  //77 / 43 = 1
    16'b01001101_00101100 : OUT <= 1;  //77 / 44 = 1
    16'b01001101_00101101 : OUT <= 1;  //77 / 45 = 1
    16'b01001101_00101110 : OUT <= 1;  //77 / 46 = 1
    16'b01001101_00101111 : OUT <= 1;  //77 / 47 = 1
    16'b01001101_00110000 : OUT <= 1;  //77 / 48 = 1
    16'b01001101_00110001 : OUT <= 1;  //77 / 49 = 1
    16'b01001101_00110010 : OUT <= 1;  //77 / 50 = 1
    16'b01001101_00110011 : OUT <= 1;  //77 / 51 = 1
    16'b01001101_00110100 : OUT <= 1;  //77 / 52 = 1
    16'b01001101_00110101 : OUT <= 1;  //77 / 53 = 1
    16'b01001101_00110110 : OUT <= 1;  //77 / 54 = 1
    16'b01001101_00110111 : OUT <= 1;  //77 / 55 = 1
    16'b01001101_00111000 : OUT <= 1;  //77 / 56 = 1
    16'b01001101_00111001 : OUT <= 1;  //77 / 57 = 1
    16'b01001101_00111010 : OUT <= 1;  //77 / 58 = 1
    16'b01001101_00111011 : OUT <= 1;  //77 / 59 = 1
    16'b01001101_00111100 : OUT <= 1;  //77 / 60 = 1
    16'b01001101_00111101 : OUT <= 1;  //77 / 61 = 1
    16'b01001101_00111110 : OUT <= 1;  //77 / 62 = 1
    16'b01001101_00111111 : OUT <= 1;  //77 / 63 = 1
    16'b01001101_01000000 : OUT <= 1;  //77 / 64 = 1
    16'b01001101_01000001 : OUT <= 1;  //77 / 65 = 1
    16'b01001101_01000010 : OUT <= 1;  //77 / 66 = 1
    16'b01001101_01000011 : OUT <= 1;  //77 / 67 = 1
    16'b01001101_01000100 : OUT <= 1;  //77 / 68 = 1
    16'b01001101_01000101 : OUT <= 1;  //77 / 69 = 1
    16'b01001101_01000110 : OUT <= 1;  //77 / 70 = 1
    16'b01001101_01000111 : OUT <= 1;  //77 / 71 = 1
    16'b01001101_01001000 : OUT <= 1;  //77 / 72 = 1
    16'b01001101_01001001 : OUT <= 1;  //77 / 73 = 1
    16'b01001101_01001010 : OUT <= 1;  //77 / 74 = 1
    16'b01001101_01001011 : OUT <= 1;  //77 / 75 = 1
    16'b01001101_01001100 : OUT <= 1;  //77 / 76 = 1
    16'b01001101_01001101 : OUT <= 1;  //77 / 77 = 1
    16'b01001101_01001110 : OUT <= 0;  //77 / 78 = 0
    16'b01001101_01001111 : OUT <= 0;  //77 / 79 = 0
    16'b01001101_01010000 : OUT <= 0;  //77 / 80 = 0
    16'b01001101_01010001 : OUT <= 0;  //77 / 81 = 0
    16'b01001101_01010010 : OUT <= 0;  //77 / 82 = 0
    16'b01001101_01010011 : OUT <= 0;  //77 / 83 = 0
    16'b01001101_01010100 : OUT <= 0;  //77 / 84 = 0
    16'b01001101_01010101 : OUT <= 0;  //77 / 85 = 0
    16'b01001101_01010110 : OUT <= 0;  //77 / 86 = 0
    16'b01001101_01010111 : OUT <= 0;  //77 / 87 = 0
    16'b01001101_01011000 : OUT <= 0;  //77 / 88 = 0
    16'b01001101_01011001 : OUT <= 0;  //77 / 89 = 0
    16'b01001101_01011010 : OUT <= 0;  //77 / 90 = 0
    16'b01001101_01011011 : OUT <= 0;  //77 / 91 = 0
    16'b01001101_01011100 : OUT <= 0;  //77 / 92 = 0
    16'b01001101_01011101 : OUT <= 0;  //77 / 93 = 0
    16'b01001101_01011110 : OUT <= 0;  //77 / 94 = 0
    16'b01001101_01011111 : OUT <= 0;  //77 / 95 = 0
    16'b01001101_01100000 : OUT <= 0;  //77 / 96 = 0
    16'b01001101_01100001 : OUT <= 0;  //77 / 97 = 0
    16'b01001101_01100010 : OUT <= 0;  //77 / 98 = 0
    16'b01001101_01100011 : OUT <= 0;  //77 / 99 = 0
    16'b01001101_01100100 : OUT <= 0;  //77 / 100 = 0
    16'b01001101_01100101 : OUT <= 0;  //77 / 101 = 0
    16'b01001101_01100110 : OUT <= 0;  //77 / 102 = 0
    16'b01001101_01100111 : OUT <= 0;  //77 / 103 = 0
    16'b01001101_01101000 : OUT <= 0;  //77 / 104 = 0
    16'b01001101_01101001 : OUT <= 0;  //77 / 105 = 0
    16'b01001101_01101010 : OUT <= 0;  //77 / 106 = 0
    16'b01001101_01101011 : OUT <= 0;  //77 / 107 = 0
    16'b01001101_01101100 : OUT <= 0;  //77 / 108 = 0
    16'b01001101_01101101 : OUT <= 0;  //77 / 109 = 0
    16'b01001101_01101110 : OUT <= 0;  //77 / 110 = 0
    16'b01001101_01101111 : OUT <= 0;  //77 / 111 = 0
    16'b01001101_01110000 : OUT <= 0;  //77 / 112 = 0
    16'b01001101_01110001 : OUT <= 0;  //77 / 113 = 0
    16'b01001101_01110010 : OUT <= 0;  //77 / 114 = 0
    16'b01001101_01110011 : OUT <= 0;  //77 / 115 = 0
    16'b01001101_01110100 : OUT <= 0;  //77 / 116 = 0
    16'b01001101_01110101 : OUT <= 0;  //77 / 117 = 0
    16'b01001101_01110110 : OUT <= 0;  //77 / 118 = 0
    16'b01001101_01110111 : OUT <= 0;  //77 / 119 = 0
    16'b01001101_01111000 : OUT <= 0;  //77 / 120 = 0
    16'b01001101_01111001 : OUT <= 0;  //77 / 121 = 0
    16'b01001101_01111010 : OUT <= 0;  //77 / 122 = 0
    16'b01001101_01111011 : OUT <= 0;  //77 / 123 = 0
    16'b01001101_01111100 : OUT <= 0;  //77 / 124 = 0
    16'b01001101_01111101 : OUT <= 0;  //77 / 125 = 0
    16'b01001101_01111110 : OUT <= 0;  //77 / 126 = 0
    16'b01001101_01111111 : OUT <= 0;  //77 / 127 = 0
    16'b01001101_10000000 : OUT <= 0;  //77 / 128 = 0
    16'b01001101_10000001 : OUT <= 0;  //77 / 129 = 0
    16'b01001101_10000010 : OUT <= 0;  //77 / 130 = 0
    16'b01001101_10000011 : OUT <= 0;  //77 / 131 = 0
    16'b01001101_10000100 : OUT <= 0;  //77 / 132 = 0
    16'b01001101_10000101 : OUT <= 0;  //77 / 133 = 0
    16'b01001101_10000110 : OUT <= 0;  //77 / 134 = 0
    16'b01001101_10000111 : OUT <= 0;  //77 / 135 = 0
    16'b01001101_10001000 : OUT <= 0;  //77 / 136 = 0
    16'b01001101_10001001 : OUT <= 0;  //77 / 137 = 0
    16'b01001101_10001010 : OUT <= 0;  //77 / 138 = 0
    16'b01001101_10001011 : OUT <= 0;  //77 / 139 = 0
    16'b01001101_10001100 : OUT <= 0;  //77 / 140 = 0
    16'b01001101_10001101 : OUT <= 0;  //77 / 141 = 0
    16'b01001101_10001110 : OUT <= 0;  //77 / 142 = 0
    16'b01001101_10001111 : OUT <= 0;  //77 / 143 = 0
    16'b01001101_10010000 : OUT <= 0;  //77 / 144 = 0
    16'b01001101_10010001 : OUT <= 0;  //77 / 145 = 0
    16'b01001101_10010010 : OUT <= 0;  //77 / 146 = 0
    16'b01001101_10010011 : OUT <= 0;  //77 / 147 = 0
    16'b01001101_10010100 : OUT <= 0;  //77 / 148 = 0
    16'b01001101_10010101 : OUT <= 0;  //77 / 149 = 0
    16'b01001101_10010110 : OUT <= 0;  //77 / 150 = 0
    16'b01001101_10010111 : OUT <= 0;  //77 / 151 = 0
    16'b01001101_10011000 : OUT <= 0;  //77 / 152 = 0
    16'b01001101_10011001 : OUT <= 0;  //77 / 153 = 0
    16'b01001101_10011010 : OUT <= 0;  //77 / 154 = 0
    16'b01001101_10011011 : OUT <= 0;  //77 / 155 = 0
    16'b01001101_10011100 : OUT <= 0;  //77 / 156 = 0
    16'b01001101_10011101 : OUT <= 0;  //77 / 157 = 0
    16'b01001101_10011110 : OUT <= 0;  //77 / 158 = 0
    16'b01001101_10011111 : OUT <= 0;  //77 / 159 = 0
    16'b01001101_10100000 : OUT <= 0;  //77 / 160 = 0
    16'b01001101_10100001 : OUT <= 0;  //77 / 161 = 0
    16'b01001101_10100010 : OUT <= 0;  //77 / 162 = 0
    16'b01001101_10100011 : OUT <= 0;  //77 / 163 = 0
    16'b01001101_10100100 : OUT <= 0;  //77 / 164 = 0
    16'b01001101_10100101 : OUT <= 0;  //77 / 165 = 0
    16'b01001101_10100110 : OUT <= 0;  //77 / 166 = 0
    16'b01001101_10100111 : OUT <= 0;  //77 / 167 = 0
    16'b01001101_10101000 : OUT <= 0;  //77 / 168 = 0
    16'b01001101_10101001 : OUT <= 0;  //77 / 169 = 0
    16'b01001101_10101010 : OUT <= 0;  //77 / 170 = 0
    16'b01001101_10101011 : OUT <= 0;  //77 / 171 = 0
    16'b01001101_10101100 : OUT <= 0;  //77 / 172 = 0
    16'b01001101_10101101 : OUT <= 0;  //77 / 173 = 0
    16'b01001101_10101110 : OUT <= 0;  //77 / 174 = 0
    16'b01001101_10101111 : OUT <= 0;  //77 / 175 = 0
    16'b01001101_10110000 : OUT <= 0;  //77 / 176 = 0
    16'b01001101_10110001 : OUT <= 0;  //77 / 177 = 0
    16'b01001101_10110010 : OUT <= 0;  //77 / 178 = 0
    16'b01001101_10110011 : OUT <= 0;  //77 / 179 = 0
    16'b01001101_10110100 : OUT <= 0;  //77 / 180 = 0
    16'b01001101_10110101 : OUT <= 0;  //77 / 181 = 0
    16'b01001101_10110110 : OUT <= 0;  //77 / 182 = 0
    16'b01001101_10110111 : OUT <= 0;  //77 / 183 = 0
    16'b01001101_10111000 : OUT <= 0;  //77 / 184 = 0
    16'b01001101_10111001 : OUT <= 0;  //77 / 185 = 0
    16'b01001101_10111010 : OUT <= 0;  //77 / 186 = 0
    16'b01001101_10111011 : OUT <= 0;  //77 / 187 = 0
    16'b01001101_10111100 : OUT <= 0;  //77 / 188 = 0
    16'b01001101_10111101 : OUT <= 0;  //77 / 189 = 0
    16'b01001101_10111110 : OUT <= 0;  //77 / 190 = 0
    16'b01001101_10111111 : OUT <= 0;  //77 / 191 = 0
    16'b01001101_11000000 : OUT <= 0;  //77 / 192 = 0
    16'b01001101_11000001 : OUT <= 0;  //77 / 193 = 0
    16'b01001101_11000010 : OUT <= 0;  //77 / 194 = 0
    16'b01001101_11000011 : OUT <= 0;  //77 / 195 = 0
    16'b01001101_11000100 : OUT <= 0;  //77 / 196 = 0
    16'b01001101_11000101 : OUT <= 0;  //77 / 197 = 0
    16'b01001101_11000110 : OUT <= 0;  //77 / 198 = 0
    16'b01001101_11000111 : OUT <= 0;  //77 / 199 = 0
    16'b01001101_11001000 : OUT <= 0;  //77 / 200 = 0
    16'b01001101_11001001 : OUT <= 0;  //77 / 201 = 0
    16'b01001101_11001010 : OUT <= 0;  //77 / 202 = 0
    16'b01001101_11001011 : OUT <= 0;  //77 / 203 = 0
    16'b01001101_11001100 : OUT <= 0;  //77 / 204 = 0
    16'b01001101_11001101 : OUT <= 0;  //77 / 205 = 0
    16'b01001101_11001110 : OUT <= 0;  //77 / 206 = 0
    16'b01001101_11001111 : OUT <= 0;  //77 / 207 = 0
    16'b01001101_11010000 : OUT <= 0;  //77 / 208 = 0
    16'b01001101_11010001 : OUT <= 0;  //77 / 209 = 0
    16'b01001101_11010010 : OUT <= 0;  //77 / 210 = 0
    16'b01001101_11010011 : OUT <= 0;  //77 / 211 = 0
    16'b01001101_11010100 : OUT <= 0;  //77 / 212 = 0
    16'b01001101_11010101 : OUT <= 0;  //77 / 213 = 0
    16'b01001101_11010110 : OUT <= 0;  //77 / 214 = 0
    16'b01001101_11010111 : OUT <= 0;  //77 / 215 = 0
    16'b01001101_11011000 : OUT <= 0;  //77 / 216 = 0
    16'b01001101_11011001 : OUT <= 0;  //77 / 217 = 0
    16'b01001101_11011010 : OUT <= 0;  //77 / 218 = 0
    16'b01001101_11011011 : OUT <= 0;  //77 / 219 = 0
    16'b01001101_11011100 : OUT <= 0;  //77 / 220 = 0
    16'b01001101_11011101 : OUT <= 0;  //77 / 221 = 0
    16'b01001101_11011110 : OUT <= 0;  //77 / 222 = 0
    16'b01001101_11011111 : OUT <= 0;  //77 / 223 = 0
    16'b01001101_11100000 : OUT <= 0;  //77 / 224 = 0
    16'b01001101_11100001 : OUT <= 0;  //77 / 225 = 0
    16'b01001101_11100010 : OUT <= 0;  //77 / 226 = 0
    16'b01001101_11100011 : OUT <= 0;  //77 / 227 = 0
    16'b01001101_11100100 : OUT <= 0;  //77 / 228 = 0
    16'b01001101_11100101 : OUT <= 0;  //77 / 229 = 0
    16'b01001101_11100110 : OUT <= 0;  //77 / 230 = 0
    16'b01001101_11100111 : OUT <= 0;  //77 / 231 = 0
    16'b01001101_11101000 : OUT <= 0;  //77 / 232 = 0
    16'b01001101_11101001 : OUT <= 0;  //77 / 233 = 0
    16'b01001101_11101010 : OUT <= 0;  //77 / 234 = 0
    16'b01001101_11101011 : OUT <= 0;  //77 / 235 = 0
    16'b01001101_11101100 : OUT <= 0;  //77 / 236 = 0
    16'b01001101_11101101 : OUT <= 0;  //77 / 237 = 0
    16'b01001101_11101110 : OUT <= 0;  //77 / 238 = 0
    16'b01001101_11101111 : OUT <= 0;  //77 / 239 = 0
    16'b01001101_11110000 : OUT <= 0;  //77 / 240 = 0
    16'b01001101_11110001 : OUT <= 0;  //77 / 241 = 0
    16'b01001101_11110010 : OUT <= 0;  //77 / 242 = 0
    16'b01001101_11110011 : OUT <= 0;  //77 / 243 = 0
    16'b01001101_11110100 : OUT <= 0;  //77 / 244 = 0
    16'b01001101_11110101 : OUT <= 0;  //77 / 245 = 0
    16'b01001101_11110110 : OUT <= 0;  //77 / 246 = 0
    16'b01001101_11110111 : OUT <= 0;  //77 / 247 = 0
    16'b01001101_11111000 : OUT <= 0;  //77 / 248 = 0
    16'b01001101_11111001 : OUT <= 0;  //77 / 249 = 0
    16'b01001101_11111010 : OUT <= 0;  //77 / 250 = 0
    16'b01001101_11111011 : OUT <= 0;  //77 / 251 = 0
    16'b01001101_11111100 : OUT <= 0;  //77 / 252 = 0
    16'b01001101_11111101 : OUT <= 0;  //77 / 253 = 0
    16'b01001101_11111110 : OUT <= 0;  //77 / 254 = 0
    16'b01001101_11111111 : OUT <= 0;  //77 / 255 = 0
    16'b01001110_00000000 : OUT <= 0;  //78 / 0 = 0
    16'b01001110_00000001 : OUT <= 78;  //78 / 1 = 78
    16'b01001110_00000010 : OUT <= 39;  //78 / 2 = 39
    16'b01001110_00000011 : OUT <= 26;  //78 / 3 = 26
    16'b01001110_00000100 : OUT <= 19;  //78 / 4 = 19
    16'b01001110_00000101 : OUT <= 15;  //78 / 5 = 15
    16'b01001110_00000110 : OUT <= 13;  //78 / 6 = 13
    16'b01001110_00000111 : OUT <= 11;  //78 / 7 = 11
    16'b01001110_00001000 : OUT <= 9;  //78 / 8 = 9
    16'b01001110_00001001 : OUT <= 8;  //78 / 9 = 8
    16'b01001110_00001010 : OUT <= 7;  //78 / 10 = 7
    16'b01001110_00001011 : OUT <= 7;  //78 / 11 = 7
    16'b01001110_00001100 : OUT <= 6;  //78 / 12 = 6
    16'b01001110_00001101 : OUT <= 6;  //78 / 13 = 6
    16'b01001110_00001110 : OUT <= 5;  //78 / 14 = 5
    16'b01001110_00001111 : OUT <= 5;  //78 / 15 = 5
    16'b01001110_00010000 : OUT <= 4;  //78 / 16 = 4
    16'b01001110_00010001 : OUT <= 4;  //78 / 17 = 4
    16'b01001110_00010010 : OUT <= 4;  //78 / 18 = 4
    16'b01001110_00010011 : OUT <= 4;  //78 / 19 = 4
    16'b01001110_00010100 : OUT <= 3;  //78 / 20 = 3
    16'b01001110_00010101 : OUT <= 3;  //78 / 21 = 3
    16'b01001110_00010110 : OUT <= 3;  //78 / 22 = 3
    16'b01001110_00010111 : OUT <= 3;  //78 / 23 = 3
    16'b01001110_00011000 : OUT <= 3;  //78 / 24 = 3
    16'b01001110_00011001 : OUT <= 3;  //78 / 25 = 3
    16'b01001110_00011010 : OUT <= 3;  //78 / 26 = 3
    16'b01001110_00011011 : OUT <= 2;  //78 / 27 = 2
    16'b01001110_00011100 : OUT <= 2;  //78 / 28 = 2
    16'b01001110_00011101 : OUT <= 2;  //78 / 29 = 2
    16'b01001110_00011110 : OUT <= 2;  //78 / 30 = 2
    16'b01001110_00011111 : OUT <= 2;  //78 / 31 = 2
    16'b01001110_00100000 : OUT <= 2;  //78 / 32 = 2
    16'b01001110_00100001 : OUT <= 2;  //78 / 33 = 2
    16'b01001110_00100010 : OUT <= 2;  //78 / 34 = 2
    16'b01001110_00100011 : OUT <= 2;  //78 / 35 = 2
    16'b01001110_00100100 : OUT <= 2;  //78 / 36 = 2
    16'b01001110_00100101 : OUT <= 2;  //78 / 37 = 2
    16'b01001110_00100110 : OUT <= 2;  //78 / 38 = 2
    16'b01001110_00100111 : OUT <= 2;  //78 / 39 = 2
    16'b01001110_00101000 : OUT <= 1;  //78 / 40 = 1
    16'b01001110_00101001 : OUT <= 1;  //78 / 41 = 1
    16'b01001110_00101010 : OUT <= 1;  //78 / 42 = 1
    16'b01001110_00101011 : OUT <= 1;  //78 / 43 = 1
    16'b01001110_00101100 : OUT <= 1;  //78 / 44 = 1
    16'b01001110_00101101 : OUT <= 1;  //78 / 45 = 1
    16'b01001110_00101110 : OUT <= 1;  //78 / 46 = 1
    16'b01001110_00101111 : OUT <= 1;  //78 / 47 = 1
    16'b01001110_00110000 : OUT <= 1;  //78 / 48 = 1
    16'b01001110_00110001 : OUT <= 1;  //78 / 49 = 1
    16'b01001110_00110010 : OUT <= 1;  //78 / 50 = 1
    16'b01001110_00110011 : OUT <= 1;  //78 / 51 = 1
    16'b01001110_00110100 : OUT <= 1;  //78 / 52 = 1
    16'b01001110_00110101 : OUT <= 1;  //78 / 53 = 1
    16'b01001110_00110110 : OUT <= 1;  //78 / 54 = 1
    16'b01001110_00110111 : OUT <= 1;  //78 / 55 = 1
    16'b01001110_00111000 : OUT <= 1;  //78 / 56 = 1
    16'b01001110_00111001 : OUT <= 1;  //78 / 57 = 1
    16'b01001110_00111010 : OUT <= 1;  //78 / 58 = 1
    16'b01001110_00111011 : OUT <= 1;  //78 / 59 = 1
    16'b01001110_00111100 : OUT <= 1;  //78 / 60 = 1
    16'b01001110_00111101 : OUT <= 1;  //78 / 61 = 1
    16'b01001110_00111110 : OUT <= 1;  //78 / 62 = 1
    16'b01001110_00111111 : OUT <= 1;  //78 / 63 = 1
    16'b01001110_01000000 : OUT <= 1;  //78 / 64 = 1
    16'b01001110_01000001 : OUT <= 1;  //78 / 65 = 1
    16'b01001110_01000010 : OUT <= 1;  //78 / 66 = 1
    16'b01001110_01000011 : OUT <= 1;  //78 / 67 = 1
    16'b01001110_01000100 : OUT <= 1;  //78 / 68 = 1
    16'b01001110_01000101 : OUT <= 1;  //78 / 69 = 1
    16'b01001110_01000110 : OUT <= 1;  //78 / 70 = 1
    16'b01001110_01000111 : OUT <= 1;  //78 / 71 = 1
    16'b01001110_01001000 : OUT <= 1;  //78 / 72 = 1
    16'b01001110_01001001 : OUT <= 1;  //78 / 73 = 1
    16'b01001110_01001010 : OUT <= 1;  //78 / 74 = 1
    16'b01001110_01001011 : OUT <= 1;  //78 / 75 = 1
    16'b01001110_01001100 : OUT <= 1;  //78 / 76 = 1
    16'b01001110_01001101 : OUT <= 1;  //78 / 77 = 1
    16'b01001110_01001110 : OUT <= 1;  //78 / 78 = 1
    16'b01001110_01001111 : OUT <= 0;  //78 / 79 = 0
    16'b01001110_01010000 : OUT <= 0;  //78 / 80 = 0
    16'b01001110_01010001 : OUT <= 0;  //78 / 81 = 0
    16'b01001110_01010010 : OUT <= 0;  //78 / 82 = 0
    16'b01001110_01010011 : OUT <= 0;  //78 / 83 = 0
    16'b01001110_01010100 : OUT <= 0;  //78 / 84 = 0
    16'b01001110_01010101 : OUT <= 0;  //78 / 85 = 0
    16'b01001110_01010110 : OUT <= 0;  //78 / 86 = 0
    16'b01001110_01010111 : OUT <= 0;  //78 / 87 = 0
    16'b01001110_01011000 : OUT <= 0;  //78 / 88 = 0
    16'b01001110_01011001 : OUT <= 0;  //78 / 89 = 0
    16'b01001110_01011010 : OUT <= 0;  //78 / 90 = 0
    16'b01001110_01011011 : OUT <= 0;  //78 / 91 = 0
    16'b01001110_01011100 : OUT <= 0;  //78 / 92 = 0
    16'b01001110_01011101 : OUT <= 0;  //78 / 93 = 0
    16'b01001110_01011110 : OUT <= 0;  //78 / 94 = 0
    16'b01001110_01011111 : OUT <= 0;  //78 / 95 = 0
    16'b01001110_01100000 : OUT <= 0;  //78 / 96 = 0
    16'b01001110_01100001 : OUT <= 0;  //78 / 97 = 0
    16'b01001110_01100010 : OUT <= 0;  //78 / 98 = 0
    16'b01001110_01100011 : OUT <= 0;  //78 / 99 = 0
    16'b01001110_01100100 : OUT <= 0;  //78 / 100 = 0
    16'b01001110_01100101 : OUT <= 0;  //78 / 101 = 0
    16'b01001110_01100110 : OUT <= 0;  //78 / 102 = 0
    16'b01001110_01100111 : OUT <= 0;  //78 / 103 = 0
    16'b01001110_01101000 : OUT <= 0;  //78 / 104 = 0
    16'b01001110_01101001 : OUT <= 0;  //78 / 105 = 0
    16'b01001110_01101010 : OUT <= 0;  //78 / 106 = 0
    16'b01001110_01101011 : OUT <= 0;  //78 / 107 = 0
    16'b01001110_01101100 : OUT <= 0;  //78 / 108 = 0
    16'b01001110_01101101 : OUT <= 0;  //78 / 109 = 0
    16'b01001110_01101110 : OUT <= 0;  //78 / 110 = 0
    16'b01001110_01101111 : OUT <= 0;  //78 / 111 = 0
    16'b01001110_01110000 : OUT <= 0;  //78 / 112 = 0
    16'b01001110_01110001 : OUT <= 0;  //78 / 113 = 0
    16'b01001110_01110010 : OUT <= 0;  //78 / 114 = 0
    16'b01001110_01110011 : OUT <= 0;  //78 / 115 = 0
    16'b01001110_01110100 : OUT <= 0;  //78 / 116 = 0
    16'b01001110_01110101 : OUT <= 0;  //78 / 117 = 0
    16'b01001110_01110110 : OUT <= 0;  //78 / 118 = 0
    16'b01001110_01110111 : OUT <= 0;  //78 / 119 = 0
    16'b01001110_01111000 : OUT <= 0;  //78 / 120 = 0
    16'b01001110_01111001 : OUT <= 0;  //78 / 121 = 0
    16'b01001110_01111010 : OUT <= 0;  //78 / 122 = 0
    16'b01001110_01111011 : OUT <= 0;  //78 / 123 = 0
    16'b01001110_01111100 : OUT <= 0;  //78 / 124 = 0
    16'b01001110_01111101 : OUT <= 0;  //78 / 125 = 0
    16'b01001110_01111110 : OUT <= 0;  //78 / 126 = 0
    16'b01001110_01111111 : OUT <= 0;  //78 / 127 = 0
    16'b01001110_10000000 : OUT <= 0;  //78 / 128 = 0
    16'b01001110_10000001 : OUT <= 0;  //78 / 129 = 0
    16'b01001110_10000010 : OUT <= 0;  //78 / 130 = 0
    16'b01001110_10000011 : OUT <= 0;  //78 / 131 = 0
    16'b01001110_10000100 : OUT <= 0;  //78 / 132 = 0
    16'b01001110_10000101 : OUT <= 0;  //78 / 133 = 0
    16'b01001110_10000110 : OUT <= 0;  //78 / 134 = 0
    16'b01001110_10000111 : OUT <= 0;  //78 / 135 = 0
    16'b01001110_10001000 : OUT <= 0;  //78 / 136 = 0
    16'b01001110_10001001 : OUT <= 0;  //78 / 137 = 0
    16'b01001110_10001010 : OUT <= 0;  //78 / 138 = 0
    16'b01001110_10001011 : OUT <= 0;  //78 / 139 = 0
    16'b01001110_10001100 : OUT <= 0;  //78 / 140 = 0
    16'b01001110_10001101 : OUT <= 0;  //78 / 141 = 0
    16'b01001110_10001110 : OUT <= 0;  //78 / 142 = 0
    16'b01001110_10001111 : OUT <= 0;  //78 / 143 = 0
    16'b01001110_10010000 : OUT <= 0;  //78 / 144 = 0
    16'b01001110_10010001 : OUT <= 0;  //78 / 145 = 0
    16'b01001110_10010010 : OUT <= 0;  //78 / 146 = 0
    16'b01001110_10010011 : OUT <= 0;  //78 / 147 = 0
    16'b01001110_10010100 : OUT <= 0;  //78 / 148 = 0
    16'b01001110_10010101 : OUT <= 0;  //78 / 149 = 0
    16'b01001110_10010110 : OUT <= 0;  //78 / 150 = 0
    16'b01001110_10010111 : OUT <= 0;  //78 / 151 = 0
    16'b01001110_10011000 : OUT <= 0;  //78 / 152 = 0
    16'b01001110_10011001 : OUT <= 0;  //78 / 153 = 0
    16'b01001110_10011010 : OUT <= 0;  //78 / 154 = 0
    16'b01001110_10011011 : OUT <= 0;  //78 / 155 = 0
    16'b01001110_10011100 : OUT <= 0;  //78 / 156 = 0
    16'b01001110_10011101 : OUT <= 0;  //78 / 157 = 0
    16'b01001110_10011110 : OUT <= 0;  //78 / 158 = 0
    16'b01001110_10011111 : OUT <= 0;  //78 / 159 = 0
    16'b01001110_10100000 : OUT <= 0;  //78 / 160 = 0
    16'b01001110_10100001 : OUT <= 0;  //78 / 161 = 0
    16'b01001110_10100010 : OUT <= 0;  //78 / 162 = 0
    16'b01001110_10100011 : OUT <= 0;  //78 / 163 = 0
    16'b01001110_10100100 : OUT <= 0;  //78 / 164 = 0
    16'b01001110_10100101 : OUT <= 0;  //78 / 165 = 0
    16'b01001110_10100110 : OUT <= 0;  //78 / 166 = 0
    16'b01001110_10100111 : OUT <= 0;  //78 / 167 = 0
    16'b01001110_10101000 : OUT <= 0;  //78 / 168 = 0
    16'b01001110_10101001 : OUT <= 0;  //78 / 169 = 0
    16'b01001110_10101010 : OUT <= 0;  //78 / 170 = 0
    16'b01001110_10101011 : OUT <= 0;  //78 / 171 = 0
    16'b01001110_10101100 : OUT <= 0;  //78 / 172 = 0
    16'b01001110_10101101 : OUT <= 0;  //78 / 173 = 0
    16'b01001110_10101110 : OUT <= 0;  //78 / 174 = 0
    16'b01001110_10101111 : OUT <= 0;  //78 / 175 = 0
    16'b01001110_10110000 : OUT <= 0;  //78 / 176 = 0
    16'b01001110_10110001 : OUT <= 0;  //78 / 177 = 0
    16'b01001110_10110010 : OUT <= 0;  //78 / 178 = 0
    16'b01001110_10110011 : OUT <= 0;  //78 / 179 = 0
    16'b01001110_10110100 : OUT <= 0;  //78 / 180 = 0
    16'b01001110_10110101 : OUT <= 0;  //78 / 181 = 0
    16'b01001110_10110110 : OUT <= 0;  //78 / 182 = 0
    16'b01001110_10110111 : OUT <= 0;  //78 / 183 = 0
    16'b01001110_10111000 : OUT <= 0;  //78 / 184 = 0
    16'b01001110_10111001 : OUT <= 0;  //78 / 185 = 0
    16'b01001110_10111010 : OUT <= 0;  //78 / 186 = 0
    16'b01001110_10111011 : OUT <= 0;  //78 / 187 = 0
    16'b01001110_10111100 : OUT <= 0;  //78 / 188 = 0
    16'b01001110_10111101 : OUT <= 0;  //78 / 189 = 0
    16'b01001110_10111110 : OUT <= 0;  //78 / 190 = 0
    16'b01001110_10111111 : OUT <= 0;  //78 / 191 = 0
    16'b01001110_11000000 : OUT <= 0;  //78 / 192 = 0
    16'b01001110_11000001 : OUT <= 0;  //78 / 193 = 0
    16'b01001110_11000010 : OUT <= 0;  //78 / 194 = 0
    16'b01001110_11000011 : OUT <= 0;  //78 / 195 = 0
    16'b01001110_11000100 : OUT <= 0;  //78 / 196 = 0
    16'b01001110_11000101 : OUT <= 0;  //78 / 197 = 0
    16'b01001110_11000110 : OUT <= 0;  //78 / 198 = 0
    16'b01001110_11000111 : OUT <= 0;  //78 / 199 = 0
    16'b01001110_11001000 : OUT <= 0;  //78 / 200 = 0
    16'b01001110_11001001 : OUT <= 0;  //78 / 201 = 0
    16'b01001110_11001010 : OUT <= 0;  //78 / 202 = 0
    16'b01001110_11001011 : OUT <= 0;  //78 / 203 = 0
    16'b01001110_11001100 : OUT <= 0;  //78 / 204 = 0
    16'b01001110_11001101 : OUT <= 0;  //78 / 205 = 0
    16'b01001110_11001110 : OUT <= 0;  //78 / 206 = 0
    16'b01001110_11001111 : OUT <= 0;  //78 / 207 = 0
    16'b01001110_11010000 : OUT <= 0;  //78 / 208 = 0
    16'b01001110_11010001 : OUT <= 0;  //78 / 209 = 0
    16'b01001110_11010010 : OUT <= 0;  //78 / 210 = 0
    16'b01001110_11010011 : OUT <= 0;  //78 / 211 = 0
    16'b01001110_11010100 : OUT <= 0;  //78 / 212 = 0
    16'b01001110_11010101 : OUT <= 0;  //78 / 213 = 0
    16'b01001110_11010110 : OUT <= 0;  //78 / 214 = 0
    16'b01001110_11010111 : OUT <= 0;  //78 / 215 = 0
    16'b01001110_11011000 : OUT <= 0;  //78 / 216 = 0
    16'b01001110_11011001 : OUT <= 0;  //78 / 217 = 0
    16'b01001110_11011010 : OUT <= 0;  //78 / 218 = 0
    16'b01001110_11011011 : OUT <= 0;  //78 / 219 = 0
    16'b01001110_11011100 : OUT <= 0;  //78 / 220 = 0
    16'b01001110_11011101 : OUT <= 0;  //78 / 221 = 0
    16'b01001110_11011110 : OUT <= 0;  //78 / 222 = 0
    16'b01001110_11011111 : OUT <= 0;  //78 / 223 = 0
    16'b01001110_11100000 : OUT <= 0;  //78 / 224 = 0
    16'b01001110_11100001 : OUT <= 0;  //78 / 225 = 0
    16'b01001110_11100010 : OUT <= 0;  //78 / 226 = 0
    16'b01001110_11100011 : OUT <= 0;  //78 / 227 = 0
    16'b01001110_11100100 : OUT <= 0;  //78 / 228 = 0
    16'b01001110_11100101 : OUT <= 0;  //78 / 229 = 0
    16'b01001110_11100110 : OUT <= 0;  //78 / 230 = 0
    16'b01001110_11100111 : OUT <= 0;  //78 / 231 = 0
    16'b01001110_11101000 : OUT <= 0;  //78 / 232 = 0
    16'b01001110_11101001 : OUT <= 0;  //78 / 233 = 0
    16'b01001110_11101010 : OUT <= 0;  //78 / 234 = 0
    16'b01001110_11101011 : OUT <= 0;  //78 / 235 = 0
    16'b01001110_11101100 : OUT <= 0;  //78 / 236 = 0
    16'b01001110_11101101 : OUT <= 0;  //78 / 237 = 0
    16'b01001110_11101110 : OUT <= 0;  //78 / 238 = 0
    16'b01001110_11101111 : OUT <= 0;  //78 / 239 = 0
    16'b01001110_11110000 : OUT <= 0;  //78 / 240 = 0
    16'b01001110_11110001 : OUT <= 0;  //78 / 241 = 0
    16'b01001110_11110010 : OUT <= 0;  //78 / 242 = 0
    16'b01001110_11110011 : OUT <= 0;  //78 / 243 = 0
    16'b01001110_11110100 : OUT <= 0;  //78 / 244 = 0
    16'b01001110_11110101 : OUT <= 0;  //78 / 245 = 0
    16'b01001110_11110110 : OUT <= 0;  //78 / 246 = 0
    16'b01001110_11110111 : OUT <= 0;  //78 / 247 = 0
    16'b01001110_11111000 : OUT <= 0;  //78 / 248 = 0
    16'b01001110_11111001 : OUT <= 0;  //78 / 249 = 0
    16'b01001110_11111010 : OUT <= 0;  //78 / 250 = 0
    16'b01001110_11111011 : OUT <= 0;  //78 / 251 = 0
    16'b01001110_11111100 : OUT <= 0;  //78 / 252 = 0
    16'b01001110_11111101 : OUT <= 0;  //78 / 253 = 0
    16'b01001110_11111110 : OUT <= 0;  //78 / 254 = 0
    16'b01001110_11111111 : OUT <= 0;  //78 / 255 = 0
    16'b01001111_00000000 : OUT <= 0;  //79 / 0 = 0
    16'b01001111_00000001 : OUT <= 79;  //79 / 1 = 79
    16'b01001111_00000010 : OUT <= 39;  //79 / 2 = 39
    16'b01001111_00000011 : OUT <= 26;  //79 / 3 = 26
    16'b01001111_00000100 : OUT <= 19;  //79 / 4 = 19
    16'b01001111_00000101 : OUT <= 15;  //79 / 5 = 15
    16'b01001111_00000110 : OUT <= 13;  //79 / 6 = 13
    16'b01001111_00000111 : OUT <= 11;  //79 / 7 = 11
    16'b01001111_00001000 : OUT <= 9;  //79 / 8 = 9
    16'b01001111_00001001 : OUT <= 8;  //79 / 9 = 8
    16'b01001111_00001010 : OUT <= 7;  //79 / 10 = 7
    16'b01001111_00001011 : OUT <= 7;  //79 / 11 = 7
    16'b01001111_00001100 : OUT <= 6;  //79 / 12 = 6
    16'b01001111_00001101 : OUT <= 6;  //79 / 13 = 6
    16'b01001111_00001110 : OUT <= 5;  //79 / 14 = 5
    16'b01001111_00001111 : OUT <= 5;  //79 / 15 = 5
    16'b01001111_00010000 : OUT <= 4;  //79 / 16 = 4
    16'b01001111_00010001 : OUT <= 4;  //79 / 17 = 4
    16'b01001111_00010010 : OUT <= 4;  //79 / 18 = 4
    16'b01001111_00010011 : OUT <= 4;  //79 / 19 = 4
    16'b01001111_00010100 : OUT <= 3;  //79 / 20 = 3
    16'b01001111_00010101 : OUT <= 3;  //79 / 21 = 3
    16'b01001111_00010110 : OUT <= 3;  //79 / 22 = 3
    16'b01001111_00010111 : OUT <= 3;  //79 / 23 = 3
    16'b01001111_00011000 : OUT <= 3;  //79 / 24 = 3
    16'b01001111_00011001 : OUT <= 3;  //79 / 25 = 3
    16'b01001111_00011010 : OUT <= 3;  //79 / 26 = 3
    16'b01001111_00011011 : OUT <= 2;  //79 / 27 = 2
    16'b01001111_00011100 : OUT <= 2;  //79 / 28 = 2
    16'b01001111_00011101 : OUT <= 2;  //79 / 29 = 2
    16'b01001111_00011110 : OUT <= 2;  //79 / 30 = 2
    16'b01001111_00011111 : OUT <= 2;  //79 / 31 = 2
    16'b01001111_00100000 : OUT <= 2;  //79 / 32 = 2
    16'b01001111_00100001 : OUT <= 2;  //79 / 33 = 2
    16'b01001111_00100010 : OUT <= 2;  //79 / 34 = 2
    16'b01001111_00100011 : OUT <= 2;  //79 / 35 = 2
    16'b01001111_00100100 : OUT <= 2;  //79 / 36 = 2
    16'b01001111_00100101 : OUT <= 2;  //79 / 37 = 2
    16'b01001111_00100110 : OUT <= 2;  //79 / 38 = 2
    16'b01001111_00100111 : OUT <= 2;  //79 / 39 = 2
    16'b01001111_00101000 : OUT <= 1;  //79 / 40 = 1
    16'b01001111_00101001 : OUT <= 1;  //79 / 41 = 1
    16'b01001111_00101010 : OUT <= 1;  //79 / 42 = 1
    16'b01001111_00101011 : OUT <= 1;  //79 / 43 = 1
    16'b01001111_00101100 : OUT <= 1;  //79 / 44 = 1
    16'b01001111_00101101 : OUT <= 1;  //79 / 45 = 1
    16'b01001111_00101110 : OUT <= 1;  //79 / 46 = 1
    16'b01001111_00101111 : OUT <= 1;  //79 / 47 = 1
    16'b01001111_00110000 : OUT <= 1;  //79 / 48 = 1
    16'b01001111_00110001 : OUT <= 1;  //79 / 49 = 1
    16'b01001111_00110010 : OUT <= 1;  //79 / 50 = 1
    16'b01001111_00110011 : OUT <= 1;  //79 / 51 = 1
    16'b01001111_00110100 : OUT <= 1;  //79 / 52 = 1
    16'b01001111_00110101 : OUT <= 1;  //79 / 53 = 1
    16'b01001111_00110110 : OUT <= 1;  //79 / 54 = 1
    16'b01001111_00110111 : OUT <= 1;  //79 / 55 = 1
    16'b01001111_00111000 : OUT <= 1;  //79 / 56 = 1
    16'b01001111_00111001 : OUT <= 1;  //79 / 57 = 1
    16'b01001111_00111010 : OUT <= 1;  //79 / 58 = 1
    16'b01001111_00111011 : OUT <= 1;  //79 / 59 = 1
    16'b01001111_00111100 : OUT <= 1;  //79 / 60 = 1
    16'b01001111_00111101 : OUT <= 1;  //79 / 61 = 1
    16'b01001111_00111110 : OUT <= 1;  //79 / 62 = 1
    16'b01001111_00111111 : OUT <= 1;  //79 / 63 = 1
    16'b01001111_01000000 : OUT <= 1;  //79 / 64 = 1
    16'b01001111_01000001 : OUT <= 1;  //79 / 65 = 1
    16'b01001111_01000010 : OUT <= 1;  //79 / 66 = 1
    16'b01001111_01000011 : OUT <= 1;  //79 / 67 = 1
    16'b01001111_01000100 : OUT <= 1;  //79 / 68 = 1
    16'b01001111_01000101 : OUT <= 1;  //79 / 69 = 1
    16'b01001111_01000110 : OUT <= 1;  //79 / 70 = 1
    16'b01001111_01000111 : OUT <= 1;  //79 / 71 = 1
    16'b01001111_01001000 : OUT <= 1;  //79 / 72 = 1
    16'b01001111_01001001 : OUT <= 1;  //79 / 73 = 1
    16'b01001111_01001010 : OUT <= 1;  //79 / 74 = 1
    16'b01001111_01001011 : OUT <= 1;  //79 / 75 = 1
    16'b01001111_01001100 : OUT <= 1;  //79 / 76 = 1
    16'b01001111_01001101 : OUT <= 1;  //79 / 77 = 1
    16'b01001111_01001110 : OUT <= 1;  //79 / 78 = 1
    16'b01001111_01001111 : OUT <= 1;  //79 / 79 = 1
    16'b01001111_01010000 : OUT <= 0;  //79 / 80 = 0
    16'b01001111_01010001 : OUT <= 0;  //79 / 81 = 0
    16'b01001111_01010010 : OUT <= 0;  //79 / 82 = 0
    16'b01001111_01010011 : OUT <= 0;  //79 / 83 = 0
    16'b01001111_01010100 : OUT <= 0;  //79 / 84 = 0
    16'b01001111_01010101 : OUT <= 0;  //79 / 85 = 0
    16'b01001111_01010110 : OUT <= 0;  //79 / 86 = 0
    16'b01001111_01010111 : OUT <= 0;  //79 / 87 = 0
    16'b01001111_01011000 : OUT <= 0;  //79 / 88 = 0
    16'b01001111_01011001 : OUT <= 0;  //79 / 89 = 0
    16'b01001111_01011010 : OUT <= 0;  //79 / 90 = 0
    16'b01001111_01011011 : OUT <= 0;  //79 / 91 = 0
    16'b01001111_01011100 : OUT <= 0;  //79 / 92 = 0
    16'b01001111_01011101 : OUT <= 0;  //79 / 93 = 0
    16'b01001111_01011110 : OUT <= 0;  //79 / 94 = 0
    16'b01001111_01011111 : OUT <= 0;  //79 / 95 = 0
    16'b01001111_01100000 : OUT <= 0;  //79 / 96 = 0
    16'b01001111_01100001 : OUT <= 0;  //79 / 97 = 0
    16'b01001111_01100010 : OUT <= 0;  //79 / 98 = 0
    16'b01001111_01100011 : OUT <= 0;  //79 / 99 = 0
    16'b01001111_01100100 : OUT <= 0;  //79 / 100 = 0
    16'b01001111_01100101 : OUT <= 0;  //79 / 101 = 0
    16'b01001111_01100110 : OUT <= 0;  //79 / 102 = 0
    16'b01001111_01100111 : OUT <= 0;  //79 / 103 = 0
    16'b01001111_01101000 : OUT <= 0;  //79 / 104 = 0
    16'b01001111_01101001 : OUT <= 0;  //79 / 105 = 0
    16'b01001111_01101010 : OUT <= 0;  //79 / 106 = 0
    16'b01001111_01101011 : OUT <= 0;  //79 / 107 = 0
    16'b01001111_01101100 : OUT <= 0;  //79 / 108 = 0
    16'b01001111_01101101 : OUT <= 0;  //79 / 109 = 0
    16'b01001111_01101110 : OUT <= 0;  //79 / 110 = 0
    16'b01001111_01101111 : OUT <= 0;  //79 / 111 = 0
    16'b01001111_01110000 : OUT <= 0;  //79 / 112 = 0
    16'b01001111_01110001 : OUT <= 0;  //79 / 113 = 0
    16'b01001111_01110010 : OUT <= 0;  //79 / 114 = 0
    16'b01001111_01110011 : OUT <= 0;  //79 / 115 = 0
    16'b01001111_01110100 : OUT <= 0;  //79 / 116 = 0
    16'b01001111_01110101 : OUT <= 0;  //79 / 117 = 0
    16'b01001111_01110110 : OUT <= 0;  //79 / 118 = 0
    16'b01001111_01110111 : OUT <= 0;  //79 / 119 = 0
    16'b01001111_01111000 : OUT <= 0;  //79 / 120 = 0
    16'b01001111_01111001 : OUT <= 0;  //79 / 121 = 0
    16'b01001111_01111010 : OUT <= 0;  //79 / 122 = 0
    16'b01001111_01111011 : OUT <= 0;  //79 / 123 = 0
    16'b01001111_01111100 : OUT <= 0;  //79 / 124 = 0
    16'b01001111_01111101 : OUT <= 0;  //79 / 125 = 0
    16'b01001111_01111110 : OUT <= 0;  //79 / 126 = 0
    16'b01001111_01111111 : OUT <= 0;  //79 / 127 = 0
    16'b01001111_10000000 : OUT <= 0;  //79 / 128 = 0
    16'b01001111_10000001 : OUT <= 0;  //79 / 129 = 0
    16'b01001111_10000010 : OUT <= 0;  //79 / 130 = 0
    16'b01001111_10000011 : OUT <= 0;  //79 / 131 = 0
    16'b01001111_10000100 : OUT <= 0;  //79 / 132 = 0
    16'b01001111_10000101 : OUT <= 0;  //79 / 133 = 0
    16'b01001111_10000110 : OUT <= 0;  //79 / 134 = 0
    16'b01001111_10000111 : OUT <= 0;  //79 / 135 = 0
    16'b01001111_10001000 : OUT <= 0;  //79 / 136 = 0
    16'b01001111_10001001 : OUT <= 0;  //79 / 137 = 0
    16'b01001111_10001010 : OUT <= 0;  //79 / 138 = 0
    16'b01001111_10001011 : OUT <= 0;  //79 / 139 = 0
    16'b01001111_10001100 : OUT <= 0;  //79 / 140 = 0
    16'b01001111_10001101 : OUT <= 0;  //79 / 141 = 0
    16'b01001111_10001110 : OUT <= 0;  //79 / 142 = 0
    16'b01001111_10001111 : OUT <= 0;  //79 / 143 = 0
    16'b01001111_10010000 : OUT <= 0;  //79 / 144 = 0
    16'b01001111_10010001 : OUT <= 0;  //79 / 145 = 0
    16'b01001111_10010010 : OUT <= 0;  //79 / 146 = 0
    16'b01001111_10010011 : OUT <= 0;  //79 / 147 = 0
    16'b01001111_10010100 : OUT <= 0;  //79 / 148 = 0
    16'b01001111_10010101 : OUT <= 0;  //79 / 149 = 0
    16'b01001111_10010110 : OUT <= 0;  //79 / 150 = 0
    16'b01001111_10010111 : OUT <= 0;  //79 / 151 = 0
    16'b01001111_10011000 : OUT <= 0;  //79 / 152 = 0
    16'b01001111_10011001 : OUT <= 0;  //79 / 153 = 0
    16'b01001111_10011010 : OUT <= 0;  //79 / 154 = 0
    16'b01001111_10011011 : OUT <= 0;  //79 / 155 = 0
    16'b01001111_10011100 : OUT <= 0;  //79 / 156 = 0
    16'b01001111_10011101 : OUT <= 0;  //79 / 157 = 0
    16'b01001111_10011110 : OUT <= 0;  //79 / 158 = 0
    16'b01001111_10011111 : OUT <= 0;  //79 / 159 = 0
    16'b01001111_10100000 : OUT <= 0;  //79 / 160 = 0
    16'b01001111_10100001 : OUT <= 0;  //79 / 161 = 0
    16'b01001111_10100010 : OUT <= 0;  //79 / 162 = 0
    16'b01001111_10100011 : OUT <= 0;  //79 / 163 = 0
    16'b01001111_10100100 : OUT <= 0;  //79 / 164 = 0
    16'b01001111_10100101 : OUT <= 0;  //79 / 165 = 0
    16'b01001111_10100110 : OUT <= 0;  //79 / 166 = 0
    16'b01001111_10100111 : OUT <= 0;  //79 / 167 = 0
    16'b01001111_10101000 : OUT <= 0;  //79 / 168 = 0
    16'b01001111_10101001 : OUT <= 0;  //79 / 169 = 0
    16'b01001111_10101010 : OUT <= 0;  //79 / 170 = 0
    16'b01001111_10101011 : OUT <= 0;  //79 / 171 = 0
    16'b01001111_10101100 : OUT <= 0;  //79 / 172 = 0
    16'b01001111_10101101 : OUT <= 0;  //79 / 173 = 0
    16'b01001111_10101110 : OUT <= 0;  //79 / 174 = 0
    16'b01001111_10101111 : OUT <= 0;  //79 / 175 = 0
    16'b01001111_10110000 : OUT <= 0;  //79 / 176 = 0
    16'b01001111_10110001 : OUT <= 0;  //79 / 177 = 0
    16'b01001111_10110010 : OUT <= 0;  //79 / 178 = 0
    16'b01001111_10110011 : OUT <= 0;  //79 / 179 = 0
    16'b01001111_10110100 : OUT <= 0;  //79 / 180 = 0
    16'b01001111_10110101 : OUT <= 0;  //79 / 181 = 0
    16'b01001111_10110110 : OUT <= 0;  //79 / 182 = 0
    16'b01001111_10110111 : OUT <= 0;  //79 / 183 = 0
    16'b01001111_10111000 : OUT <= 0;  //79 / 184 = 0
    16'b01001111_10111001 : OUT <= 0;  //79 / 185 = 0
    16'b01001111_10111010 : OUT <= 0;  //79 / 186 = 0
    16'b01001111_10111011 : OUT <= 0;  //79 / 187 = 0
    16'b01001111_10111100 : OUT <= 0;  //79 / 188 = 0
    16'b01001111_10111101 : OUT <= 0;  //79 / 189 = 0
    16'b01001111_10111110 : OUT <= 0;  //79 / 190 = 0
    16'b01001111_10111111 : OUT <= 0;  //79 / 191 = 0
    16'b01001111_11000000 : OUT <= 0;  //79 / 192 = 0
    16'b01001111_11000001 : OUT <= 0;  //79 / 193 = 0
    16'b01001111_11000010 : OUT <= 0;  //79 / 194 = 0
    16'b01001111_11000011 : OUT <= 0;  //79 / 195 = 0
    16'b01001111_11000100 : OUT <= 0;  //79 / 196 = 0
    16'b01001111_11000101 : OUT <= 0;  //79 / 197 = 0
    16'b01001111_11000110 : OUT <= 0;  //79 / 198 = 0
    16'b01001111_11000111 : OUT <= 0;  //79 / 199 = 0
    16'b01001111_11001000 : OUT <= 0;  //79 / 200 = 0
    16'b01001111_11001001 : OUT <= 0;  //79 / 201 = 0
    16'b01001111_11001010 : OUT <= 0;  //79 / 202 = 0
    16'b01001111_11001011 : OUT <= 0;  //79 / 203 = 0
    16'b01001111_11001100 : OUT <= 0;  //79 / 204 = 0
    16'b01001111_11001101 : OUT <= 0;  //79 / 205 = 0
    16'b01001111_11001110 : OUT <= 0;  //79 / 206 = 0
    16'b01001111_11001111 : OUT <= 0;  //79 / 207 = 0
    16'b01001111_11010000 : OUT <= 0;  //79 / 208 = 0
    16'b01001111_11010001 : OUT <= 0;  //79 / 209 = 0
    16'b01001111_11010010 : OUT <= 0;  //79 / 210 = 0
    16'b01001111_11010011 : OUT <= 0;  //79 / 211 = 0
    16'b01001111_11010100 : OUT <= 0;  //79 / 212 = 0
    16'b01001111_11010101 : OUT <= 0;  //79 / 213 = 0
    16'b01001111_11010110 : OUT <= 0;  //79 / 214 = 0
    16'b01001111_11010111 : OUT <= 0;  //79 / 215 = 0
    16'b01001111_11011000 : OUT <= 0;  //79 / 216 = 0
    16'b01001111_11011001 : OUT <= 0;  //79 / 217 = 0
    16'b01001111_11011010 : OUT <= 0;  //79 / 218 = 0
    16'b01001111_11011011 : OUT <= 0;  //79 / 219 = 0
    16'b01001111_11011100 : OUT <= 0;  //79 / 220 = 0
    16'b01001111_11011101 : OUT <= 0;  //79 / 221 = 0
    16'b01001111_11011110 : OUT <= 0;  //79 / 222 = 0
    16'b01001111_11011111 : OUT <= 0;  //79 / 223 = 0
    16'b01001111_11100000 : OUT <= 0;  //79 / 224 = 0
    16'b01001111_11100001 : OUT <= 0;  //79 / 225 = 0
    16'b01001111_11100010 : OUT <= 0;  //79 / 226 = 0
    16'b01001111_11100011 : OUT <= 0;  //79 / 227 = 0
    16'b01001111_11100100 : OUT <= 0;  //79 / 228 = 0
    16'b01001111_11100101 : OUT <= 0;  //79 / 229 = 0
    16'b01001111_11100110 : OUT <= 0;  //79 / 230 = 0
    16'b01001111_11100111 : OUT <= 0;  //79 / 231 = 0
    16'b01001111_11101000 : OUT <= 0;  //79 / 232 = 0
    16'b01001111_11101001 : OUT <= 0;  //79 / 233 = 0
    16'b01001111_11101010 : OUT <= 0;  //79 / 234 = 0
    16'b01001111_11101011 : OUT <= 0;  //79 / 235 = 0
    16'b01001111_11101100 : OUT <= 0;  //79 / 236 = 0
    16'b01001111_11101101 : OUT <= 0;  //79 / 237 = 0
    16'b01001111_11101110 : OUT <= 0;  //79 / 238 = 0
    16'b01001111_11101111 : OUT <= 0;  //79 / 239 = 0
    16'b01001111_11110000 : OUT <= 0;  //79 / 240 = 0
    16'b01001111_11110001 : OUT <= 0;  //79 / 241 = 0
    16'b01001111_11110010 : OUT <= 0;  //79 / 242 = 0
    16'b01001111_11110011 : OUT <= 0;  //79 / 243 = 0
    16'b01001111_11110100 : OUT <= 0;  //79 / 244 = 0
    16'b01001111_11110101 : OUT <= 0;  //79 / 245 = 0
    16'b01001111_11110110 : OUT <= 0;  //79 / 246 = 0
    16'b01001111_11110111 : OUT <= 0;  //79 / 247 = 0
    16'b01001111_11111000 : OUT <= 0;  //79 / 248 = 0
    16'b01001111_11111001 : OUT <= 0;  //79 / 249 = 0
    16'b01001111_11111010 : OUT <= 0;  //79 / 250 = 0
    16'b01001111_11111011 : OUT <= 0;  //79 / 251 = 0
    16'b01001111_11111100 : OUT <= 0;  //79 / 252 = 0
    16'b01001111_11111101 : OUT <= 0;  //79 / 253 = 0
    16'b01001111_11111110 : OUT <= 0;  //79 / 254 = 0
    16'b01001111_11111111 : OUT <= 0;  //79 / 255 = 0
    16'b01010000_00000000 : OUT <= 0;  //80 / 0 = 0
    16'b01010000_00000001 : OUT <= 80;  //80 / 1 = 80
    16'b01010000_00000010 : OUT <= 40;  //80 / 2 = 40
    16'b01010000_00000011 : OUT <= 26;  //80 / 3 = 26
    16'b01010000_00000100 : OUT <= 20;  //80 / 4 = 20
    16'b01010000_00000101 : OUT <= 16;  //80 / 5 = 16
    16'b01010000_00000110 : OUT <= 13;  //80 / 6 = 13
    16'b01010000_00000111 : OUT <= 11;  //80 / 7 = 11
    16'b01010000_00001000 : OUT <= 10;  //80 / 8 = 10
    16'b01010000_00001001 : OUT <= 8;  //80 / 9 = 8
    16'b01010000_00001010 : OUT <= 8;  //80 / 10 = 8
    16'b01010000_00001011 : OUT <= 7;  //80 / 11 = 7
    16'b01010000_00001100 : OUT <= 6;  //80 / 12 = 6
    16'b01010000_00001101 : OUT <= 6;  //80 / 13 = 6
    16'b01010000_00001110 : OUT <= 5;  //80 / 14 = 5
    16'b01010000_00001111 : OUT <= 5;  //80 / 15 = 5
    16'b01010000_00010000 : OUT <= 5;  //80 / 16 = 5
    16'b01010000_00010001 : OUT <= 4;  //80 / 17 = 4
    16'b01010000_00010010 : OUT <= 4;  //80 / 18 = 4
    16'b01010000_00010011 : OUT <= 4;  //80 / 19 = 4
    16'b01010000_00010100 : OUT <= 4;  //80 / 20 = 4
    16'b01010000_00010101 : OUT <= 3;  //80 / 21 = 3
    16'b01010000_00010110 : OUT <= 3;  //80 / 22 = 3
    16'b01010000_00010111 : OUT <= 3;  //80 / 23 = 3
    16'b01010000_00011000 : OUT <= 3;  //80 / 24 = 3
    16'b01010000_00011001 : OUT <= 3;  //80 / 25 = 3
    16'b01010000_00011010 : OUT <= 3;  //80 / 26 = 3
    16'b01010000_00011011 : OUT <= 2;  //80 / 27 = 2
    16'b01010000_00011100 : OUT <= 2;  //80 / 28 = 2
    16'b01010000_00011101 : OUT <= 2;  //80 / 29 = 2
    16'b01010000_00011110 : OUT <= 2;  //80 / 30 = 2
    16'b01010000_00011111 : OUT <= 2;  //80 / 31 = 2
    16'b01010000_00100000 : OUT <= 2;  //80 / 32 = 2
    16'b01010000_00100001 : OUT <= 2;  //80 / 33 = 2
    16'b01010000_00100010 : OUT <= 2;  //80 / 34 = 2
    16'b01010000_00100011 : OUT <= 2;  //80 / 35 = 2
    16'b01010000_00100100 : OUT <= 2;  //80 / 36 = 2
    16'b01010000_00100101 : OUT <= 2;  //80 / 37 = 2
    16'b01010000_00100110 : OUT <= 2;  //80 / 38 = 2
    16'b01010000_00100111 : OUT <= 2;  //80 / 39 = 2
    16'b01010000_00101000 : OUT <= 2;  //80 / 40 = 2
    16'b01010000_00101001 : OUT <= 1;  //80 / 41 = 1
    16'b01010000_00101010 : OUT <= 1;  //80 / 42 = 1
    16'b01010000_00101011 : OUT <= 1;  //80 / 43 = 1
    16'b01010000_00101100 : OUT <= 1;  //80 / 44 = 1
    16'b01010000_00101101 : OUT <= 1;  //80 / 45 = 1
    16'b01010000_00101110 : OUT <= 1;  //80 / 46 = 1
    16'b01010000_00101111 : OUT <= 1;  //80 / 47 = 1
    16'b01010000_00110000 : OUT <= 1;  //80 / 48 = 1
    16'b01010000_00110001 : OUT <= 1;  //80 / 49 = 1
    16'b01010000_00110010 : OUT <= 1;  //80 / 50 = 1
    16'b01010000_00110011 : OUT <= 1;  //80 / 51 = 1
    16'b01010000_00110100 : OUT <= 1;  //80 / 52 = 1
    16'b01010000_00110101 : OUT <= 1;  //80 / 53 = 1
    16'b01010000_00110110 : OUT <= 1;  //80 / 54 = 1
    16'b01010000_00110111 : OUT <= 1;  //80 / 55 = 1
    16'b01010000_00111000 : OUT <= 1;  //80 / 56 = 1
    16'b01010000_00111001 : OUT <= 1;  //80 / 57 = 1
    16'b01010000_00111010 : OUT <= 1;  //80 / 58 = 1
    16'b01010000_00111011 : OUT <= 1;  //80 / 59 = 1
    16'b01010000_00111100 : OUT <= 1;  //80 / 60 = 1
    16'b01010000_00111101 : OUT <= 1;  //80 / 61 = 1
    16'b01010000_00111110 : OUT <= 1;  //80 / 62 = 1
    16'b01010000_00111111 : OUT <= 1;  //80 / 63 = 1
    16'b01010000_01000000 : OUT <= 1;  //80 / 64 = 1
    16'b01010000_01000001 : OUT <= 1;  //80 / 65 = 1
    16'b01010000_01000010 : OUT <= 1;  //80 / 66 = 1
    16'b01010000_01000011 : OUT <= 1;  //80 / 67 = 1
    16'b01010000_01000100 : OUT <= 1;  //80 / 68 = 1
    16'b01010000_01000101 : OUT <= 1;  //80 / 69 = 1
    16'b01010000_01000110 : OUT <= 1;  //80 / 70 = 1
    16'b01010000_01000111 : OUT <= 1;  //80 / 71 = 1
    16'b01010000_01001000 : OUT <= 1;  //80 / 72 = 1
    16'b01010000_01001001 : OUT <= 1;  //80 / 73 = 1
    16'b01010000_01001010 : OUT <= 1;  //80 / 74 = 1
    16'b01010000_01001011 : OUT <= 1;  //80 / 75 = 1
    16'b01010000_01001100 : OUT <= 1;  //80 / 76 = 1
    16'b01010000_01001101 : OUT <= 1;  //80 / 77 = 1
    16'b01010000_01001110 : OUT <= 1;  //80 / 78 = 1
    16'b01010000_01001111 : OUT <= 1;  //80 / 79 = 1
    16'b01010000_01010000 : OUT <= 1;  //80 / 80 = 1
    16'b01010000_01010001 : OUT <= 0;  //80 / 81 = 0
    16'b01010000_01010010 : OUT <= 0;  //80 / 82 = 0
    16'b01010000_01010011 : OUT <= 0;  //80 / 83 = 0
    16'b01010000_01010100 : OUT <= 0;  //80 / 84 = 0
    16'b01010000_01010101 : OUT <= 0;  //80 / 85 = 0
    16'b01010000_01010110 : OUT <= 0;  //80 / 86 = 0
    16'b01010000_01010111 : OUT <= 0;  //80 / 87 = 0
    16'b01010000_01011000 : OUT <= 0;  //80 / 88 = 0
    16'b01010000_01011001 : OUT <= 0;  //80 / 89 = 0
    16'b01010000_01011010 : OUT <= 0;  //80 / 90 = 0
    16'b01010000_01011011 : OUT <= 0;  //80 / 91 = 0
    16'b01010000_01011100 : OUT <= 0;  //80 / 92 = 0
    16'b01010000_01011101 : OUT <= 0;  //80 / 93 = 0
    16'b01010000_01011110 : OUT <= 0;  //80 / 94 = 0
    16'b01010000_01011111 : OUT <= 0;  //80 / 95 = 0
    16'b01010000_01100000 : OUT <= 0;  //80 / 96 = 0
    16'b01010000_01100001 : OUT <= 0;  //80 / 97 = 0
    16'b01010000_01100010 : OUT <= 0;  //80 / 98 = 0
    16'b01010000_01100011 : OUT <= 0;  //80 / 99 = 0
    16'b01010000_01100100 : OUT <= 0;  //80 / 100 = 0
    16'b01010000_01100101 : OUT <= 0;  //80 / 101 = 0
    16'b01010000_01100110 : OUT <= 0;  //80 / 102 = 0
    16'b01010000_01100111 : OUT <= 0;  //80 / 103 = 0
    16'b01010000_01101000 : OUT <= 0;  //80 / 104 = 0
    16'b01010000_01101001 : OUT <= 0;  //80 / 105 = 0
    16'b01010000_01101010 : OUT <= 0;  //80 / 106 = 0
    16'b01010000_01101011 : OUT <= 0;  //80 / 107 = 0
    16'b01010000_01101100 : OUT <= 0;  //80 / 108 = 0
    16'b01010000_01101101 : OUT <= 0;  //80 / 109 = 0
    16'b01010000_01101110 : OUT <= 0;  //80 / 110 = 0
    16'b01010000_01101111 : OUT <= 0;  //80 / 111 = 0
    16'b01010000_01110000 : OUT <= 0;  //80 / 112 = 0
    16'b01010000_01110001 : OUT <= 0;  //80 / 113 = 0
    16'b01010000_01110010 : OUT <= 0;  //80 / 114 = 0
    16'b01010000_01110011 : OUT <= 0;  //80 / 115 = 0
    16'b01010000_01110100 : OUT <= 0;  //80 / 116 = 0
    16'b01010000_01110101 : OUT <= 0;  //80 / 117 = 0
    16'b01010000_01110110 : OUT <= 0;  //80 / 118 = 0
    16'b01010000_01110111 : OUT <= 0;  //80 / 119 = 0
    16'b01010000_01111000 : OUT <= 0;  //80 / 120 = 0
    16'b01010000_01111001 : OUT <= 0;  //80 / 121 = 0
    16'b01010000_01111010 : OUT <= 0;  //80 / 122 = 0
    16'b01010000_01111011 : OUT <= 0;  //80 / 123 = 0
    16'b01010000_01111100 : OUT <= 0;  //80 / 124 = 0
    16'b01010000_01111101 : OUT <= 0;  //80 / 125 = 0
    16'b01010000_01111110 : OUT <= 0;  //80 / 126 = 0
    16'b01010000_01111111 : OUT <= 0;  //80 / 127 = 0
    16'b01010000_10000000 : OUT <= 0;  //80 / 128 = 0
    16'b01010000_10000001 : OUT <= 0;  //80 / 129 = 0
    16'b01010000_10000010 : OUT <= 0;  //80 / 130 = 0
    16'b01010000_10000011 : OUT <= 0;  //80 / 131 = 0
    16'b01010000_10000100 : OUT <= 0;  //80 / 132 = 0
    16'b01010000_10000101 : OUT <= 0;  //80 / 133 = 0
    16'b01010000_10000110 : OUT <= 0;  //80 / 134 = 0
    16'b01010000_10000111 : OUT <= 0;  //80 / 135 = 0
    16'b01010000_10001000 : OUT <= 0;  //80 / 136 = 0
    16'b01010000_10001001 : OUT <= 0;  //80 / 137 = 0
    16'b01010000_10001010 : OUT <= 0;  //80 / 138 = 0
    16'b01010000_10001011 : OUT <= 0;  //80 / 139 = 0
    16'b01010000_10001100 : OUT <= 0;  //80 / 140 = 0
    16'b01010000_10001101 : OUT <= 0;  //80 / 141 = 0
    16'b01010000_10001110 : OUT <= 0;  //80 / 142 = 0
    16'b01010000_10001111 : OUT <= 0;  //80 / 143 = 0
    16'b01010000_10010000 : OUT <= 0;  //80 / 144 = 0
    16'b01010000_10010001 : OUT <= 0;  //80 / 145 = 0
    16'b01010000_10010010 : OUT <= 0;  //80 / 146 = 0
    16'b01010000_10010011 : OUT <= 0;  //80 / 147 = 0
    16'b01010000_10010100 : OUT <= 0;  //80 / 148 = 0
    16'b01010000_10010101 : OUT <= 0;  //80 / 149 = 0
    16'b01010000_10010110 : OUT <= 0;  //80 / 150 = 0
    16'b01010000_10010111 : OUT <= 0;  //80 / 151 = 0
    16'b01010000_10011000 : OUT <= 0;  //80 / 152 = 0
    16'b01010000_10011001 : OUT <= 0;  //80 / 153 = 0
    16'b01010000_10011010 : OUT <= 0;  //80 / 154 = 0
    16'b01010000_10011011 : OUT <= 0;  //80 / 155 = 0
    16'b01010000_10011100 : OUT <= 0;  //80 / 156 = 0
    16'b01010000_10011101 : OUT <= 0;  //80 / 157 = 0
    16'b01010000_10011110 : OUT <= 0;  //80 / 158 = 0
    16'b01010000_10011111 : OUT <= 0;  //80 / 159 = 0
    16'b01010000_10100000 : OUT <= 0;  //80 / 160 = 0
    16'b01010000_10100001 : OUT <= 0;  //80 / 161 = 0
    16'b01010000_10100010 : OUT <= 0;  //80 / 162 = 0
    16'b01010000_10100011 : OUT <= 0;  //80 / 163 = 0
    16'b01010000_10100100 : OUT <= 0;  //80 / 164 = 0
    16'b01010000_10100101 : OUT <= 0;  //80 / 165 = 0
    16'b01010000_10100110 : OUT <= 0;  //80 / 166 = 0
    16'b01010000_10100111 : OUT <= 0;  //80 / 167 = 0
    16'b01010000_10101000 : OUT <= 0;  //80 / 168 = 0
    16'b01010000_10101001 : OUT <= 0;  //80 / 169 = 0
    16'b01010000_10101010 : OUT <= 0;  //80 / 170 = 0
    16'b01010000_10101011 : OUT <= 0;  //80 / 171 = 0
    16'b01010000_10101100 : OUT <= 0;  //80 / 172 = 0
    16'b01010000_10101101 : OUT <= 0;  //80 / 173 = 0
    16'b01010000_10101110 : OUT <= 0;  //80 / 174 = 0
    16'b01010000_10101111 : OUT <= 0;  //80 / 175 = 0
    16'b01010000_10110000 : OUT <= 0;  //80 / 176 = 0
    16'b01010000_10110001 : OUT <= 0;  //80 / 177 = 0
    16'b01010000_10110010 : OUT <= 0;  //80 / 178 = 0
    16'b01010000_10110011 : OUT <= 0;  //80 / 179 = 0
    16'b01010000_10110100 : OUT <= 0;  //80 / 180 = 0
    16'b01010000_10110101 : OUT <= 0;  //80 / 181 = 0
    16'b01010000_10110110 : OUT <= 0;  //80 / 182 = 0
    16'b01010000_10110111 : OUT <= 0;  //80 / 183 = 0
    16'b01010000_10111000 : OUT <= 0;  //80 / 184 = 0
    16'b01010000_10111001 : OUT <= 0;  //80 / 185 = 0
    16'b01010000_10111010 : OUT <= 0;  //80 / 186 = 0
    16'b01010000_10111011 : OUT <= 0;  //80 / 187 = 0
    16'b01010000_10111100 : OUT <= 0;  //80 / 188 = 0
    16'b01010000_10111101 : OUT <= 0;  //80 / 189 = 0
    16'b01010000_10111110 : OUT <= 0;  //80 / 190 = 0
    16'b01010000_10111111 : OUT <= 0;  //80 / 191 = 0
    16'b01010000_11000000 : OUT <= 0;  //80 / 192 = 0
    16'b01010000_11000001 : OUT <= 0;  //80 / 193 = 0
    16'b01010000_11000010 : OUT <= 0;  //80 / 194 = 0
    16'b01010000_11000011 : OUT <= 0;  //80 / 195 = 0
    16'b01010000_11000100 : OUT <= 0;  //80 / 196 = 0
    16'b01010000_11000101 : OUT <= 0;  //80 / 197 = 0
    16'b01010000_11000110 : OUT <= 0;  //80 / 198 = 0
    16'b01010000_11000111 : OUT <= 0;  //80 / 199 = 0
    16'b01010000_11001000 : OUT <= 0;  //80 / 200 = 0
    16'b01010000_11001001 : OUT <= 0;  //80 / 201 = 0
    16'b01010000_11001010 : OUT <= 0;  //80 / 202 = 0
    16'b01010000_11001011 : OUT <= 0;  //80 / 203 = 0
    16'b01010000_11001100 : OUT <= 0;  //80 / 204 = 0
    16'b01010000_11001101 : OUT <= 0;  //80 / 205 = 0
    16'b01010000_11001110 : OUT <= 0;  //80 / 206 = 0
    16'b01010000_11001111 : OUT <= 0;  //80 / 207 = 0
    16'b01010000_11010000 : OUT <= 0;  //80 / 208 = 0
    16'b01010000_11010001 : OUT <= 0;  //80 / 209 = 0
    16'b01010000_11010010 : OUT <= 0;  //80 / 210 = 0
    16'b01010000_11010011 : OUT <= 0;  //80 / 211 = 0
    16'b01010000_11010100 : OUT <= 0;  //80 / 212 = 0
    16'b01010000_11010101 : OUT <= 0;  //80 / 213 = 0
    16'b01010000_11010110 : OUT <= 0;  //80 / 214 = 0
    16'b01010000_11010111 : OUT <= 0;  //80 / 215 = 0
    16'b01010000_11011000 : OUT <= 0;  //80 / 216 = 0
    16'b01010000_11011001 : OUT <= 0;  //80 / 217 = 0
    16'b01010000_11011010 : OUT <= 0;  //80 / 218 = 0
    16'b01010000_11011011 : OUT <= 0;  //80 / 219 = 0
    16'b01010000_11011100 : OUT <= 0;  //80 / 220 = 0
    16'b01010000_11011101 : OUT <= 0;  //80 / 221 = 0
    16'b01010000_11011110 : OUT <= 0;  //80 / 222 = 0
    16'b01010000_11011111 : OUT <= 0;  //80 / 223 = 0
    16'b01010000_11100000 : OUT <= 0;  //80 / 224 = 0
    16'b01010000_11100001 : OUT <= 0;  //80 / 225 = 0
    16'b01010000_11100010 : OUT <= 0;  //80 / 226 = 0
    16'b01010000_11100011 : OUT <= 0;  //80 / 227 = 0
    16'b01010000_11100100 : OUT <= 0;  //80 / 228 = 0
    16'b01010000_11100101 : OUT <= 0;  //80 / 229 = 0
    16'b01010000_11100110 : OUT <= 0;  //80 / 230 = 0
    16'b01010000_11100111 : OUT <= 0;  //80 / 231 = 0
    16'b01010000_11101000 : OUT <= 0;  //80 / 232 = 0
    16'b01010000_11101001 : OUT <= 0;  //80 / 233 = 0
    16'b01010000_11101010 : OUT <= 0;  //80 / 234 = 0
    16'b01010000_11101011 : OUT <= 0;  //80 / 235 = 0
    16'b01010000_11101100 : OUT <= 0;  //80 / 236 = 0
    16'b01010000_11101101 : OUT <= 0;  //80 / 237 = 0
    16'b01010000_11101110 : OUT <= 0;  //80 / 238 = 0
    16'b01010000_11101111 : OUT <= 0;  //80 / 239 = 0
    16'b01010000_11110000 : OUT <= 0;  //80 / 240 = 0
    16'b01010000_11110001 : OUT <= 0;  //80 / 241 = 0
    16'b01010000_11110010 : OUT <= 0;  //80 / 242 = 0
    16'b01010000_11110011 : OUT <= 0;  //80 / 243 = 0
    16'b01010000_11110100 : OUT <= 0;  //80 / 244 = 0
    16'b01010000_11110101 : OUT <= 0;  //80 / 245 = 0
    16'b01010000_11110110 : OUT <= 0;  //80 / 246 = 0
    16'b01010000_11110111 : OUT <= 0;  //80 / 247 = 0
    16'b01010000_11111000 : OUT <= 0;  //80 / 248 = 0
    16'b01010000_11111001 : OUT <= 0;  //80 / 249 = 0
    16'b01010000_11111010 : OUT <= 0;  //80 / 250 = 0
    16'b01010000_11111011 : OUT <= 0;  //80 / 251 = 0
    16'b01010000_11111100 : OUT <= 0;  //80 / 252 = 0
    16'b01010000_11111101 : OUT <= 0;  //80 / 253 = 0
    16'b01010000_11111110 : OUT <= 0;  //80 / 254 = 0
    16'b01010000_11111111 : OUT <= 0;  //80 / 255 = 0
    16'b01010001_00000000 : OUT <= 0;  //81 / 0 = 0
    16'b01010001_00000001 : OUT <= 81;  //81 / 1 = 81
    16'b01010001_00000010 : OUT <= 40;  //81 / 2 = 40
    16'b01010001_00000011 : OUT <= 27;  //81 / 3 = 27
    16'b01010001_00000100 : OUT <= 20;  //81 / 4 = 20
    16'b01010001_00000101 : OUT <= 16;  //81 / 5 = 16
    16'b01010001_00000110 : OUT <= 13;  //81 / 6 = 13
    16'b01010001_00000111 : OUT <= 11;  //81 / 7 = 11
    16'b01010001_00001000 : OUT <= 10;  //81 / 8 = 10
    16'b01010001_00001001 : OUT <= 9;  //81 / 9 = 9
    16'b01010001_00001010 : OUT <= 8;  //81 / 10 = 8
    16'b01010001_00001011 : OUT <= 7;  //81 / 11 = 7
    16'b01010001_00001100 : OUT <= 6;  //81 / 12 = 6
    16'b01010001_00001101 : OUT <= 6;  //81 / 13 = 6
    16'b01010001_00001110 : OUT <= 5;  //81 / 14 = 5
    16'b01010001_00001111 : OUT <= 5;  //81 / 15 = 5
    16'b01010001_00010000 : OUT <= 5;  //81 / 16 = 5
    16'b01010001_00010001 : OUT <= 4;  //81 / 17 = 4
    16'b01010001_00010010 : OUT <= 4;  //81 / 18 = 4
    16'b01010001_00010011 : OUT <= 4;  //81 / 19 = 4
    16'b01010001_00010100 : OUT <= 4;  //81 / 20 = 4
    16'b01010001_00010101 : OUT <= 3;  //81 / 21 = 3
    16'b01010001_00010110 : OUT <= 3;  //81 / 22 = 3
    16'b01010001_00010111 : OUT <= 3;  //81 / 23 = 3
    16'b01010001_00011000 : OUT <= 3;  //81 / 24 = 3
    16'b01010001_00011001 : OUT <= 3;  //81 / 25 = 3
    16'b01010001_00011010 : OUT <= 3;  //81 / 26 = 3
    16'b01010001_00011011 : OUT <= 3;  //81 / 27 = 3
    16'b01010001_00011100 : OUT <= 2;  //81 / 28 = 2
    16'b01010001_00011101 : OUT <= 2;  //81 / 29 = 2
    16'b01010001_00011110 : OUT <= 2;  //81 / 30 = 2
    16'b01010001_00011111 : OUT <= 2;  //81 / 31 = 2
    16'b01010001_00100000 : OUT <= 2;  //81 / 32 = 2
    16'b01010001_00100001 : OUT <= 2;  //81 / 33 = 2
    16'b01010001_00100010 : OUT <= 2;  //81 / 34 = 2
    16'b01010001_00100011 : OUT <= 2;  //81 / 35 = 2
    16'b01010001_00100100 : OUT <= 2;  //81 / 36 = 2
    16'b01010001_00100101 : OUT <= 2;  //81 / 37 = 2
    16'b01010001_00100110 : OUT <= 2;  //81 / 38 = 2
    16'b01010001_00100111 : OUT <= 2;  //81 / 39 = 2
    16'b01010001_00101000 : OUT <= 2;  //81 / 40 = 2
    16'b01010001_00101001 : OUT <= 1;  //81 / 41 = 1
    16'b01010001_00101010 : OUT <= 1;  //81 / 42 = 1
    16'b01010001_00101011 : OUT <= 1;  //81 / 43 = 1
    16'b01010001_00101100 : OUT <= 1;  //81 / 44 = 1
    16'b01010001_00101101 : OUT <= 1;  //81 / 45 = 1
    16'b01010001_00101110 : OUT <= 1;  //81 / 46 = 1
    16'b01010001_00101111 : OUT <= 1;  //81 / 47 = 1
    16'b01010001_00110000 : OUT <= 1;  //81 / 48 = 1
    16'b01010001_00110001 : OUT <= 1;  //81 / 49 = 1
    16'b01010001_00110010 : OUT <= 1;  //81 / 50 = 1
    16'b01010001_00110011 : OUT <= 1;  //81 / 51 = 1
    16'b01010001_00110100 : OUT <= 1;  //81 / 52 = 1
    16'b01010001_00110101 : OUT <= 1;  //81 / 53 = 1
    16'b01010001_00110110 : OUT <= 1;  //81 / 54 = 1
    16'b01010001_00110111 : OUT <= 1;  //81 / 55 = 1
    16'b01010001_00111000 : OUT <= 1;  //81 / 56 = 1
    16'b01010001_00111001 : OUT <= 1;  //81 / 57 = 1
    16'b01010001_00111010 : OUT <= 1;  //81 / 58 = 1
    16'b01010001_00111011 : OUT <= 1;  //81 / 59 = 1
    16'b01010001_00111100 : OUT <= 1;  //81 / 60 = 1
    16'b01010001_00111101 : OUT <= 1;  //81 / 61 = 1
    16'b01010001_00111110 : OUT <= 1;  //81 / 62 = 1
    16'b01010001_00111111 : OUT <= 1;  //81 / 63 = 1
    16'b01010001_01000000 : OUT <= 1;  //81 / 64 = 1
    16'b01010001_01000001 : OUT <= 1;  //81 / 65 = 1
    16'b01010001_01000010 : OUT <= 1;  //81 / 66 = 1
    16'b01010001_01000011 : OUT <= 1;  //81 / 67 = 1
    16'b01010001_01000100 : OUT <= 1;  //81 / 68 = 1
    16'b01010001_01000101 : OUT <= 1;  //81 / 69 = 1
    16'b01010001_01000110 : OUT <= 1;  //81 / 70 = 1
    16'b01010001_01000111 : OUT <= 1;  //81 / 71 = 1
    16'b01010001_01001000 : OUT <= 1;  //81 / 72 = 1
    16'b01010001_01001001 : OUT <= 1;  //81 / 73 = 1
    16'b01010001_01001010 : OUT <= 1;  //81 / 74 = 1
    16'b01010001_01001011 : OUT <= 1;  //81 / 75 = 1
    16'b01010001_01001100 : OUT <= 1;  //81 / 76 = 1
    16'b01010001_01001101 : OUT <= 1;  //81 / 77 = 1
    16'b01010001_01001110 : OUT <= 1;  //81 / 78 = 1
    16'b01010001_01001111 : OUT <= 1;  //81 / 79 = 1
    16'b01010001_01010000 : OUT <= 1;  //81 / 80 = 1
    16'b01010001_01010001 : OUT <= 1;  //81 / 81 = 1
    16'b01010001_01010010 : OUT <= 0;  //81 / 82 = 0
    16'b01010001_01010011 : OUT <= 0;  //81 / 83 = 0
    16'b01010001_01010100 : OUT <= 0;  //81 / 84 = 0
    16'b01010001_01010101 : OUT <= 0;  //81 / 85 = 0
    16'b01010001_01010110 : OUT <= 0;  //81 / 86 = 0
    16'b01010001_01010111 : OUT <= 0;  //81 / 87 = 0
    16'b01010001_01011000 : OUT <= 0;  //81 / 88 = 0
    16'b01010001_01011001 : OUT <= 0;  //81 / 89 = 0
    16'b01010001_01011010 : OUT <= 0;  //81 / 90 = 0
    16'b01010001_01011011 : OUT <= 0;  //81 / 91 = 0
    16'b01010001_01011100 : OUT <= 0;  //81 / 92 = 0
    16'b01010001_01011101 : OUT <= 0;  //81 / 93 = 0
    16'b01010001_01011110 : OUT <= 0;  //81 / 94 = 0
    16'b01010001_01011111 : OUT <= 0;  //81 / 95 = 0
    16'b01010001_01100000 : OUT <= 0;  //81 / 96 = 0
    16'b01010001_01100001 : OUT <= 0;  //81 / 97 = 0
    16'b01010001_01100010 : OUT <= 0;  //81 / 98 = 0
    16'b01010001_01100011 : OUT <= 0;  //81 / 99 = 0
    16'b01010001_01100100 : OUT <= 0;  //81 / 100 = 0
    16'b01010001_01100101 : OUT <= 0;  //81 / 101 = 0
    16'b01010001_01100110 : OUT <= 0;  //81 / 102 = 0
    16'b01010001_01100111 : OUT <= 0;  //81 / 103 = 0
    16'b01010001_01101000 : OUT <= 0;  //81 / 104 = 0
    16'b01010001_01101001 : OUT <= 0;  //81 / 105 = 0
    16'b01010001_01101010 : OUT <= 0;  //81 / 106 = 0
    16'b01010001_01101011 : OUT <= 0;  //81 / 107 = 0
    16'b01010001_01101100 : OUT <= 0;  //81 / 108 = 0
    16'b01010001_01101101 : OUT <= 0;  //81 / 109 = 0
    16'b01010001_01101110 : OUT <= 0;  //81 / 110 = 0
    16'b01010001_01101111 : OUT <= 0;  //81 / 111 = 0
    16'b01010001_01110000 : OUT <= 0;  //81 / 112 = 0
    16'b01010001_01110001 : OUT <= 0;  //81 / 113 = 0
    16'b01010001_01110010 : OUT <= 0;  //81 / 114 = 0
    16'b01010001_01110011 : OUT <= 0;  //81 / 115 = 0
    16'b01010001_01110100 : OUT <= 0;  //81 / 116 = 0
    16'b01010001_01110101 : OUT <= 0;  //81 / 117 = 0
    16'b01010001_01110110 : OUT <= 0;  //81 / 118 = 0
    16'b01010001_01110111 : OUT <= 0;  //81 / 119 = 0
    16'b01010001_01111000 : OUT <= 0;  //81 / 120 = 0
    16'b01010001_01111001 : OUT <= 0;  //81 / 121 = 0
    16'b01010001_01111010 : OUT <= 0;  //81 / 122 = 0
    16'b01010001_01111011 : OUT <= 0;  //81 / 123 = 0
    16'b01010001_01111100 : OUT <= 0;  //81 / 124 = 0
    16'b01010001_01111101 : OUT <= 0;  //81 / 125 = 0
    16'b01010001_01111110 : OUT <= 0;  //81 / 126 = 0
    16'b01010001_01111111 : OUT <= 0;  //81 / 127 = 0
    16'b01010001_10000000 : OUT <= 0;  //81 / 128 = 0
    16'b01010001_10000001 : OUT <= 0;  //81 / 129 = 0
    16'b01010001_10000010 : OUT <= 0;  //81 / 130 = 0
    16'b01010001_10000011 : OUT <= 0;  //81 / 131 = 0
    16'b01010001_10000100 : OUT <= 0;  //81 / 132 = 0
    16'b01010001_10000101 : OUT <= 0;  //81 / 133 = 0
    16'b01010001_10000110 : OUT <= 0;  //81 / 134 = 0
    16'b01010001_10000111 : OUT <= 0;  //81 / 135 = 0
    16'b01010001_10001000 : OUT <= 0;  //81 / 136 = 0
    16'b01010001_10001001 : OUT <= 0;  //81 / 137 = 0
    16'b01010001_10001010 : OUT <= 0;  //81 / 138 = 0
    16'b01010001_10001011 : OUT <= 0;  //81 / 139 = 0
    16'b01010001_10001100 : OUT <= 0;  //81 / 140 = 0
    16'b01010001_10001101 : OUT <= 0;  //81 / 141 = 0
    16'b01010001_10001110 : OUT <= 0;  //81 / 142 = 0
    16'b01010001_10001111 : OUT <= 0;  //81 / 143 = 0
    16'b01010001_10010000 : OUT <= 0;  //81 / 144 = 0
    16'b01010001_10010001 : OUT <= 0;  //81 / 145 = 0
    16'b01010001_10010010 : OUT <= 0;  //81 / 146 = 0
    16'b01010001_10010011 : OUT <= 0;  //81 / 147 = 0
    16'b01010001_10010100 : OUT <= 0;  //81 / 148 = 0
    16'b01010001_10010101 : OUT <= 0;  //81 / 149 = 0
    16'b01010001_10010110 : OUT <= 0;  //81 / 150 = 0
    16'b01010001_10010111 : OUT <= 0;  //81 / 151 = 0
    16'b01010001_10011000 : OUT <= 0;  //81 / 152 = 0
    16'b01010001_10011001 : OUT <= 0;  //81 / 153 = 0
    16'b01010001_10011010 : OUT <= 0;  //81 / 154 = 0
    16'b01010001_10011011 : OUT <= 0;  //81 / 155 = 0
    16'b01010001_10011100 : OUT <= 0;  //81 / 156 = 0
    16'b01010001_10011101 : OUT <= 0;  //81 / 157 = 0
    16'b01010001_10011110 : OUT <= 0;  //81 / 158 = 0
    16'b01010001_10011111 : OUT <= 0;  //81 / 159 = 0
    16'b01010001_10100000 : OUT <= 0;  //81 / 160 = 0
    16'b01010001_10100001 : OUT <= 0;  //81 / 161 = 0
    16'b01010001_10100010 : OUT <= 0;  //81 / 162 = 0
    16'b01010001_10100011 : OUT <= 0;  //81 / 163 = 0
    16'b01010001_10100100 : OUT <= 0;  //81 / 164 = 0
    16'b01010001_10100101 : OUT <= 0;  //81 / 165 = 0
    16'b01010001_10100110 : OUT <= 0;  //81 / 166 = 0
    16'b01010001_10100111 : OUT <= 0;  //81 / 167 = 0
    16'b01010001_10101000 : OUT <= 0;  //81 / 168 = 0
    16'b01010001_10101001 : OUT <= 0;  //81 / 169 = 0
    16'b01010001_10101010 : OUT <= 0;  //81 / 170 = 0
    16'b01010001_10101011 : OUT <= 0;  //81 / 171 = 0
    16'b01010001_10101100 : OUT <= 0;  //81 / 172 = 0
    16'b01010001_10101101 : OUT <= 0;  //81 / 173 = 0
    16'b01010001_10101110 : OUT <= 0;  //81 / 174 = 0
    16'b01010001_10101111 : OUT <= 0;  //81 / 175 = 0
    16'b01010001_10110000 : OUT <= 0;  //81 / 176 = 0
    16'b01010001_10110001 : OUT <= 0;  //81 / 177 = 0
    16'b01010001_10110010 : OUT <= 0;  //81 / 178 = 0
    16'b01010001_10110011 : OUT <= 0;  //81 / 179 = 0
    16'b01010001_10110100 : OUT <= 0;  //81 / 180 = 0
    16'b01010001_10110101 : OUT <= 0;  //81 / 181 = 0
    16'b01010001_10110110 : OUT <= 0;  //81 / 182 = 0
    16'b01010001_10110111 : OUT <= 0;  //81 / 183 = 0
    16'b01010001_10111000 : OUT <= 0;  //81 / 184 = 0
    16'b01010001_10111001 : OUT <= 0;  //81 / 185 = 0
    16'b01010001_10111010 : OUT <= 0;  //81 / 186 = 0
    16'b01010001_10111011 : OUT <= 0;  //81 / 187 = 0
    16'b01010001_10111100 : OUT <= 0;  //81 / 188 = 0
    16'b01010001_10111101 : OUT <= 0;  //81 / 189 = 0
    16'b01010001_10111110 : OUT <= 0;  //81 / 190 = 0
    16'b01010001_10111111 : OUT <= 0;  //81 / 191 = 0
    16'b01010001_11000000 : OUT <= 0;  //81 / 192 = 0
    16'b01010001_11000001 : OUT <= 0;  //81 / 193 = 0
    16'b01010001_11000010 : OUT <= 0;  //81 / 194 = 0
    16'b01010001_11000011 : OUT <= 0;  //81 / 195 = 0
    16'b01010001_11000100 : OUT <= 0;  //81 / 196 = 0
    16'b01010001_11000101 : OUT <= 0;  //81 / 197 = 0
    16'b01010001_11000110 : OUT <= 0;  //81 / 198 = 0
    16'b01010001_11000111 : OUT <= 0;  //81 / 199 = 0
    16'b01010001_11001000 : OUT <= 0;  //81 / 200 = 0
    16'b01010001_11001001 : OUT <= 0;  //81 / 201 = 0
    16'b01010001_11001010 : OUT <= 0;  //81 / 202 = 0
    16'b01010001_11001011 : OUT <= 0;  //81 / 203 = 0
    16'b01010001_11001100 : OUT <= 0;  //81 / 204 = 0
    16'b01010001_11001101 : OUT <= 0;  //81 / 205 = 0
    16'b01010001_11001110 : OUT <= 0;  //81 / 206 = 0
    16'b01010001_11001111 : OUT <= 0;  //81 / 207 = 0
    16'b01010001_11010000 : OUT <= 0;  //81 / 208 = 0
    16'b01010001_11010001 : OUT <= 0;  //81 / 209 = 0
    16'b01010001_11010010 : OUT <= 0;  //81 / 210 = 0
    16'b01010001_11010011 : OUT <= 0;  //81 / 211 = 0
    16'b01010001_11010100 : OUT <= 0;  //81 / 212 = 0
    16'b01010001_11010101 : OUT <= 0;  //81 / 213 = 0
    16'b01010001_11010110 : OUT <= 0;  //81 / 214 = 0
    16'b01010001_11010111 : OUT <= 0;  //81 / 215 = 0
    16'b01010001_11011000 : OUT <= 0;  //81 / 216 = 0
    16'b01010001_11011001 : OUT <= 0;  //81 / 217 = 0
    16'b01010001_11011010 : OUT <= 0;  //81 / 218 = 0
    16'b01010001_11011011 : OUT <= 0;  //81 / 219 = 0
    16'b01010001_11011100 : OUT <= 0;  //81 / 220 = 0
    16'b01010001_11011101 : OUT <= 0;  //81 / 221 = 0
    16'b01010001_11011110 : OUT <= 0;  //81 / 222 = 0
    16'b01010001_11011111 : OUT <= 0;  //81 / 223 = 0
    16'b01010001_11100000 : OUT <= 0;  //81 / 224 = 0
    16'b01010001_11100001 : OUT <= 0;  //81 / 225 = 0
    16'b01010001_11100010 : OUT <= 0;  //81 / 226 = 0
    16'b01010001_11100011 : OUT <= 0;  //81 / 227 = 0
    16'b01010001_11100100 : OUT <= 0;  //81 / 228 = 0
    16'b01010001_11100101 : OUT <= 0;  //81 / 229 = 0
    16'b01010001_11100110 : OUT <= 0;  //81 / 230 = 0
    16'b01010001_11100111 : OUT <= 0;  //81 / 231 = 0
    16'b01010001_11101000 : OUT <= 0;  //81 / 232 = 0
    16'b01010001_11101001 : OUT <= 0;  //81 / 233 = 0
    16'b01010001_11101010 : OUT <= 0;  //81 / 234 = 0
    16'b01010001_11101011 : OUT <= 0;  //81 / 235 = 0
    16'b01010001_11101100 : OUT <= 0;  //81 / 236 = 0
    16'b01010001_11101101 : OUT <= 0;  //81 / 237 = 0
    16'b01010001_11101110 : OUT <= 0;  //81 / 238 = 0
    16'b01010001_11101111 : OUT <= 0;  //81 / 239 = 0
    16'b01010001_11110000 : OUT <= 0;  //81 / 240 = 0
    16'b01010001_11110001 : OUT <= 0;  //81 / 241 = 0
    16'b01010001_11110010 : OUT <= 0;  //81 / 242 = 0
    16'b01010001_11110011 : OUT <= 0;  //81 / 243 = 0
    16'b01010001_11110100 : OUT <= 0;  //81 / 244 = 0
    16'b01010001_11110101 : OUT <= 0;  //81 / 245 = 0
    16'b01010001_11110110 : OUT <= 0;  //81 / 246 = 0
    16'b01010001_11110111 : OUT <= 0;  //81 / 247 = 0
    16'b01010001_11111000 : OUT <= 0;  //81 / 248 = 0
    16'b01010001_11111001 : OUT <= 0;  //81 / 249 = 0
    16'b01010001_11111010 : OUT <= 0;  //81 / 250 = 0
    16'b01010001_11111011 : OUT <= 0;  //81 / 251 = 0
    16'b01010001_11111100 : OUT <= 0;  //81 / 252 = 0
    16'b01010001_11111101 : OUT <= 0;  //81 / 253 = 0
    16'b01010001_11111110 : OUT <= 0;  //81 / 254 = 0
    16'b01010001_11111111 : OUT <= 0;  //81 / 255 = 0
    16'b01010010_00000000 : OUT <= 0;  //82 / 0 = 0
    16'b01010010_00000001 : OUT <= 82;  //82 / 1 = 82
    16'b01010010_00000010 : OUT <= 41;  //82 / 2 = 41
    16'b01010010_00000011 : OUT <= 27;  //82 / 3 = 27
    16'b01010010_00000100 : OUT <= 20;  //82 / 4 = 20
    16'b01010010_00000101 : OUT <= 16;  //82 / 5 = 16
    16'b01010010_00000110 : OUT <= 13;  //82 / 6 = 13
    16'b01010010_00000111 : OUT <= 11;  //82 / 7 = 11
    16'b01010010_00001000 : OUT <= 10;  //82 / 8 = 10
    16'b01010010_00001001 : OUT <= 9;  //82 / 9 = 9
    16'b01010010_00001010 : OUT <= 8;  //82 / 10 = 8
    16'b01010010_00001011 : OUT <= 7;  //82 / 11 = 7
    16'b01010010_00001100 : OUT <= 6;  //82 / 12 = 6
    16'b01010010_00001101 : OUT <= 6;  //82 / 13 = 6
    16'b01010010_00001110 : OUT <= 5;  //82 / 14 = 5
    16'b01010010_00001111 : OUT <= 5;  //82 / 15 = 5
    16'b01010010_00010000 : OUT <= 5;  //82 / 16 = 5
    16'b01010010_00010001 : OUT <= 4;  //82 / 17 = 4
    16'b01010010_00010010 : OUT <= 4;  //82 / 18 = 4
    16'b01010010_00010011 : OUT <= 4;  //82 / 19 = 4
    16'b01010010_00010100 : OUT <= 4;  //82 / 20 = 4
    16'b01010010_00010101 : OUT <= 3;  //82 / 21 = 3
    16'b01010010_00010110 : OUT <= 3;  //82 / 22 = 3
    16'b01010010_00010111 : OUT <= 3;  //82 / 23 = 3
    16'b01010010_00011000 : OUT <= 3;  //82 / 24 = 3
    16'b01010010_00011001 : OUT <= 3;  //82 / 25 = 3
    16'b01010010_00011010 : OUT <= 3;  //82 / 26 = 3
    16'b01010010_00011011 : OUT <= 3;  //82 / 27 = 3
    16'b01010010_00011100 : OUT <= 2;  //82 / 28 = 2
    16'b01010010_00011101 : OUT <= 2;  //82 / 29 = 2
    16'b01010010_00011110 : OUT <= 2;  //82 / 30 = 2
    16'b01010010_00011111 : OUT <= 2;  //82 / 31 = 2
    16'b01010010_00100000 : OUT <= 2;  //82 / 32 = 2
    16'b01010010_00100001 : OUT <= 2;  //82 / 33 = 2
    16'b01010010_00100010 : OUT <= 2;  //82 / 34 = 2
    16'b01010010_00100011 : OUT <= 2;  //82 / 35 = 2
    16'b01010010_00100100 : OUT <= 2;  //82 / 36 = 2
    16'b01010010_00100101 : OUT <= 2;  //82 / 37 = 2
    16'b01010010_00100110 : OUT <= 2;  //82 / 38 = 2
    16'b01010010_00100111 : OUT <= 2;  //82 / 39 = 2
    16'b01010010_00101000 : OUT <= 2;  //82 / 40 = 2
    16'b01010010_00101001 : OUT <= 2;  //82 / 41 = 2
    16'b01010010_00101010 : OUT <= 1;  //82 / 42 = 1
    16'b01010010_00101011 : OUT <= 1;  //82 / 43 = 1
    16'b01010010_00101100 : OUT <= 1;  //82 / 44 = 1
    16'b01010010_00101101 : OUT <= 1;  //82 / 45 = 1
    16'b01010010_00101110 : OUT <= 1;  //82 / 46 = 1
    16'b01010010_00101111 : OUT <= 1;  //82 / 47 = 1
    16'b01010010_00110000 : OUT <= 1;  //82 / 48 = 1
    16'b01010010_00110001 : OUT <= 1;  //82 / 49 = 1
    16'b01010010_00110010 : OUT <= 1;  //82 / 50 = 1
    16'b01010010_00110011 : OUT <= 1;  //82 / 51 = 1
    16'b01010010_00110100 : OUT <= 1;  //82 / 52 = 1
    16'b01010010_00110101 : OUT <= 1;  //82 / 53 = 1
    16'b01010010_00110110 : OUT <= 1;  //82 / 54 = 1
    16'b01010010_00110111 : OUT <= 1;  //82 / 55 = 1
    16'b01010010_00111000 : OUT <= 1;  //82 / 56 = 1
    16'b01010010_00111001 : OUT <= 1;  //82 / 57 = 1
    16'b01010010_00111010 : OUT <= 1;  //82 / 58 = 1
    16'b01010010_00111011 : OUT <= 1;  //82 / 59 = 1
    16'b01010010_00111100 : OUT <= 1;  //82 / 60 = 1
    16'b01010010_00111101 : OUT <= 1;  //82 / 61 = 1
    16'b01010010_00111110 : OUT <= 1;  //82 / 62 = 1
    16'b01010010_00111111 : OUT <= 1;  //82 / 63 = 1
    16'b01010010_01000000 : OUT <= 1;  //82 / 64 = 1
    16'b01010010_01000001 : OUT <= 1;  //82 / 65 = 1
    16'b01010010_01000010 : OUT <= 1;  //82 / 66 = 1
    16'b01010010_01000011 : OUT <= 1;  //82 / 67 = 1
    16'b01010010_01000100 : OUT <= 1;  //82 / 68 = 1
    16'b01010010_01000101 : OUT <= 1;  //82 / 69 = 1
    16'b01010010_01000110 : OUT <= 1;  //82 / 70 = 1
    16'b01010010_01000111 : OUT <= 1;  //82 / 71 = 1
    16'b01010010_01001000 : OUT <= 1;  //82 / 72 = 1
    16'b01010010_01001001 : OUT <= 1;  //82 / 73 = 1
    16'b01010010_01001010 : OUT <= 1;  //82 / 74 = 1
    16'b01010010_01001011 : OUT <= 1;  //82 / 75 = 1
    16'b01010010_01001100 : OUT <= 1;  //82 / 76 = 1
    16'b01010010_01001101 : OUT <= 1;  //82 / 77 = 1
    16'b01010010_01001110 : OUT <= 1;  //82 / 78 = 1
    16'b01010010_01001111 : OUT <= 1;  //82 / 79 = 1
    16'b01010010_01010000 : OUT <= 1;  //82 / 80 = 1
    16'b01010010_01010001 : OUT <= 1;  //82 / 81 = 1
    16'b01010010_01010010 : OUT <= 1;  //82 / 82 = 1
    16'b01010010_01010011 : OUT <= 0;  //82 / 83 = 0
    16'b01010010_01010100 : OUT <= 0;  //82 / 84 = 0
    16'b01010010_01010101 : OUT <= 0;  //82 / 85 = 0
    16'b01010010_01010110 : OUT <= 0;  //82 / 86 = 0
    16'b01010010_01010111 : OUT <= 0;  //82 / 87 = 0
    16'b01010010_01011000 : OUT <= 0;  //82 / 88 = 0
    16'b01010010_01011001 : OUT <= 0;  //82 / 89 = 0
    16'b01010010_01011010 : OUT <= 0;  //82 / 90 = 0
    16'b01010010_01011011 : OUT <= 0;  //82 / 91 = 0
    16'b01010010_01011100 : OUT <= 0;  //82 / 92 = 0
    16'b01010010_01011101 : OUT <= 0;  //82 / 93 = 0
    16'b01010010_01011110 : OUT <= 0;  //82 / 94 = 0
    16'b01010010_01011111 : OUT <= 0;  //82 / 95 = 0
    16'b01010010_01100000 : OUT <= 0;  //82 / 96 = 0
    16'b01010010_01100001 : OUT <= 0;  //82 / 97 = 0
    16'b01010010_01100010 : OUT <= 0;  //82 / 98 = 0
    16'b01010010_01100011 : OUT <= 0;  //82 / 99 = 0
    16'b01010010_01100100 : OUT <= 0;  //82 / 100 = 0
    16'b01010010_01100101 : OUT <= 0;  //82 / 101 = 0
    16'b01010010_01100110 : OUT <= 0;  //82 / 102 = 0
    16'b01010010_01100111 : OUT <= 0;  //82 / 103 = 0
    16'b01010010_01101000 : OUT <= 0;  //82 / 104 = 0
    16'b01010010_01101001 : OUT <= 0;  //82 / 105 = 0
    16'b01010010_01101010 : OUT <= 0;  //82 / 106 = 0
    16'b01010010_01101011 : OUT <= 0;  //82 / 107 = 0
    16'b01010010_01101100 : OUT <= 0;  //82 / 108 = 0
    16'b01010010_01101101 : OUT <= 0;  //82 / 109 = 0
    16'b01010010_01101110 : OUT <= 0;  //82 / 110 = 0
    16'b01010010_01101111 : OUT <= 0;  //82 / 111 = 0
    16'b01010010_01110000 : OUT <= 0;  //82 / 112 = 0
    16'b01010010_01110001 : OUT <= 0;  //82 / 113 = 0
    16'b01010010_01110010 : OUT <= 0;  //82 / 114 = 0
    16'b01010010_01110011 : OUT <= 0;  //82 / 115 = 0
    16'b01010010_01110100 : OUT <= 0;  //82 / 116 = 0
    16'b01010010_01110101 : OUT <= 0;  //82 / 117 = 0
    16'b01010010_01110110 : OUT <= 0;  //82 / 118 = 0
    16'b01010010_01110111 : OUT <= 0;  //82 / 119 = 0
    16'b01010010_01111000 : OUT <= 0;  //82 / 120 = 0
    16'b01010010_01111001 : OUT <= 0;  //82 / 121 = 0
    16'b01010010_01111010 : OUT <= 0;  //82 / 122 = 0
    16'b01010010_01111011 : OUT <= 0;  //82 / 123 = 0
    16'b01010010_01111100 : OUT <= 0;  //82 / 124 = 0
    16'b01010010_01111101 : OUT <= 0;  //82 / 125 = 0
    16'b01010010_01111110 : OUT <= 0;  //82 / 126 = 0
    16'b01010010_01111111 : OUT <= 0;  //82 / 127 = 0
    16'b01010010_10000000 : OUT <= 0;  //82 / 128 = 0
    16'b01010010_10000001 : OUT <= 0;  //82 / 129 = 0
    16'b01010010_10000010 : OUT <= 0;  //82 / 130 = 0
    16'b01010010_10000011 : OUT <= 0;  //82 / 131 = 0
    16'b01010010_10000100 : OUT <= 0;  //82 / 132 = 0
    16'b01010010_10000101 : OUT <= 0;  //82 / 133 = 0
    16'b01010010_10000110 : OUT <= 0;  //82 / 134 = 0
    16'b01010010_10000111 : OUT <= 0;  //82 / 135 = 0
    16'b01010010_10001000 : OUT <= 0;  //82 / 136 = 0
    16'b01010010_10001001 : OUT <= 0;  //82 / 137 = 0
    16'b01010010_10001010 : OUT <= 0;  //82 / 138 = 0
    16'b01010010_10001011 : OUT <= 0;  //82 / 139 = 0
    16'b01010010_10001100 : OUT <= 0;  //82 / 140 = 0
    16'b01010010_10001101 : OUT <= 0;  //82 / 141 = 0
    16'b01010010_10001110 : OUT <= 0;  //82 / 142 = 0
    16'b01010010_10001111 : OUT <= 0;  //82 / 143 = 0
    16'b01010010_10010000 : OUT <= 0;  //82 / 144 = 0
    16'b01010010_10010001 : OUT <= 0;  //82 / 145 = 0
    16'b01010010_10010010 : OUT <= 0;  //82 / 146 = 0
    16'b01010010_10010011 : OUT <= 0;  //82 / 147 = 0
    16'b01010010_10010100 : OUT <= 0;  //82 / 148 = 0
    16'b01010010_10010101 : OUT <= 0;  //82 / 149 = 0
    16'b01010010_10010110 : OUT <= 0;  //82 / 150 = 0
    16'b01010010_10010111 : OUT <= 0;  //82 / 151 = 0
    16'b01010010_10011000 : OUT <= 0;  //82 / 152 = 0
    16'b01010010_10011001 : OUT <= 0;  //82 / 153 = 0
    16'b01010010_10011010 : OUT <= 0;  //82 / 154 = 0
    16'b01010010_10011011 : OUT <= 0;  //82 / 155 = 0
    16'b01010010_10011100 : OUT <= 0;  //82 / 156 = 0
    16'b01010010_10011101 : OUT <= 0;  //82 / 157 = 0
    16'b01010010_10011110 : OUT <= 0;  //82 / 158 = 0
    16'b01010010_10011111 : OUT <= 0;  //82 / 159 = 0
    16'b01010010_10100000 : OUT <= 0;  //82 / 160 = 0
    16'b01010010_10100001 : OUT <= 0;  //82 / 161 = 0
    16'b01010010_10100010 : OUT <= 0;  //82 / 162 = 0
    16'b01010010_10100011 : OUT <= 0;  //82 / 163 = 0
    16'b01010010_10100100 : OUT <= 0;  //82 / 164 = 0
    16'b01010010_10100101 : OUT <= 0;  //82 / 165 = 0
    16'b01010010_10100110 : OUT <= 0;  //82 / 166 = 0
    16'b01010010_10100111 : OUT <= 0;  //82 / 167 = 0
    16'b01010010_10101000 : OUT <= 0;  //82 / 168 = 0
    16'b01010010_10101001 : OUT <= 0;  //82 / 169 = 0
    16'b01010010_10101010 : OUT <= 0;  //82 / 170 = 0
    16'b01010010_10101011 : OUT <= 0;  //82 / 171 = 0
    16'b01010010_10101100 : OUT <= 0;  //82 / 172 = 0
    16'b01010010_10101101 : OUT <= 0;  //82 / 173 = 0
    16'b01010010_10101110 : OUT <= 0;  //82 / 174 = 0
    16'b01010010_10101111 : OUT <= 0;  //82 / 175 = 0
    16'b01010010_10110000 : OUT <= 0;  //82 / 176 = 0
    16'b01010010_10110001 : OUT <= 0;  //82 / 177 = 0
    16'b01010010_10110010 : OUT <= 0;  //82 / 178 = 0
    16'b01010010_10110011 : OUT <= 0;  //82 / 179 = 0
    16'b01010010_10110100 : OUT <= 0;  //82 / 180 = 0
    16'b01010010_10110101 : OUT <= 0;  //82 / 181 = 0
    16'b01010010_10110110 : OUT <= 0;  //82 / 182 = 0
    16'b01010010_10110111 : OUT <= 0;  //82 / 183 = 0
    16'b01010010_10111000 : OUT <= 0;  //82 / 184 = 0
    16'b01010010_10111001 : OUT <= 0;  //82 / 185 = 0
    16'b01010010_10111010 : OUT <= 0;  //82 / 186 = 0
    16'b01010010_10111011 : OUT <= 0;  //82 / 187 = 0
    16'b01010010_10111100 : OUT <= 0;  //82 / 188 = 0
    16'b01010010_10111101 : OUT <= 0;  //82 / 189 = 0
    16'b01010010_10111110 : OUT <= 0;  //82 / 190 = 0
    16'b01010010_10111111 : OUT <= 0;  //82 / 191 = 0
    16'b01010010_11000000 : OUT <= 0;  //82 / 192 = 0
    16'b01010010_11000001 : OUT <= 0;  //82 / 193 = 0
    16'b01010010_11000010 : OUT <= 0;  //82 / 194 = 0
    16'b01010010_11000011 : OUT <= 0;  //82 / 195 = 0
    16'b01010010_11000100 : OUT <= 0;  //82 / 196 = 0
    16'b01010010_11000101 : OUT <= 0;  //82 / 197 = 0
    16'b01010010_11000110 : OUT <= 0;  //82 / 198 = 0
    16'b01010010_11000111 : OUT <= 0;  //82 / 199 = 0
    16'b01010010_11001000 : OUT <= 0;  //82 / 200 = 0
    16'b01010010_11001001 : OUT <= 0;  //82 / 201 = 0
    16'b01010010_11001010 : OUT <= 0;  //82 / 202 = 0
    16'b01010010_11001011 : OUT <= 0;  //82 / 203 = 0
    16'b01010010_11001100 : OUT <= 0;  //82 / 204 = 0
    16'b01010010_11001101 : OUT <= 0;  //82 / 205 = 0
    16'b01010010_11001110 : OUT <= 0;  //82 / 206 = 0
    16'b01010010_11001111 : OUT <= 0;  //82 / 207 = 0
    16'b01010010_11010000 : OUT <= 0;  //82 / 208 = 0
    16'b01010010_11010001 : OUT <= 0;  //82 / 209 = 0
    16'b01010010_11010010 : OUT <= 0;  //82 / 210 = 0
    16'b01010010_11010011 : OUT <= 0;  //82 / 211 = 0
    16'b01010010_11010100 : OUT <= 0;  //82 / 212 = 0
    16'b01010010_11010101 : OUT <= 0;  //82 / 213 = 0
    16'b01010010_11010110 : OUT <= 0;  //82 / 214 = 0
    16'b01010010_11010111 : OUT <= 0;  //82 / 215 = 0
    16'b01010010_11011000 : OUT <= 0;  //82 / 216 = 0
    16'b01010010_11011001 : OUT <= 0;  //82 / 217 = 0
    16'b01010010_11011010 : OUT <= 0;  //82 / 218 = 0
    16'b01010010_11011011 : OUT <= 0;  //82 / 219 = 0
    16'b01010010_11011100 : OUT <= 0;  //82 / 220 = 0
    16'b01010010_11011101 : OUT <= 0;  //82 / 221 = 0
    16'b01010010_11011110 : OUT <= 0;  //82 / 222 = 0
    16'b01010010_11011111 : OUT <= 0;  //82 / 223 = 0
    16'b01010010_11100000 : OUT <= 0;  //82 / 224 = 0
    16'b01010010_11100001 : OUT <= 0;  //82 / 225 = 0
    16'b01010010_11100010 : OUT <= 0;  //82 / 226 = 0
    16'b01010010_11100011 : OUT <= 0;  //82 / 227 = 0
    16'b01010010_11100100 : OUT <= 0;  //82 / 228 = 0
    16'b01010010_11100101 : OUT <= 0;  //82 / 229 = 0
    16'b01010010_11100110 : OUT <= 0;  //82 / 230 = 0
    16'b01010010_11100111 : OUT <= 0;  //82 / 231 = 0
    16'b01010010_11101000 : OUT <= 0;  //82 / 232 = 0
    16'b01010010_11101001 : OUT <= 0;  //82 / 233 = 0
    16'b01010010_11101010 : OUT <= 0;  //82 / 234 = 0
    16'b01010010_11101011 : OUT <= 0;  //82 / 235 = 0
    16'b01010010_11101100 : OUT <= 0;  //82 / 236 = 0
    16'b01010010_11101101 : OUT <= 0;  //82 / 237 = 0
    16'b01010010_11101110 : OUT <= 0;  //82 / 238 = 0
    16'b01010010_11101111 : OUT <= 0;  //82 / 239 = 0
    16'b01010010_11110000 : OUT <= 0;  //82 / 240 = 0
    16'b01010010_11110001 : OUT <= 0;  //82 / 241 = 0
    16'b01010010_11110010 : OUT <= 0;  //82 / 242 = 0
    16'b01010010_11110011 : OUT <= 0;  //82 / 243 = 0
    16'b01010010_11110100 : OUT <= 0;  //82 / 244 = 0
    16'b01010010_11110101 : OUT <= 0;  //82 / 245 = 0
    16'b01010010_11110110 : OUT <= 0;  //82 / 246 = 0
    16'b01010010_11110111 : OUT <= 0;  //82 / 247 = 0
    16'b01010010_11111000 : OUT <= 0;  //82 / 248 = 0
    16'b01010010_11111001 : OUT <= 0;  //82 / 249 = 0
    16'b01010010_11111010 : OUT <= 0;  //82 / 250 = 0
    16'b01010010_11111011 : OUT <= 0;  //82 / 251 = 0
    16'b01010010_11111100 : OUT <= 0;  //82 / 252 = 0
    16'b01010010_11111101 : OUT <= 0;  //82 / 253 = 0
    16'b01010010_11111110 : OUT <= 0;  //82 / 254 = 0
    16'b01010010_11111111 : OUT <= 0;  //82 / 255 = 0
    16'b01010011_00000000 : OUT <= 0;  //83 / 0 = 0
    16'b01010011_00000001 : OUT <= 83;  //83 / 1 = 83
    16'b01010011_00000010 : OUT <= 41;  //83 / 2 = 41
    16'b01010011_00000011 : OUT <= 27;  //83 / 3 = 27
    16'b01010011_00000100 : OUT <= 20;  //83 / 4 = 20
    16'b01010011_00000101 : OUT <= 16;  //83 / 5 = 16
    16'b01010011_00000110 : OUT <= 13;  //83 / 6 = 13
    16'b01010011_00000111 : OUT <= 11;  //83 / 7 = 11
    16'b01010011_00001000 : OUT <= 10;  //83 / 8 = 10
    16'b01010011_00001001 : OUT <= 9;  //83 / 9 = 9
    16'b01010011_00001010 : OUT <= 8;  //83 / 10 = 8
    16'b01010011_00001011 : OUT <= 7;  //83 / 11 = 7
    16'b01010011_00001100 : OUT <= 6;  //83 / 12 = 6
    16'b01010011_00001101 : OUT <= 6;  //83 / 13 = 6
    16'b01010011_00001110 : OUT <= 5;  //83 / 14 = 5
    16'b01010011_00001111 : OUT <= 5;  //83 / 15 = 5
    16'b01010011_00010000 : OUT <= 5;  //83 / 16 = 5
    16'b01010011_00010001 : OUT <= 4;  //83 / 17 = 4
    16'b01010011_00010010 : OUT <= 4;  //83 / 18 = 4
    16'b01010011_00010011 : OUT <= 4;  //83 / 19 = 4
    16'b01010011_00010100 : OUT <= 4;  //83 / 20 = 4
    16'b01010011_00010101 : OUT <= 3;  //83 / 21 = 3
    16'b01010011_00010110 : OUT <= 3;  //83 / 22 = 3
    16'b01010011_00010111 : OUT <= 3;  //83 / 23 = 3
    16'b01010011_00011000 : OUT <= 3;  //83 / 24 = 3
    16'b01010011_00011001 : OUT <= 3;  //83 / 25 = 3
    16'b01010011_00011010 : OUT <= 3;  //83 / 26 = 3
    16'b01010011_00011011 : OUT <= 3;  //83 / 27 = 3
    16'b01010011_00011100 : OUT <= 2;  //83 / 28 = 2
    16'b01010011_00011101 : OUT <= 2;  //83 / 29 = 2
    16'b01010011_00011110 : OUT <= 2;  //83 / 30 = 2
    16'b01010011_00011111 : OUT <= 2;  //83 / 31 = 2
    16'b01010011_00100000 : OUT <= 2;  //83 / 32 = 2
    16'b01010011_00100001 : OUT <= 2;  //83 / 33 = 2
    16'b01010011_00100010 : OUT <= 2;  //83 / 34 = 2
    16'b01010011_00100011 : OUT <= 2;  //83 / 35 = 2
    16'b01010011_00100100 : OUT <= 2;  //83 / 36 = 2
    16'b01010011_00100101 : OUT <= 2;  //83 / 37 = 2
    16'b01010011_00100110 : OUT <= 2;  //83 / 38 = 2
    16'b01010011_00100111 : OUT <= 2;  //83 / 39 = 2
    16'b01010011_00101000 : OUT <= 2;  //83 / 40 = 2
    16'b01010011_00101001 : OUT <= 2;  //83 / 41 = 2
    16'b01010011_00101010 : OUT <= 1;  //83 / 42 = 1
    16'b01010011_00101011 : OUT <= 1;  //83 / 43 = 1
    16'b01010011_00101100 : OUT <= 1;  //83 / 44 = 1
    16'b01010011_00101101 : OUT <= 1;  //83 / 45 = 1
    16'b01010011_00101110 : OUT <= 1;  //83 / 46 = 1
    16'b01010011_00101111 : OUT <= 1;  //83 / 47 = 1
    16'b01010011_00110000 : OUT <= 1;  //83 / 48 = 1
    16'b01010011_00110001 : OUT <= 1;  //83 / 49 = 1
    16'b01010011_00110010 : OUT <= 1;  //83 / 50 = 1
    16'b01010011_00110011 : OUT <= 1;  //83 / 51 = 1
    16'b01010011_00110100 : OUT <= 1;  //83 / 52 = 1
    16'b01010011_00110101 : OUT <= 1;  //83 / 53 = 1
    16'b01010011_00110110 : OUT <= 1;  //83 / 54 = 1
    16'b01010011_00110111 : OUT <= 1;  //83 / 55 = 1
    16'b01010011_00111000 : OUT <= 1;  //83 / 56 = 1
    16'b01010011_00111001 : OUT <= 1;  //83 / 57 = 1
    16'b01010011_00111010 : OUT <= 1;  //83 / 58 = 1
    16'b01010011_00111011 : OUT <= 1;  //83 / 59 = 1
    16'b01010011_00111100 : OUT <= 1;  //83 / 60 = 1
    16'b01010011_00111101 : OUT <= 1;  //83 / 61 = 1
    16'b01010011_00111110 : OUT <= 1;  //83 / 62 = 1
    16'b01010011_00111111 : OUT <= 1;  //83 / 63 = 1
    16'b01010011_01000000 : OUT <= 1;  //83 / 64 = 1
    16'b01010011_01000001 : OUT <= 1;  //83 / 65 = 1
    16'b01010011_01000010 : OUT <= 1;  //83 / 66 = 1
    16'b01010011_01000011 : OUT <= 1;  //83 / 67 = 1
    16'b01010011_01000100 : OUT <= 1;  //83 / 68 = 1
    16'b01010011_01000101 : OUT <= 1;  //83 / 69 = 1
    16'b01010011_01000110 : OUT <= 1;  //83 / 70 = 1
    16'b01010011_01000111 : OUT <= 1;  //83 / 71 = 1
    16'b01010011_01001000 : OUT <= 1;  //83 / 72 = 1
    16'b01010011_01001001 : OUT <= 1;  //83 / 73 = 1
    16'b01010011_01001010 : OUT <= 1;  //83 / 74 = 1
    16'b01010011_01001011 : OUT <= 1;  //83 / 75 = 1
    16'b01010011_01001100 : OUT <= 1;  //83 / 76 = 1
    16'b01010011_01001101 : OUT <= 1;  //83 / 77 = 1
    16'b01010011_01001110 : OUT <= 1;  //83 / 78 = 1
    16'b01010011_01001111 : OUT <= 1;  //83 / 79 = 1
    16'b01010011_01010000 : OUT <= 1;  //83 / 80 = 1
    16'b01010011_01010001 : OUT <= 1;  //83 / 81 = 1
    16'b01010011_01010010 : OUT <= 1;  //83 / 82 = 1
    16'b01010011_01010011 : OUT <= 1;  //83 / 83 = 1
    16'b01010011_01010100 : OUT <= 0;  //83 / 84 = 0
    16'b01010011_01010101 : OUT <= 0;  //83 / 85 = 0
    16'b01010011_01010110 : OUT <= 0;  //83 / 86 = 0
    16'b01010011_01010111 : OUT <= 0;  //83 / 87 = 0
    16'b01010011_01011000 : OUT <= 0;  //83 / 88 = 0
    16'b01010011_01011001 : OUT <= 0;  //83 / 89 = 0
    16'b01010011_01011010 : OUT <= 0;  //83 / 90 = 0
    16'b01010011_01011011 : OUT <= 0;  //83 / 91 = 0
    16'b01010011_01011100 : OUT <= 0;  //83 / 92 = 0
    16'b01010011_01011101 : OUT <= 0;  //83 / 93 = 0
    16'b01010011_01011110 : OUT <= 0;  //83 / 94 = 0
    16'b01010011_01011111 : OUT <= 0;  //83 / 95 = 0
    16'b01010011_01100000 : OUT <= 0;  //83 / 96 = 0
    16'b01010011_01100001 : OUT <= 0;  //83 / 97 = 0
    16'b01010011_01100010 : OUT <= 0;  //83 / 98 = 0
    16'b01010011_01100011 : OUT <= 0;  //83 / 99 = 0
    16'b01010011_01100100 : OUT <= 0;  //83 / 100 = 0
    16'b01010011_01100101 : OUT <= 0;  //83 / 101 = 0
    16'b01010011_01100110 : OUT <= 0;  //83 / 102 = 0
    16'b01010011_01100111 : OUT <= 0;  //83 / 103 = 0
    16'b01010011_01101000 : OUT <= 0;  //83 / 104 = 0
    16'b01010011_01101001 : OUT <= 0;  //83 / 105 = 0
    16'b01010011_01101010 : OUT <= 0;  //83 / 106 = 0
    16'b01010011_01101011 : OUT <= 0;  //83 / 107 = 0
    16'b01010011_01101100 : OUT <= 0;  //83 / 108 = 0
    16'b01010011_01101101 : OUT <= 0;  //83 / 109 = 0
    16'b01010011_01101110 : OUT <= 0;  //83 / 110 = 0
    16'b01010011_01101111 : OUT <= 0;  //83 / 111 = 0
    16'b01010011_01110000 : OUT <= 0;  //83 / 112 = 0
    16'b01010011_01110001 : OUT <= 0;  //83 / 113 = 0
    16'b01010011_01110010 : OUT <= 0;  //83 / 114 = 0
    16'b01010011_01110011 : OUT <= 0;  //83 / 115 = 0
    16'b01010011_01110100 : OUT <= 0;  //83 / 116 = 0
    16'b01010011_01110101 : OUT <= 0;  //83 / 117 = 0
    16'b01010011_01110110 : OUT <= 0;  //83 / 118 = 0
    16'b01010011_01110111 : OUT <= 0;  //83 / 119 = 0
    16'b01010011_01111000 : OUT <= 0;  //83 / 120 = 0
    16'b01010011_01111001 : OUT <= 0;  //83 / 121 = 0
    16'b01010011_01111010 : OUT <= 0;  //83 / 122 = 0
    16'b01010011_01111011 : OUT <= 0;  //83 / 123 = 0
    16'b01010011_01111100 : OUT <= 0;  //83 / 124 = 0
    16'b01010011_01111101 : OUT <= 0;  //83 / 125 = 0
    16'b01010011_01111110 : OUT <= 0;  //83 / 126 = 0
    16'b01010011_01111111 : OUT <= 0;  //83 / 127 = 0
    16'b01010011_10000000 : OUT <= 0;  //83 / 128 = 0
    16'b01010011_10000001 : OUT <= 0;  //83 / 129 = 0
    16'b01010011_10000010 : OUT <= 0;  //83 / 130 = 0
    16'b01010011_10000011 : OUT <= 0;  //83 / 131 = 0
    16'b01010011_10000100 : OUT <= 0;  //83 / 132 = 0
    16'b01010011_10000101 : OUT <= 0;  //83 / 133 = 0
    16'b01010011_10000110 : OUT <= 0;  //83 / 134 = 0
    16'b01010011_10000111 : OUT <= 0;  //83 / 135 = 0
    16'b01010011_10001000 : OUT <= 0;  //83 / 136 = 0
    16'b01010011_10001001 : OUT <= 0;  //83 / 137 = 0
    16'b01010011_10001010 : OUT <= 0;  //83 / 138 = 0
    16'b01010011_10001011 : OUT <= 0;  //83 / 139 = 0
    16'b01010011_10001100 : OUT <= 0;  //83 / 140 = 0
    16'b01010011_10001101 : OUT <= 0;  //83 / 141 = 0
    16'b01010011_10001110 : OUT <= 0;  //83 / 142 = 0
    16'b01010011_10001111 : OUT <= 0;  //83 / 143 = 0
    16'b01010011_10010000 : OUT <= 0;  //83 / 144 = 0
    16'b01010011_10010001 : OUT <= 0;  //83 / 145 = 0
    16'b01010011_10010010 : OUT <= 0;  //83 / 146 = 0
    16'b01010011_10010011 : OUT <= 0;  //83 / 147 = 0
    16'b01010011_10010100 : OUT <= 0;  //83 / 148 = 0
    16'b01010011_10010101 : OUT <= 0;  //83 / 149 = 0
    16'b01010011_10010110 : OUT <= 0;  //83 / 150 = 0
    16'b01010011_10010111 : OUT <= 0;  //83 / 151 = 0
    16'b01010011_10011000 : OUT <= 0;  //83 / 152 = 0
    16'b01010011_10011001 : OUT <= 0;  //83 / 153 = 0
    16'b01010011_10011010 : OUT <= 0;  //83 / 154 = 0
    16'b01010011_10011011 : OUT <= 0;  //83 / 155 = 0
    16'b01010011_10011100 : OUT <= 0;  //83 / 156 = 0
    16'b01010011_10011101 : OUT <= 0;  //83 / 157 = 0
    16'b01010011_10011110 : OUT <= 0;  //83 / 158 = 0
    16'b01010011_10011111 : OUT <= 0;  //83 / 159 = 0
    16'b01010011_10100000 : OUT <= 0;  //83 / 160 = 0
    16'b01010011_10100001 : OUT <= 0;  //83 / 161 = 0
    16'b01010011_10100010 : OUT <= 0;  //83 / 162 = 0
    16'b01010011_10100011 : OUT <= 0;  //83 / 163 = 0
    16'b01010011_10100100 : OUT <= 0;  //83 / 164 = 0
    16'b01010011_10100101 : OUT <= 0;  //83 / 165 = 0
    16'b01010011_10100110 : OUT <= 0;  //83 / 166 = 0
    16'b01010011_10100111 : OUT <= 0;  //83 / 167 = 0
    16'b01010011_10101000 : OUT <= 0;  //83 / 168 = 0
    16'b01010011_10101001 : OUT <= 0;  //83 / 169 = 0
    16'b01010011_10101010 : OUT <= 0;  //83 / 170 = 0
    16'b01010011_10101011 : OUT <= 0;  //83 / 171 = 0
    16'b01010011_10101100 : OUT <= 0;  //83 / 172 = 0
    16'b01010011_10101101 : OUT <= 0;  //83 / 173 = 0
    16'b01010011_10101110 : OUT <= 0;  //83 / 174 = 0
    16'b01010011_10101111 : OUT <= 0;  //83 / 175 = 0
    16'b01010011_10110000 : OUT <= 0;  //83 / 176 = 0
    16'b01010011_10110001 : OUT <= 0;  //83 / 177 = 0
    16'b01010011_10110010 : OUT <= 0;  //83 / 178 = 0
    16'b01010011_10110011 : OUT <= 0;  //83 / 179 = 0
    16'b01010011_10110100 : OUT <= 0;  //83 / 180 = 0
    16'b01010011_10110101 : OUT <= 0;  //83 / 181 = 0
    16'b01010011_10110110 : OUT <= 0;  //83 / 182 = 0
    16'b01010011_10110111 : OUT <= 0;  //83 / 183 = 0
    16'b01010011_10111000 : OUT <= 0;  //83 / 184 = 0
    16'b01010011_10111001 : OUT <= 0;  //83 / 185 = 0
    16'b01010011_10111010 : OUT <= 0;  //83 / 186 = 0
    16'b01010011_10111011 : OUT <= 0;  //83 / 187 = 0
    16'b01010011_10111100 : OUT <= 0;  //83 / 188 = 0
    16'b01010011_10111101 : OUT <= 0;  //83 / 189 = 0
    16'b01010011_10111110 : OUT <= 0;  //83 / 190 = 0
    16'b01010011_10111111 : OUT <= 0;  //83 / 191 = 0
    16'b01010011_11000000 : OUT <= 0;  //83 / 192 = 0
    16'b01010011_11000001 : OUT <= 0;  //83 / 193 = 0
    16'b01010011_11000010 : OUT <= 0;  //83 / 194 = 0
    16'b01010011_11000011 : OUT <= 0;  //83 / 195 = 0
    16'b01010011_11000100 : OUT <= 0;  //83 / 196 = 0
    16'b01010011_11000101 : OUT <= 0;  //83 / 197 = 0
    16'b01010011_11000110 : OUT <= 0;  //83 / 198 = 0
    16'b01010011_11000111 : OUT <= 0;  //83 / 199 = 0
    16'b01010011_11001000 : OUT <= 0;  //83 / 200 = 0
    16'b01010011_11001001 : OUT <= 0;  //83 / 201 = 0
    16'b01010011_11001010 : OUT <= 0;  //83 / 202 = 0
    16'b01010011_11001011 : OUT <= 0;  //83 / 203 = 0
    16'b01010011_11001100 : OUT <= 0;  //83 / 204 = 0
    16'b01010011_11001101 : OUT <= 0;  //83 / 205 = 0
    16'b01010011_11001110 : OUT <= 0;  //83 / 206 = 0
    16'b01010011_11001111 : OUT <= 0;  //83 / 207 = 0
    16'b01010011_11010000 : OUT <= 0;  //83 / 208 = 0
    16'b01010011_11010001 : OUT <= 0;  //83 / 209 = 0
    16'b01010011_11010010 : OUT <= 0;  //83 / 210 = 0
    16'b01010011_11010011 : OUT <= 0;  //83 / 211 = 0
    16'b01010011_11010100 : OUT <= 0;  //83 / 212 = 0
    16'b01010011_11010101 : OUT <= 0;  //83 / 213 = 0
    16'b01010011_11010110 : OUT <= 0;  //83 / 214 = 0
    16'b01010011_11010111 : OUT <= 0;  //83 / 215 = 0
    16'b01010011_11011000 : OUT <= 0;  //83 / 216 = 0
    16'b01010011_11011001 : OUT <= 0;  //83 / 217 = 0
    16'b01010011_11011010 : OUT <= 0;  //83 / 218 = 0
    16'b01010011_11011011 : OUT <= 0;  //83 / 219 = 0
    16'b01010011_11011100 : OUT <= 0;  //83 / 220 = 0
    16'b01010011_11011101 : OUT <= 0;  //83 / 221 = 0
    16'b01010011_11011110 : OUT <= 0;  //83 / 222 = 0
    16'b01010011_11011111 : OUT <= 0;  //83 / 223 = 0
    16'b01010011_11100000 : OUT <= 0;  //83 / 224 = 0
    16'b01010011_11100001 : OUT <= 0;  //83 / 225 = 0
    16'b01010011_11100010 : OUT <= 0;  //83 / 226 = 0
    16'b01010011_11100011 : OUT <= 0;  //83 / 227 = 0
    16'b01010011_11100100 : OUT <= 0;  //83 / 228 = 0
    16'b01010011_11100101 : OUT <= 0;  //83 / 229 = 0
    16'b01010011_11100110 : OUT <= 0;  //83 / 230 = 0
    16'b01010011_11100111 : OUT <= 0;  //83 / 231 = 0
    16'b01010011_11101000 : OUT <= 0;  //83 / 232 = 0
    16'b01010011_11101001 : OUT <= 0;  //83 / 233 = 0
    16'b01010011_11101010 : OUT <= 0;  //83 / 234 = 0
    16'b01010011_11101011 : OUT <= 0;  //83 / 235 = 0
    16'b01010011_11101100 : OUT <= 0;  //83 / 236 = 0
    16'b01010011_11101101 : OUT <= 0;  //83 / 237 = 0
    16'b01010011_11101110 : OUT <= 0;  //83 / 238 = 0
    16'b01010011_11101111 : OUT <= 0;  //83 / 239 = 0
    16'b01010011_11110000 : OUT <= 0;  //83 / 240 = 0
    16'b01010011_11110001 : OUT <= 0;  //83 / 241 = 0
    16'b01010011_11110010 : OUT <= 0;  //83 / 242 = 0
    16'b01010011_11110011 : OUT <= 0;  //83 / 243 = 0
    16'b01010011_11110100 : OUT <= 0;  //83 / 244 = 0
    16'b01010011_11110101 : OUT <= 0;  //83 / 245 = 0
    16'b01010011_11110110 : OUT <= 0;  //83 / 246 = 0
    16'b01010011_11110111 : OUT <= 0;  //83 / 247 = 0
    16'b01010011_11111000 : OUT <= 0;  //83 / 248 = 0
    16'b01010011_11111001 : OUT <= 0;  //83 / 249 = 0
    16'b01010011_11111010 : OUT <= 0;  //83 / 250 = 0
    16'b01010011_11111011 : OUT <= 0;  //83 / 251 = 0
    16'b01010011_11111100 : OUT <= 0;  //83 / 252 = 0
    16'b01010011_11111101 : OUT <= 0;  //83 / 253 = 0
    16'b01010011_11111110 : OUT <= 0;  //83 / 254 = 0
    16'b01010011_11111111 : OUT <= 0;  //83 / 255 = 0
    16'b01010100_00000000 : OUT <= 0;  //84 / 0 = 0
    16'b01010100_00000001 : OUT <= 84;  //84 / 1 = 84
    16'b01010100_00000010 : OUT <= 42;  //84 / 2 = 42
    16'b01010100_00000011 : OUT <= 28;  //84 / 3 = 28
    16'b01010100_00000100 : OUT <= 21;  //84 / 4 = 21
    16'b01010100_00000101 : OUT <= 16;  //84 / 5 = 16
    16'b01010100_00000110 : OUT <= 14;  //84 / 6 = 14
    16'b01010100_00000111 : OUT <= 12;  //84 / 7 = 12
    16'b01010100_00001000 : OUT <= 10;  //84 / 8 = 10
    16'b01010100_00001001 : OUT <= 9;  //84 / 9 = 9
    16'b01010100_00001010 : OUT <= 8;  //84 / 10 = 8
    16'b01010100_00001011 : OUT <= 7;  //84 / 11 = 7
    16'b01010100_00001100 : OUT <= 7;  //84 / 12 = 7
    16'b01010100_00001101 : OUT <= 6;  //84 / 13 = 6
    16'b01010100_00001110 : OUT <= 6;  //84 / 14 = 6
    16'b01010100_00001111 : OUT <= 5;  //84 / 15 = 5
    16'b01010100_00010000 : OUT <= 5;  //84 / 16 = 5
    16'b01010100_00010001 : OUT <= 4;  //84 / 17 = 4
    16'b01010100_00010010 : OUT <= 4;  //84 / 18 = 4
    16'b01010100_00010011 : OUT <= 4;  //84 / 19 = 4
    16'b01010100_00010100 : OUT <= 4;  //84 / 20 = 4
    16'b01010100_00010101 : OUT <= 4;  //84 / 21 = 4
    16'b01010100_00010110 : OUT <= 3;  //84 / 22 = 3
    16'b01010100_00010111 : OUT <= 3;  //84 / 23 = 3
    16'b01010100_00011000 : OUT <= 3;  //84 / 24 = 3
    16'b01010100_00011001 : OUT <= 3;  //84 / 25 = 3
    16'b01010100_00011010 : OUT <= 3;  //84 / 26 = 3
    16'b01010100_00011011 : OUT <= 3;  //84 / 27 = 3
    16'b01010100_00011100 : OUT <= 3;  //84 / 28 = 3
    16'b01010100_00011101 : OUT <= 2;  //84 / 29 = 2
    16'b01010100_00011110 : OUT <= 2;  //84 / 30 = 2
    16'b01010100_00011111 : OUT <= 2;  //84 / 31 = 2
    16'b01010100_00100000 : OUT <= 2;  //84 / 32 = 2
    16'b01010100_00100001 : OUT <= 2;  //84 / 33 = 2
    16'b01010100_00100010 : OUT <= 2;  //84 / 34 = 2
    16'b01010100_00100011 : OUT <= 2;  //84 / 35 = 2
    16'b01010100_00100100 : OUT <= 2;  //84 / 36 = 2
    16'b01010100_00100101 : OUT <= 2;  //84 / 37 = 2
    16'b01010100_00100110 : OUT <= 2;  //84 / 38 = 2
    16'b01010100_00100111 : OUT <= 2;  //84 / 39 = 2
    16'b01010100_00101000 : OUT <= 2;  //84 / 40 = 2
    16'b01010100_00101001 : OUT <= 2;  //84 / 41 = 2
    16'b01010100_00101010 : OUT <= 2;  //84 / 42 = 2
    16'b01010100_00101011 : OUT <= 1;  //84 / 43 = 1
    16'b01010100_00101100 : OUT <= 1;  //84 / 44 = 1
    16'b01010100_00101101 : OUT <= 1;  //84 / 45 = 1
    16'b01010100_00101110 : OUT <= 1;  //84 / 46 = 1
    16'b01010100_00101111 : OUT <= 1;  //84 / 47 = 1
    16'b01010100_00110000 : OUT <= 1;  //84 / 48 = 1
    16'b01010100_00110001 : OUT <= 1;  //84 / 49 = 1
    16'b01010100_00110010 : OUT <= 1;  //84 / 50 = 1
    16'b01010100_00110011 : OUT <= 1;  //84 / 51 = 1
    16'b01010100_00110100 : OUT <= 1;  //84 / 52 = 1
    16'b01010100_00110101 : OUT <= 1;  //84 / 53 = 1
    16'b01010100_00110110 : OUT <= 1;  //84 / 54 = 1
    16'b01010100_00110111 : OUT <= 1;  //84 / 55 = 1
    16'b01010100_00111000 : OUT <= 1;  //84 / 56 = 1
    16'b01010100_00111001 : OUT <= 1;  //84 / 57 = 1
    16'b01010100_00111010 : OUT <= 1;  //84 / 58 = 1
    16'b01010100_00111011 : OUT <= 1;  //84 / 59 = 1
    16'b01010100_00111100 : OUT <= 1;  //84 / 60 = 1
    16'b01010100_00111101 : OUT <= 1;  //84 / 61 = 1
    16'b01010100_00111110 : OUT <= 1;  //84 / 62 = 1
    16'b01010100_00111111 : OUT <= 1;  //84 / 63 = 1
    16'b01010100_01000000 : OUT <= 1;  //84 / 64 = 1
    16'b01010100_01000001 : OUT <= 1;  //84 / 65 = 1
    16'b01010100_01000010 : OUT <= 1;  //84 / 66 = 1
    16'b01010100_01000011 : OUT <= 1;  //84 / 67 = 1
    16'b01010100_01000100 : OUT <= 1;  //84 / 68 = 1
    16'b01010100_01000101 : OUT <= 1;  //84 / 69 = 1
    16'b01010100_01000110 : OUT <= 1;  //84 / 70 = 1
    16'b01010100_01000111 : OUT <= 1;  //84 / 71 = 1
    16'b01010100_01001000 : OUT <= 1;  //84 / 72 = 1
    16'b01010100_01001001 : OUT <= 1;  //84 / 73 = 1
    16'b01010100_01001010 : OUT <= 1;  //84 / 74 = 1
    16'b01010100_01001011 : OUT <= 1;  //84 / 75 = 1
    16'b01010100_01001100 : OUT <= 1;  //84 / 76 = 1
    16'b01010100_01001101 : OUT <= 1;  //84 / 77 = 1
    16'b01010100_01001110 : OUT <= 1;  //84 / 78 = 1
    16'b01010100_01001111 : OUT <= 1;  //84 / 79 = 1
    16'b01010100_01010000 : OUT <= 1;  //84 / 80 = 1
    16'b01010100_01010001 : OUT <= 1;  //84 / 81 = 1
    16'b01010100_01010010 : OUT <= 1;  //84 / 82 = 1
    16'b01010100_01010011 : OUT <= 1;  //84 / 83 = 1
    16'b01010100_01010100 : OUT <= 1;  //84 / 84 = 1
    16'b01010100_01010101 : OUT <= 0;  //84 / 85 = 0
    16'b01010100_01010110 : OUT <= 0;  //84 / 86 = 0
    16'b01010100_01010111 : OUT <= 0;  //84 / 87 = 0
    16'b01010100_01011000 : OUT <= 0;  //84 / 88 = 0
    16'b01010100_01011001 : OUT <= 0;  //84 / 89 = 0
    16'b01010100_01011010 : OUT <= 0;  //84 / 90 = 0
    16'b01010100_01011011 : OUT <= 0;  //84 / 91 = 0
    16'b01010100_01011100 : OUT <= 0;  //84 / 92 = 0
    16'b01010100_01011101 : OUT <= 0;  //84 / 93 = 0
    16'b01010100_01011110 : OUT <= 0;  //84 / 94 = 0
    16'b01010100_01011111 : OUT <= 0;  //84 / 95 = 0
    16'b01010100_01100000 : OUT <= 0;  //84 / 96 = 0
    16'b01010100_01100001 : OUT <= 0;  //84 / 97 = 0
    16'b01010100_01100010 : OUT <= 0;  //84 / 98 = 0
    16'b01010100_01100011 : OUT <= 0;  //84 / 99 = 0
    16'b01010100_01100100 : OUT <= 0;  //84 / 100 = 0
    16'b01010100_01100101 : OUT <= 0;  //84 / 101 = 0
    16'b01010100_01100110 : OUT <= 0;  //84 / 102 = 0
    16'b01010100_01100111 : OUT <= 0;  //84 / 103 = 0
    16'b01010100_01101000 : OUT <= 0;  //84 / 104 = 0
    16'b01010100_01101001 : OUT <= 0;  //84 / 105 = 0
    16'b01010100_01101010 : OUT <= 0;  //84 / 106 = 0
    16'b01010100_01101011 : OUT <= 0;  //84 / 107 = 0
    16'b01010100_01101100 : OUT <= 0;  //84 / 108 = 0
    16'b01010100_01101101 : OUT <= 0;  //84 / 109 = 0
    16'b01010100_01101110 : OUT <= 0;  //84 / 110 = 0
    16'b01010100_01101111 : OUT <= 0;  //84 / 111 = 0
    16'b01010100_01110000 : OUT <= 0;  //84 / 112 = 0
    16'b01010100_01110001 : OUT <= 0;  //84 / 113 = 0
    16'b01010100_01110010 : OUT <= 0;  //84 / 114 = 0
    16'b01010100_01110011 : OUT <= 0;  //84 / 115 = 0
    16'b01010100_01110100 : OUT <= 0;  //84 / 116 = 0
    16'b01010100_01110101 : OUT <= 0;  //84 / 117 = 0
    16'b01010100_01110110 : OUT <= 0;  //84 / 118 = 0
    16'b01010100_01110111 : OUT <= 0;  //84 / 119 = 0
    16'b01010100_01111000 : OUT <= 0;  //84 / 120 = 0
    16'b01010100_01111001 : OUT <= 0;  //84 / 121 = 0
    16'b01010100_01111010 : OUT <= 0;  //84 / 122 = 0
    16'b01010100_01111011 : OUT <= 0;  //84 / 123 = 0
    16'b01010100_01111100 : OUT <= 0;  //84 / 124 = 0
    16'b01010100_01111101 : OUT <= 0;  //84 / 125 = 0
    16'b01010100_01111110 : OUT <= 0;  //84 / 126 = 0
    16'b01010100_01111111 : OUT <= 0;  //84 / 127 = 0
    16'b01010100_10000000 : OUT <= 0;  //84 / 128 = 0
    16'b01010100_10000001 : OUT <= 0;  //84 / 129 = 0
    16'b01010100_10000010 : OUT <= 0;  //84 / 130 = 0
    16'b01010100_10000011 : OUT <= 0;  //84 / 131 = 0
    16'b01010100_10000100 : OUT <= 0;  //84 / 132 = 0
    16'b01010100_10000101 : OUT <= 0;  //84 / 133 = 0
    16'b01010100_10000110 : OUT <= 0;  //84 / 134 = 0
    16'b01010100_10000111 : OUT <= 0;  //84 / 135 = 0
    16'b01010100_10001000 : OUT <= 0;  //84 / 136 = 0
    16'b01010100_10001001 : OUT <= 0;  //84 / 137 = 0
    16'b01010100_10001010 : OUT <= 0;  //84 / 138 = 0
    16'b01010100_10001011 : OUT <= 0;  //84 / 139 = 0
    16'b01010100_10001100 : OUT <= 0;  //84 / 140 = 0
    16'b01010100_10001101 : OUT <= 0;  //84 / 141 = 0
    16'b01010100_10001110 : OUT <= 0;  //84 / 142 = 0
    16'b01010100_10001111 : OUT <= 0;  //84 / 143 = 0
    16'b01010100_10010000 : OUT <= 0;  //84 / 144 = 0
    16'b01010100_10010001 : OUT <= 0;  //84 / 145 = 0
    16'b01010100_10010010 : OUT <= 0;  //84 / 146 = 0
    16'b01010100_10010011 : OUT <= 0;  //84 / 147 = 0
    16'b01010100_10010100 : OUT <= 0;  //84 / 148 = 0
    16'b01010100_10010101 : OUT <= 0;  //84 / 149 = 0
    16'b01010100_10010110 : OUT <= 0;  //84 / 150 = 0
    16'b01010100_10010111 : OUT <= 0;  //84 / 151 = 0
    16'b01010100_10011000 : OUT <= 0;  //84 / 152 = 0
    16'b01010100_10011001 : OUT <= 0;  //84 / 153 = 0
    16'b01010100_10011010 : OUT <= 0;  //84 / 154 = 0
    16'b01010100_10011011 : OUT <= 0;  //84 / 155 = 0
    16'b01010100_10011100 : OUT <= 0;  //84 / 156 = 0
    16'b01010100_10011101 : OUT <= 0;  //84 / 157 = 0
    16'b01010100_10011110 : OUT <= 0;  //84 / 158 = 0
    16'b01010100_10011111 : OUT <= 0;  //84 / 159 = 0
    16'b01010100_10100000 : OUT <= 0;  //84 / 160 = 0
    16'b01010100_10100001 : OUT <= 0;  //84 / 161 = 0
    16'b01010100_10100010 : OUT <= 0;  //84 / 162 = 0
    16'b01010100_10100011 : OUT <= 0;  //84 / 163 = 0
    16'b01010100_10100100 : OUT <= 0;  //84 / 164 = 0
    16'b01010100_10100101 : OUT <= 0;  //84 / 165 = 0
    16'b01010100_10100110 : OUT <= 0;  //84 / 166 = 0
    16'b01010100_10100111 : OUT <= 0;  //84 / 167 = 0
    16'b01010100_10101000 : OUT <= 0;  //84 / 168 = 0
    16'b01010100_10101001 : OUT <= 0;  //84 / 169 = 0
    16'b01010100_10101010 : OUT <= 0;  //84 / 170 = 0
    16'b01010100_10101011 : OUT <= 0;  //84 / 171 = 0
    16'b01010100_10101100 : OUT <= 0;  //84 / 172 = 0
    16'b01010100_10101101 : OUT <= 0;  //84 / 173 = 0
    16'b01010100_10101110 : OUT <= 0;  //84 / 174 = 0
    16'b01010100_10101111 : OUT <= 0;  //84 / 175 = 0
    16'b01010100_10110000 : OUT <= 0;  //84 / 176 = 0
    16'b01010100_10110001 : OUT <= 0;  //84 / 177 = 0
    16'b01010100_10110010 : OUT <= 0;  //84 / 178 = 0
    16'b01010100_10110011 : OUT <= 0;  //84 / 179 = 0
    16'b01010100_10110100 : OUT <= 0;  //84 / 180 = 0
    16'b01010100_10110101 : OUT <= 0;  //84 / 181 = 0
    16'b01010100_10110110 : OUT <= 0;  //84 / 182 = 0
    16'b01010100_10110111 : OUT <= 0;  //84 / 183 = 0
    16'b01010100_10111000 : OUT <= 0;  //84 / 184 = 0
    16'b01010100_10111001 : OUT <= 0;  //84 / 185 = 0
    16'b01010100_10111010 : OUT <= 0;  //84 / 186 = 0
    16'b01010100_10111011 : OUT <= 0;  //84 / 187 = 0
    16'b01010100_10111100 : OUT <= 0;  //84 / 188 = 0
    16'b01010100_10111101 : OUT <= 0;  //84 / 189 = 0
    16'b01010100_10111110 : OUT <= 0;  //84 / 190 = 0
    16'b01010100_10111111 : OUT <= 0;  //84 / 191 = 0
    16'b01010100_11000000 : OUT <= 0;  //84 / 192 = 0
    16'b01010100_11000001 : OUT <= 0;  //84 / 193 = 0
    16'b01010100_11000010 : OUT <= 0;  //84 / 194 = 0
    16'b01010100_11000011 : OUT <= 0;  //84 / 195 = 0
    16'b01010100_11000100 : OUT <= 0;  //84 / 196 = 0
    16'b01010100_11000101 : OUT <= 0;  //84 / 197 = 0
    16'b01010100_11000110 : OUT <= 0;  //84 / 198 = 0
    16'b01010100_11000111 : OUT <= 0;  //84 / 199 = 0
    16'b01010100_11001000 : OUT <= 0;  //84 / 200 = 0
    16'b01010100_11001001 : OUT <= 0;  //84 / 201 = 0
    16'b01010100_11001010 : OUT <= 0;  //84 / 202 = 0
    16'b01010100_11001011 : OUT <= 0;  //84 / 203 = 0
    16'b01010100_11001100 : OUT <= 0;  //84 / 204 = 0
    16'b01010100_11001101 : OUT <= 0;  //84 / 205 = 0
    16'b01010100_11001110 : OUT <= 0;  //84 / 206 = 0
    16'b01010100_11001111 : OUT <= 0;  //84 / 207 = 0
    16'b01010100_11010000 : OUT <= 0;  //84 / 208 = 0
    16'b01010100_11010001 : OUT <= 0;  //84 / 209 = 0
    16'b01010100_11010010 : OUT <= 0;  //84 / 210 = 0
    16'b01010100_11010011 : OUT <= 0;  //84 / 211 = 0
    16'b01010100_11010100 : OUT <= 0;  //84 / 212 = 0
    16'b01010100_11010101 : OUT <= 0;  //84 / 213 = 0
    16'b01010100_11010110 : OUT <= 0;  //84 / 214 = 0
    16'b01010100_11010111 : OUT <= 0;  //84 / 215 = 0
    16'b01010100_11011000 : OUT <= 0;  //84 / 216 = 0
    16'b01010100_11011001 : OUT <= 0;  //84 / 217 = 0
    16'b01010100_11011010 : OUT <= 0;  //84 / 218 = 0
    16'b01010100_11011011 : OUT <= 0;  //84 / 219 = 0
    16'b01010100_11011100 : OUT <= 0;  //84 / 220 = 0
    16'b01010100_11011101 : OUT <= 0;  //84 / 221 = 0
    16'b01010100_11011110 : OUT <= 0;  //84 / 222 = 0
    16'b01010100_11011111 : OUT <= 0;  //84 / 223 = 0
    16'b01010100_11100000 : OUT <= 0;  //84 / 224 = 0
    16'b01010100_11100001 : OUT <= 0;  //84 / 225 = 0
    16'b01010100_11100010 : OUT <= 0;  //84 / 226 = 0
    16'b01010100_11100011 : OUT <= 0;  //84 / 227 = 0
    16'b01010100_11100100 : OUT <= 0;  //84 / 228 = 0
    16'b01010100_11100101 : OUT <= 0;  //84 / 229 = 0
    16'b01010100_11100110 : OUT <= 0;  //84 / 230 = 0
    16'b01010100_11100111 : OUT <= 0;  //84 / 231 = 0
    16'b01010100_11101000 : OUT <= 0;  //84 / 232 = 0
    16'b01010100_11101001 : OUT <= 0;  //84 / 233 = 0
    16'b01010100_11101010 : OUT <= 0;  //84 / 234 = 0
    16'b01010100_11101011 : OUT <= 0;  //84 / 235 = 0
    16'b01010100_11101100 : OUT <= 0;  //84 / 236 = 0
    16'b01010100_11101101 : OUT <= 0;  //84 / 237 = 0
    16'b01010100_11101110 : OUT <= 0;  //84 / 238 = 0
    16'b01010100_11101111 : OUT <= 0;  //84 / 239 = 0
    16'b01010100_11110000 : OUT <= 0;  //84 / 240 = 0
    16'b01010100_11110001 : OUT <= 0;  //84 / 241 = 0
    16'b01010100_11110010 : OUT <= 0;  //84 / 242 = 0
    16'b01010100_11110011 : OUT <= 0;  //84 / 243 = 0
    16'b01010100_11110100 : OUT <= 0;  //84 / 244 = 0
    16'b01010100_11110101 : OUT <= 0;  //84 / 245 = 0
    16'b01010100_11110110 : OUT <= 0;  //84 / 246 = 0
    16'b01010100_11110111 : OUT <= 0;  //84 / 247 = 0
    16'b01010100_11111000 : OUT <= 0;  //84 / 248 = 0
    16'b01010100_11111001 : OUT <= 0;  //84 / 249 = 0
    16'b01010100_11111010 : OUT <= 0;  //84 / 250 = 0
    16'b01010100_11111011 : OUT <= 0;  //84 / 251 = 0
    16'b01010100_11111100 : OUT <= 0;  //84 / 252 = 0
    16'b01010100_11111101 : OUT <= 0;  //84 / 253 = 0
    16'b01010100_11111110 : OUT <= 0;  //84 / 254 = 0
    16'b01010100_11111111 : OUT <= 0;  //84 / 255 = 0
    16'b01010101_00000000 : OUT <= 0;  //85 / 0 = 0
    16'b01010101_00000001 : OUT <= 85;  //85 / 1 = 85
    16'b01010101_00000010 : OUT <= 42;  //85 / 2 = 42
    16'b01010101_00000011 : OUT <= 28;  //85 / 3 = 28
    16'b01010101_00000100 : OUT <= 21;  //85 / 4 = 21
    16'b01010101_00000101 : OUT <= 17;  //85 / 5 = 17
    16'b01010101_00000110 : OUT <= 14;  //85 / 6 = 14
    16'b01010101_00000111 : OUT <= 12;  //85 / 7 = 12
    16'b01010101_00001000 : OUT <= 10;  //85 / 8 = 10
    16'b01010101_00001001 : OUT <= 9;  //85 / 9 = 9
    16'b01010101_00001010 : OUT <= 8;  //85 / 10 = 8
    16'b01010101_00001011 : OUT <= 7;  //85 / 11 = 7
    16'b01010101_00001100 : OUT <= 7;  //85 / 12 = 7
    16'b01010101_00001101 : OUT <= 6;  //85 / 13 = 6
    16'b01010101_00001110 : OUT <= 6;  //85 / 14 = 6
    16'b01010101_00001111 : OUT <= 5;  //85 / 15 = 5
    16'b01010101_00010000 : OUT <= 5;  //85 / 16 = 5
    16'b01010101_00010001 : OUT <= 5;  //85 / 17 = 5
    16'b01010101_00010010 : OUT <= 4;  //85 / 18 = 4
    16'b01010101_00010011 : OUT <= 4;  //85 / 19 = 4
    16'b01010101_00010100 : OUT <= 4;  //85 / 20 = 4
    16'b01010101_00010101 : OUT <= 4;  //85 / 21 = 4
    16'b01010101_00010110 : OUT <= 3;  //85 / 22 = 3
    16'b01010101_00010111 : OUT <= 3;  //85 / 23 = 3
    16'b01010101_00011000 : OUT <= 3;  //85 / 24 = 3
    16'b01010101_00011001 : OUT <= 3;  //85 / 25 = 3
    16'b01010101_00011010 : OUT <= 3;  //85 / 26 = 3
    16'b01010101_00011011 : OUT <= 3;  //85 / 27 = 3
    16'b01010101_00011100 : OUT <= 3;  //85 / 28 = 3
    16'b01010101_00011101 : OUT <= 2;  //85 / 29 = 2
    16'b01010101_00011110 : OUT <= 2;  //85 / 30 = 2
    16'b01010101_00011111 : OUT <= 2;  //85 / 31 = 2
    16'b01010101_00100000 : OUT <= 2;  //85 / 32 = 2
    16'b01010101_00100001 : OUT <= 2;  //85 / 33 = 2
    16'b01010101_00100010 : OUT <= 2;  //85 / 34 = 2
    16'b01010101_00100011 : OUT <= 2;  //85 / 35 = 2
    16'b01010101_00100100 : OUT <= 2;  //85 / 36 = 2
    16'b01010101_00100101 : OUT <= 2;  //85 / 37 = 2
    16'b01010101_00100110 : OUT <= 2;  //85 / 38 = 2
    16'b01010101_00100111 : OUT <= 2;  //85 / 39 = 2
    16'b01010101_00101000 : OUT <= 2;  //85 / 40 = 2
    16'b01010101_00101001 : OUT <= 2;  //85 / 41 = 2
    16'b01010101_00101010 : OUT <= 2;  //85 / 42 = 2
    16'b01010101_00101011 : OUT <= 1;  //85 / 43 = 1
    16'b01010101_00101100 : OUT <= 1;  //85 / 44 = 1
    16'b01010101_00101101 : OUT <= 1;  //85 / 45 = 1
    16'b01010101_00101110 : OUT <= 1;  //85 / 46 = 1
    16'b01010101_00101111 : OUT <= 1;  //85 / 47 = 1
    16'b01010101_00110000 : OUT <= 1;  //85 / 48 = 1
    16'b01010101_00110001 : OUT <= 1;  //85 / 49 = 1
    16'b01010101_00110010 : OUT <= 1;  //85 / 50 = 1
    16'b01010101_00110011 : OUT <= 1;  //85 / 51 = 1
    16'b01010101_00110100 : OUT <= 1;  //85 / 52 = 1
    16'b01010101_00110101 : OUT <= 1;  //85 / 53 = 1
    16'b01010101_00110110 : OUT <= 1;  //85 / 54 = 1
    16'b01010101_00110111 : OUT <= 1;  //85 / 55 = 1
    16'b01010101_00111000 : OUT <= 1;  //85 / 56 = 1
    16'b01010101_00111001 : OUT <= 1;  //85 / 57 = 1
    16'b01010101_00111010 : OUT <= 1;  //85 / 58 = 1
    16'b01010101_00111011 : OUT <= 1;  //85 / 59 = 1
    16'b01010101_00111100 : OUT <= 1;  //85 / 60 = 1
    16'b01010101_00111101 : OUT <= 1;  //85 / 61 = 1
    16'b01010101_00111110 : OUT <= 1;  //85 / 62 = 1
    16'b01010101_00111111 : OUT <= 1;  //85 / 63 = 1
    16'b01010101_01000000 : OUT <= 1;  //85 / 64 = 1
    16'b01010101_01000001 : OUT <= 1;  //85 / 65 = 1
    16'b01010101_01000010 : OUT <= 1;  //85 / 66 = 1
    16'b01010101_01000011 : OUT <= 1;  //85 / 67 = 1
    16'b01010101_01000100 : OUT <= 1;  //85 / 68 = 1
    16'b01010101_01000101 : OUT <= 1;  //85 / 69 = 1
    16'b01010101_01000110 : OUT <= 1;  //85 / 70 = 1
    16'b01010101_01000111 : OUT <= 1;  //85 / 71 = 1
    16'b01010101_01001000 : OUT <= 1;  //85 / 72 = 1
    16'b01010101_01001001 : OUT <= 1;  //85 / 73 = 1
    16'b01010101_01001010 : OUT <= 1;  //85 / 74 = 1
    16'b01010101_01001011 : OUT <= 1;  //85 / 75 = 1
    16'b01010101_01001100 : OUT <= 1;  //85 / 76 = 1
    16'b01010101_01001101 : OUT <= 1;  //85 / 77 = 1
    16'b01010101_01001110 : OUT <= 1;  //85 / 78 = 1
    16'b01010101_01001111 : OUT <= 1;  //85 / 79 = 1
    16'b01010101_01010000 : OUT <= 1;  //85 / 80 = 1
    16'b01010101_01010001 : OUT <= 1;  //85 / 81 = 1
    16'b01010101_01010010 : OUT <= 1;  //85 / 82 = 1
    16'b01010101_01010011 : OUT <= 1;  //85 / 83 = 1
    16'b01010101_01010100 : OUT <= 1;  //85 / 84 = 1
    16'b01010101_01010101 : OUT <= 1;  //85 / 85 = 1
    16'b01010101_01010110 : OUT <= 0;  //85 / 86 = 0
    16'b01010101_01010111 : OUT <= 0;  //85 / 87 = 0
    16'b01010101_01011000 : OUT <= 0;  //85 / 88 = 0
    16'b01010101_01011001 : OUT <= 0;  //85 / 89 = 0
    16'b01010101_01011010 : OUT <= 0;  //85 / 90 = 0
    16'b01010101_01011011 : OUT <= 0;  //85 / 91 = 0
    16'b01010101_01011100 : OUT <= 0;  //85 / 92 = 0
    16'b01010101_01011101 : OUT <= 0;  //85 / 93 = 0
    16'b01010101_01011110 : OUT <= 0;  //85 / 94 = 0
    16'b01010101_01011111 : OUT <= 0;  //85 / 95 = 0
    16'b01010101_01100000 : OUT <= 0;  //85 / 96 = 0
    16'b01010101_01100001 : OUT <= 0;  //85 / 97 = 0
    16'b01010101_01100010 : OUT <= 0;  //85 / 98 = 0
    16'b01010101_01100011 : OUT <= 0;  //85 / 99 = 0
    16'b01010101_01100100 : OUT <= 0;  //85 / 100 = 0
    16'b01010101_01100101 : OUT <= 0;  //85 / 101 = 0
    16'b01010101_01100110 : OUT <= 0;  //85 / 102 = 0
    16'b01010101_01100111 : OUT <= 0;  //85 / 103 = 0
    16'b01010101_01101000 : OUT <= 0;  //85 / 104 = 0
    16'b01010101_01101001 : OUT <= 0;  //85 / 105 = 0
    16'b01010101_01101010 : OUT <= 0;  //85 / 106 = 0
    16'b01010101_01101011 : OUT <= 0;  //85 / 107 = 0
    16'b01010101_01101100 : OUT <= 0;  //85 / 108 = 0
    16'b01010101_01101101 : OUT <= 0;  //85 / 109 = 0
    16'b01010101_01101110 : OUT <= 0;  //85 / 110 = 0
    16'b01010101_01101111 : OUT <= 0;  //85 / 111 = 0
    16'b01010101_01110000 : OUT <= 0;  //85 / 112 = 0
    16'b01010101_01110001 : OUT <= 0;  //85 / 113 = 0
    16'b01010101_01110010 : OUT <= 0;  //85 / 114 = 0
    16'b01010101_01110011 : OUT <= 0;  //85 / 115 = 0
    16'b01010101_01110100 : OUT <= 0;  //85 / 116 = 0
    16'b01010101_01110101 : OUT <= 0;  //85 / 117 = 0
    16'b01010101_01110110 : OUT <= 0;  //85 / 118 = 0
    16'b01010101_01110111 : OUT <= 0;  //85 / 119 = 0
    16'b01010101_01111000 : OUT <= 0;  //85 / 120 = 0
    16'b01010101_01111001 : OUT <= 0;  //85 / 121 = 0
    16'b01010101_01111010 : OUT <= 0;  //85 / 122 = 0
    16'b01010101_01111011 : OUT <= 0;  //85 / 123 = 0
    16'b01010101_01111100 : OUT <= 0;  //85 / 124 = 0
    16'b01010101_01111101 : OUT <= 0;  //85 / 125 = 0
    16'b01010101_01111110 : OUT <= 0;  //85 / 126 = 0
    16'b01010101_01111111 : OUT <= 0;  //85 / 127 = 0
    16'b01010101_10000000 : OUT <= 0;  //85 / 128 = 0
    16'b01010101_10000001 : OUT <= 0;  //85 / 129 = 0
    16'b01010101_10000010 : OUT <= 0;  //85 / 130 = 0
    16'b01010101_10000011 : OUT <= 0;  //85 / 131 = 0
    16'b01010101_10000100 : OUT <= 0;  //85 / 132 = 0
    16'b01010101_10000101 : OUT <= 0;  //85 / 133 = 0
    16'b01010101_10000110 : OUT <= 0;  //85 / 134 = 0
    16'b01010101_10000111 : OUT <= 0;  //85 / 135 = 0
    16'b01010101_10001000 : OUT <= 0;  //85 / 136 = 0
    16'b01010101_10001001 : OUT <= 0;  //85 / 137 = 0
    16'b01010101_10001010 : OUT <= 0;  //85 / 138 = 0
    16'b01010101_10001011 : OUT <= 0;  //85 / 139 = 0
    16'b01010101_10001100 : OUT <= 0;  //85 / 140 = 0
    16'b01010101_10001101 : OUT <= 0;  //85 / 141 = 0
    16'b01010101_10001110 : OUT <= 0;  //85 / 142 = 0
    16'b01010101_10001111 : OUT <= 0;  //85 / 143 = 0
    16'b01010101_10010000 : OUT <= 0;  //85 / 144 = 0
    16'b01010101_10010001 : OUT <= 0;  //85 / 145 = 0
    16'b01010101_10010010 : OUT <= 0;  //85 / 146 = 0
    16'b01010101_10010011 : OUT <= 0;  //85 / 147 = 0
    16'b01010101_10010100 : OUT <= 0;  //85 / 148 = 0
    16'b01010101_10010101 : OUT <= 0;  //85 / 149 = 0
    16'b01010101_10010110 : OUT <= 0;  //85 / 150 = 0
    16'b01010101_10010111 : OUT <= 0;  //85 / 151 = 0
    16'b01010101_10011000 : OUT <= 0;  //85 / 152 = 0
    16'b01010101_10011001 : OUT <= 0;  //85 / 153 = 0
    16'b01010101_10011010 : OUT <= 0;  //85 / 154 = 0
    16'b01010101_10011011 : OUT <= 0;  //85 / 155 = 0
    16'b01010101_10011100 : OUT <= 0;  //85 / 156 = 0
    16'b01010101_10011101 : OUT <= 0;  //85 / 157 = 0
    16'b01010101_10011110 : OUT <= 0;  //85 / 158 = 0
    16'b01010101_10011111 : OUT <= 0;  //85 / 159 = 0
    16'b01010101_10100000 : OUT <= 0;  //85 / 160 = 0
    16'b01010101_10100001 : OUT <= 0;  //85 / 161 = 0
    16'b01010101_10100010 : OUT <= 0;  //85 / 162 = 0
    16'b01010101_10100011 : OUT <= 0;  //85 / 163 = 0
    16'b01010101_10100100 : OUT <= 0;  //85 / 164 = 0
    16'b01010101_10100101 : OUT <= 0;  //85 / 165 = 0
    16'b01010101_10100110 : OUT <= 0;  //85 / 166 = 0
    16'b01010101_10100111 : OUT <= 0;  //85 / 167 = 0
    16'b01010101_10101000 : OUT <= 0;  //85 / 168 = 0
    16'b01010101_10101001 : OUT <= 0;  //85 / 169 = 0
    16'b01010101_10101010 : OUT <= 0;  //85 / 170 = 0
    16'b01010101_10101011 : OUT <= 0;  //85 / 171 = 0
    16'b01010101_10101100 : OUT <= 0;  //85 / 172 = 0
    16'b01010101_10101101 : OUT <= 0;  //85 / 173 = 0
    16'b01010101_10101110 : OUT <= 0;  //85 / 174 = 0
    16'b01010101_10101111 : OUT <= 0;  //85 / 175 = 0
    16'b01010101_10110000 : OUT <= 0;  //85 / 176 = 0
    16'b01010101_10110001 : OUT <= 0;  //85 / 177 = 0
    16'b01010101_10110010 : OUT <= 0;  //85 / 178 = 0
    16'b01010101_10110011 : OUT <= 0;  //85 / 179 = 0
    16'b01010101_10110100 : OUT <= 0;  //85 / 180 = 0
    16'b01010101_10110101 : OUT <= 0;  //85 / 181 = 0
    16'b01010101_10110110 : OUT <= 0;  //85 / 182 = 0
    16'b01010101_10110111 : OUT <= 0;  //85 / 183 = 0
    16'b01010101_10111000 : OUT <= 0;  //85 / 184 = 0
    16'b01010101_10111001 : OUT <= 0;  //85 / 185 = 0
    16'b01010101_10111010 : OUT <= 0;  //85 / 186 = 0
    16'b01010101_10111011 : OUT <= 0;  //85 / 187 = 0
    16'b01010101_10111100 : OUT <= 0;  //85 / 188 = 0
    16'b01010101_10111101 : OUT <= 0;  //85 / 189 = 0
    16'b01010101_10111110 : OUT <= 0;  //85 / 190 = 0
    16'b01010101_10111111 : OUT <= 0;  //85 / 191 = 0
    16'b01010101_11000000 : OUT <= 0;  //85 / 192 = 0
    16'b01010101_11000001 : OUT <= 0;  //85 / 193 = 0
    16'b01010101_11000010 : OUT <= 0;  //85 / 194 = 0
    16'b01010101_11000011 : OUT <= 0;  //85 / 195 = 0
    16'b01010101_11000100 : OUT <= 0;  //85 / 196 = 0
    16'b01010101_11000101 : OUT <= 0;  //85 / 197 = 0
    16'b01010101_11000110 : OUT <= 0;  //85 / 198 = 0
    16'b01010101_11000111 : OUT <= 0;  //85 / 199 = 0
    16'b01010101_11001000 : OUT <= 0;  //85 / 200 = 0
    16'b01010101_11001001 : OUT <= 0;  //85 / 201 = 0
    16'b01010101_11001010 : OUT <= 0;  //85 / 202 = 0
    16'b01010101_11001011 : OUT <= 0;  //85 / 203 = 0
    16'b01010101_11001100 : OUT <= 0;  //85 / 204 = 0
    16'b01010101_11001101 : OUT <= 0;  //85 / 205 = 0
    16'b01010101_11001110 : OUT <= 0;  //85 / 206 = 0
    16'b01010101_11001111 : OUT <= 0;  //85 / 207 = 0
    16'b01010101_11010000 : OUT <= 0;  //85 / 208 = 0
    16'b01010101_11010001 : OUT <= 0;  //85 / 209 = 0
    16'b01010101_11010010 : OUT <= 0;  //85 / 210 = 0
    16'b01010101_11010011 : OUT <= 0;  //85 / 211 = 0
    16'b01010101_11010100 : OUT <= 0;  //85 / 212 = 0
    16'b01010101_11010101 : OUT <= 0;  //85 / 213 = 0
    16'b01010101_11010110 : OUT <= 0;  //85 / 214 = 0
    16'b01010101_11010111 : OUT <= 0;  //85 / 215 = 0
    16'b01010101_11011000 : OUT <= 0;  //85 / 216 = 0
    16'b01010101_11011001 : OUT <= 0;  //85 / 217 = 0
    16'b01010101_11011010 : OUT <= 0;  //85 / 218 = 0
    16'b01010101_11011011 : OUT <= 0;  //85 / 219 = 0
    16'b01010101_11011100 : OUT <= 0;  //85 / 220 = 0
    16'b01010101_11011101 : OUT <= 0;  //85 / 221 = 0
    16'b01010101_11011110 : OUT <= 0;  //85 / 222 = 0
    16'b01010101_11011111 : OUT <= 0;  //85 / 223 = 0
    16'b01010101_11100000 : OUT <= 0;  //85 / 224 = 0
    16'b01010101_11100001 : OUT <= 0;  //85 / 225 = 0
    16'b01010101_11100010 : OUT <= 0;  //85 / 226 = 0
    16'b01010101_11100011 : OUT <= 0;  //85 / 227 = 0
    16'b01010101_11100100 : OUT <= 0;  //85 / 228 = 0
    16'b01010101_11100101 : OUT <= 0;  //85 / 229 = 0
    16'b01010101_11100110 : OUT <= 0;  //85 / 230 = 0
    16'b01010101_11100111 : OUT <= 0;  //85 / 231 = 0
    16'b01010101_11101000 : OUT <= 0;  //85 / 232 = 0
    16'b01010101_11101001 : OUT <= 0;  //85 / 233 = 0
    16'b01010101_11101010 : OUT <= 0;  //85 / 234 = 0
    16'b01010101_11101011 : OUT <= 0;  //85 / 235 = 0
    16'b01010101_11101100 : OUT <= 0;  //85 / 236 = 0
    16'b01010101_11101101 : OUT <= 0;  //85 / 237 = 0
    16'b01010101_11101110 : OUT <= 0;  //85 / 238 = 0
    16'b01010101_11101111 : OUT <= 0;  //85 / 239 = 0
    16'b01010101_11110000 : OUT <= 0;  //85 / 240 = 0
    16'b01010101_11110001 : OUT <= 0;  //85 / 241 = 0
    16'b01010101_11110010 : OUT <= 0;  //85 / 242 = 0
    16'b01010101_11110011 : OUT <= 0;  //85 / 243 = 0
    16'b01010101_11110100 : OUT <= 0;  //85 / 244 = 0
    16'b01010101_11110101 : OUT <= 0;  //85 / 245 = 0
    16'b01010101_11110110 : OUT <= 0;  //85 / 246 = 0
    16'b01010101_11110111 : OUT <= 0;  //85 / 247 = 0
    16'b01010101_11111000 : OUT <= 0;  //85 / 248 = 0
    16'b01010101_11111001 : OUT <= 0;  //85 / 249 = 0
    16'b01010101_11111010 : OUT <= 0;  //85 / 250 = 0
    16'b01010101_11111011 : OUT <= 0;  //85 / 251 = 0
    16'b01010101_11111100 : OUT <= 0;  //85 / 252 = 0
    16'b01010101_11111101 : OUT <= 0;  //85 / 253 = 0
    16'b01010101_11111110 : OUT <= 0;  //85 / 254 = 0
    16'b01010101_11111111 : OUT <= 0;  //85 / 255 = 0
    16'b01010110_00000000 : OUT <= 0;  //86 / 0 = 0
    16'b01010110_00000001 : OUT <= 86;  //86 / 1 = 86
    16'b01010110_00000010 : OUT <= 43;  //86 / 2 = 43
    16'b01010110_00000011 : OUT <= 28;  //86 / 3 = 28
    16'b01010110_00000100 : OUT <= 21;  //86 / 4 = 21
    16'b01010110_00000101 : OUT <= 17;  //86 / 5 = 17
    16'b01010110_00000110 : OUT <= 14;  //86 / 6 = 14
    16'b01010110_00000111 : OUT <= 12;  //86 / 7 = 12
    16'b01010110_00001000 : OUT <= 10;  //86 / 8 = 10
    16'b01010110_00001001 : OUT <= 9;  //86 / 9 = 9
    16'b01010110_00001010 : OUT <= 8;  //86 / 10 = 8
    16'b01010110_00001011 : OUT <= 7;  //86 / 11 = 7
    16'b01010110_00001100 : OUT <= 7;  //86 / 12 = 7
    16'b01010110_00001101 : OUT <= 6;  //86 / 13 = 6
    16'b01010110_00001110 : OUT <= 6;  //86 / 14 = 6
    16'b01010110_00001111 : OUT <= 5;  //86 / 15 = 5
    16'b01010110_00010000 : OUT <= 5;  //86 / 16 = 5
    16'b01010110_00010001 : OUT <= 5;  //86 / 17 = 5
    16'b01010110_00010010 : OUT <= 4;  //86 / 18 = 4
    16'b01010110_00010011 : OUT <= 4;  //86 / 19 = 4
    16'b01010110_00010100 : OUT <= 4;  //86 / 20 = 4
    16'b01010110_00010101 : OUT <= 4;  //86 / 21 = 4
    16'b01010110_00010110 : OUT <= 3;  //86 / 22 = 3
    16'b01010110_00010111 : OUT <= 3;  //86 / 23 = 3
    16'b01010110_00011000 : OUT <= 3;  //86 / 24 = 3
    16'b01010110_00011001 : OUT <= 3;  //86 / 25 = 3
    16'b01010110_00011010 : OUT <= 3;  //86 / 26 = 3
    16'b01010110_00011011 : OUT <= 3;  //86 / 27 = 3
    16'b01010110_00011100 : OUT <= 3;  //86 / 28 = 3
    16'b01010110_00011101 : OUT <= 2;  //86 / 29 = 2
    16'b01010110_00011110 : OUT <= 2;  //86 / 30 = 2
    16'b01010110_00011111 : OUT <= 2;  //86 / 31 = 2
    16'b01010110_00100000 : OUT <= 2;  //86 / 32 = 2
    16'b01010110_00100001 : OUT <= 2;  //86 / 33 = 2
    16'b01010110_00100010 : OUT <= 2;  //86 / 34 = 2
    16'b01010110_00100011 : OUT <= 2;  //86 / 35 = 2
    16'b01010110_00100100 : OUT <= 2;  //86 / 36 = 2
    16'b01010110_00100101 : OUT <= 2;  //86 / 37 = 2
    16'b01010110_00100110 : OUT <= 2;  //86 / 38 = 2
    16'b01010110_00100111 : OUT <= 2;  //86 / 39 = 2
    16'b01010110_00101000 : OUT <= 2;  //86 / 40 = 2
    16'b01010110_00101001 : OUT <= 2;  //86 / 41 = 2
    16'b01010110_00101010 : OUT <= 2;  //86 / 42 = 2
    16'b01010110_00101011 : OUT <= 2;  //86 / 43 = 2
    16'b01010110_00101100 : OUT <= 1;  //86 / 44 = 1
    16'b01010110_00101101 : OUT <= 1;  //86 / 45 = 1
    16'b01010110_00101110 : OUT <= 1;  //86 / 46 = 1
    16'b01010110_00101111 : OUT <= 1;  //86 / 47 = 1
    16'b01010110_00110000 : OUT <= 1;  //86 / 48 = 1
    16'b01010110_00110001 : OUT <= 1;  //86 / 49 = 1
    16'b01010110_00110010 : OUT <= 1;  //86 / 50 = 1
    16'b01010110_00110011 : OUT <= 1;  //86 / 51 = 1
    16'b01010110_00110100 : OUT <= 1;  //86 / 52 = 1
    16'b01010110_00110101 : OUT <= 1;  //86 / 53 = 1
    16'b01010110_00110110 : OUT <= 1;  //86 / 54 = 1
    16'b01010110_00110111 : OUT <= 1;  //86 / 55 = 1
    16'b01010110_00111000 : OUT <= 1;  //86 / 56 = 1
    16'b01010110_00111001 : OUT <= 1;  //86 / 57 = 1
    16'b01010110_00111010 : OUT <= 1;  //86 / 58 = 1
    16'b01010110_00111011 : OUT <= 1;  //86 / 59 = 1
    16'b01010110_00111100 : OUT <= 1;  //86 / 60 = 1
    16'b01010110_00111101 : OUT <= 1;  //86 / 61 = 1
    16'b01010110_00111110 : OUT <= 1;  //86 / 62 = 1
    16'b01010110_00111111 : OUT <= 1;  //86 / 63 = 1
    16'b01010110_01000000 : OUT <= 1;  //86 / 64 = 1
    16'b01010110_01000001 : OUT <= 1;  //86 / 65 = 1
    16'b01010110_01000010 : OUT <= 1;  //86 / 66 = 1
    16'b01010110_01000011 : OUT <= 1;  //86 / 67 = 1
    16'b01010110_01000100 : OUT <= 1;  //86 / 68 = 1
    16'b01010110_01000101 : OUT <= 1;  //86 / 69 = 1
    16'b01010110_01000110 : OUT <= 1;  //86 / 70 = 1
    16'b01010110_01000111 : OUT <= 1;  //86 / 71 = 1
    16'b01010110_01001000 : OUT <= 1;  //86 / 72 = 1
    16'b01010110_01001001 : OUT <= 1;  //86 / 73 = 1
    16'b01010110_01001010 : OUT <= 1;  //86 / 74 = 1
    16'b01010110_01001011 : OUT <= 1;  //86 / 75 = 1
    16'b01010110_01001100 : OUT <= 1;  //86 / 76 = 1
    16'b01010110_01001101 : OUT <= 1;  //86 / 77 = 1
    16'b01010110_01001110 : OUT <= 1;  //86 / 78 = 1
    16'b01010110_01001111 : OUT <= 1;  //86 / 79 = 1
    16'b01010110_01010000 : OUT <= 1;  //86 / 80 = 1
    16'b01010110_01010001 : OUT <= 1;  //86 / 81 = 1
    16'b01010110_01010010 : OUT <= 1;  //86 / 82 = 1
    16'b01010110_01010011 : OUT <= 1;  //86 / 83 = 1
    16'b01010110_01010100 : OUT <= 1;  //86 / 84 = 1
    16'b01010110_01010101 : OUT <= 1;  //86 / 85 = 1
    16'b01010110_01010110 : OUT <= 1;  //86 / 86 = 1
    16'b01010110_01010111 : OUT <= 0;  //86 / 87 = 0
    16'b01010110_01011000 : OUT <= 0;  //86 / 88 = 0
    16'b01010110_01011001 : OUT <= 0;  //86 / 89 = 0
    16'b01010110_01011010 : OUT <= 0;  //86 / 90 = 0
    16'b01010110_01011011 : OUT <= 0;  //86 / 91 = 0
    16'b01010110_01011100 : OUT <= 0;  //86 / 92 = 0
    16'b01010110_01011101 : OUT <= 0;  //86 / 93 = 0
    16'b01010110_01011110 : OUT <= 0;  //86 / 94 = 0
    16'b01010110_01011111 : OUT <= 0;  //86 / 95 = 0
    16'b01010110_01100000 : OUT <= 0;  //86 / 96 = 0
    16'b01010110_01100001 : OUT <= 0;  //86 / 97 = 0
    16'b01010110_01100010 : OUT <= 0;  //86 / 98 = 0
    16'b01010110_01100011 : OUT <= 0;  //86 / 99 = 0
    16'b01010110_01100100 : OUT <= 0;  //86 / 100 = 0
    16'b01010110_01100101 : OUT <= 0;  //86 / 101 = 0
    16'b01010110_01100110 : OUT <= 0;  //86 / 102 = 0
    16'b01010110_01100111 : OUT <= 0;  //86 / 103 = 0
    16'b01010110_01101000 : OUT <= 0;  //86 / 104 = 0
    16'b01010110_01101001 : OUT <= 0;  //86 / 105 = 0
    16'b01010110_01101010 : OUT <= 0;  //86 / 106 = 0
    16'b01010110_01101011 : OUT <= 0;  //86 / 107 = 0
    16'b01010110_01101100 : OUT <= 0;  //86 / 108 = 0
    16'b01010110_01101101 : OUT <= 0;  //86 / 109 = 0
    16'b01010110_01101110 : OUT <= 0;  //86 / 110 = 0
    16'b01010110_01101111 : OUT <= 0;  //86 / 111 = 0
    16'b01010110_01110000 : OUT <= 0;  //86 / 112 = 0
    16'b01010110_01110001 : OUT <= 0;  //86 / 113 = 0
    16'b01010110_01110010 : OUT <= 0;  //86 / 114 = 0
    16'b01010110_01110011 : OUT <= 0;  //86 / 115 = 0
    16'b01010110_01110100 : OUT <= 0;  //86 / 116 = 0
    16'b01010110_01110101 : OUT <= 0;  //86 / 117 = 0
    16'b01010110_01110110 : OUT <= 0;  //86 / 118 = 0
    16'b01010110_01110111 : OUT <= 0;  //86 / 119 = 0
    16'b01010110_01111000 : OUT <= 0;  //86 / 120 = 0
    16'b01010110_01111001 : OUT <= 0;  //86 / 121 = 0
    16'b01010110_01111010 : OUT <= 0;  //86 / 122 = 0
    16'b01010110_01111011 : OUT <= 0;  //86 / 123 = 0
    16'b01010110_01111100 : OUT <= 0;  //86 / 124 = 0
    16'b01010110_01111101 : OUT <= 0;  //86 / 125 = 0
    16'b01010110_01111110 : OUT <= 0;  //86 / 126 = 0
    16'b01010110_01111111 : OUT <= 0;  //86 / 127 = 0
    16'b01010110_10000000 : OUT <= 0;  //86 / 128 = 0
    16'b01010110_10000001 : OUT <= 0;  //86 / 129 = 0
    16'b01010110_10000010 : OUT <= 0;  //86 / 130 = 0
    16'b01010110_10000011 : OUT <= 0;  //86 / 131 = 0
    16'b01010110_10000100 : OUT <= 0;  //86 / 132 = 0
    16'b01010110_10000101 : OUT <= 0;  //86 / 133 = 0
    16'b01010110_10000110 : OUT <= 0;  //86 / 134 = 0
    16'b01010110_10000111 : OUT <= 0;  //86 / 135 = 0
    16'b01010110_10001000 : OUT <= 0;  //86 / 136 = 0
    16'b01010110_10001001 : OUT <= 0;  //86 / 137 = 0
    16'b01010110_10001010 : OUT <= 0;  //86 / 138 = 0
    16'b01010110_10001011 : OUT <= 0;  //86 / 139 = 0
    16'b01010110_10001100 : OUT <= 0;  //86 / 140 = 0
    16'b01010110_10001101 : OUT <= 0;  //86 / 141 = 0
    16'b01010110_10001110 : OUT <= 0;  //86 / 142 = 0
    16'b01010110_10001111 : OUT <= 0;  //86 / 143 = 0
    16'b01010110_10010000 : OUT <= 0;  //86 / 144 = 0
    16'b01010110_10010001 : OUT <= 0;  //86 / 145 = 0
    16'b01010110_10010010 : OUT <= 0;  //86 / 146 = 0
    16'b01010110_10010011 : OUT <= 0;  //86 / 147 = 0
    16'b01010110_10010100 : OUT <= 0;  //86 / 148 = 0
    16'b01010110_10010101 : OUT <= 0;  //86 / 149 = 0
    16'b01010110_10010110 : OUT <= 0;  //86 / 150 = 0
    16'b01010110_10010111 : OUT <= 0;  //86 / 151 = 0
    16'b01010110_10011000 : OUT <= 0;  //86 / 152 = 0
    16'b01010110_10011001 : OUT <= 0;  //86 / 153 = 0
    16'b01010110_10011010 : OUT <= 0;  //86 / 154 = 0
    16'b01010110_10011011 : OUT <= 0;  //86 / 155 = 0
    16'b01010110_10011100 : OUT <= 0;  //86 / 156 = 0
    16'b01010110_10011101 : OUT <= 0;  //86 / 157 = 0
    16'b01010110_10011110 : OUT <= 0;  //86 / 158 = 0
    16'b01010110_10011111 : OUT <= 0;  //86 / 159 = 0
    16'b01010110_10100000 : OUT <= 0;  //86 / 160 = 0
    16'b01010110_10100001 : OUT <= 0;  //86 / 161 = 0
    16'b01010110_10100010 : OUT <= 0;  //86 / 162 = 0
    16'b01010110_10100011 : OUT <= 0;  //86 / 163 = 0
    16'b01010110_10100100 : OUT <= 0;  //86 / 164 = 0
    16'b01010110_10100101 : OUT <= 0;  //86 / 165 = 0
    16'b01010110_10100110 : OUT <= 0;  //86 / 166 = 0
    16'b01010110_10100111 : OUT <= 0;  //86 / 167 = 0
    16'b01010110_10101000 : OUT <= 0;  //86 / 168 = 0
    16'b01010110_10101001 : OUT <= 0;  //86 / 169 = 0
    16'b01010110_10101010 : OUT <= 0;  //86 / 170 = 0
    16'b01010110_10101011 : OUT <= 0;  //86 / 171 = 0
    16'b01010110_10101100 : OUT <= 0;  //86 / 172 = 0
    16'b01010110_10101101 : OUT <= 0;  //86 / 173 = 0
    16'b01010110_10101110 : OUT <= 0;  //86 / 174 = 0
    16'b01010110_10101111 : OUT <= 0;  //86 / 175 = 0
    16'b01010110_10110000 : OUT <= 0;  //86 / 176 = 0
    16'b01010110_10110001 : OUT <= 0;  //86 / 177 = 0
    16'b01010110_10110010 : OUT <= 0;  //86 / 178 = 0
    16'b01010110_10110011 : OUT <= 0;  //86 / 179 = 0
    16'b01010110_10110100 : OUT <= 0;  //86 / 180 = 0
    16'b01010110_10110101 : OUT <= 0;  //86 / 181 = 0
    16'b01010110_10110110 : OUT <= 0;  //86 / 182 = 0
    16'b01010110_10110111 : OUT <= 0;  //86 / 183 = 0
    16'b01010110_10111000 : OUT <= 0;  //86 / 184 = 0
    16'b01010110_10111001 : OUT <= 0;  //86 / 185 = 0
    16'b01010110_10111010 : OUT <= 0;  //86 / 186 = 0
    16'b01010110_10111011 : OUT <= 0;  //86 / 187 = 0
    16'b01010110_10111100 : OUT <= 0;  //86 / 188 = 0
    16'b01010110_10111101 : OUT <= 0;  //86 / 189 = 0
    16'b01010110_10111110 : OUT <= 0;  //86 / 190 = 0
    16'b01010110_10111111 : OUT <= 0;  //86 / 191 = 0
    16'b01010110_11000000 : OUT <= 0;  //86 / 192 = 0
    16'b01010110_11000001 : OUT <= 0;  //86 / 193 = 0
    16'b01010110_11000010 : OUT <= 0;  //86 / 194 = 0
    16'b01010110_11000011 : OUT <= 0;  //86 / 195 = 0
    16'b01010110_11000100 : OUT <= 0;  //86 / 196 = 0
    16'b01010110_11000101 : OUT <= 0;  //86 / 197 = 0
    16'b01010110_11000110 : OUT <= 0;  //86 / 198 = 0
    16'b01010110_11000111 : OUT <= 0;  //86 / 199 = 0
    16'b01010110_11001000 : OUT <= 0;  //86 / 200 = 0
    16'b01010110_11001001 : OUT <= 0;  //86 / 201 = 0
    16'b01010110_11001010 : OUT <= 0;  //86 / 202 = 0
    16'b01010110_11001011 : OUT <= 0;  //86 / 203 = 0
    16'b01010110_11001100 : OUT <= 0;  //86 / 204 = 0
    16'b01010110_11001101 : OUT <= 0;  //86 / 205 = 0
    16'b01010110_11001110 : OUT <= 0;  //86 / 206 = 0
    16'b01010110_11001111 : OUT <= 0;  //86 / 207 = 0
    16'b01010110_11010000 : OUT <= 0;  //86 / 208 = 0
    16'b01010110_11010001 : OUT <= 0;  //86 / 209 = 0
    16'b01010110_11010010 : OUT <= 0;  //86 / 210 = 0
    16'b01010110_11010011 : OUT <= 0;  //86 / 211 = 0
    16'b01010110_11010100 : OUT <= 0;  //86 / 212 = 0
    16'b01010110_11010101 : OUT <= 0;  //86 / 213 = 0
    16'b01010110_11010110 : OUT <= 0;  //86 / 214 = 0
    16'b01010110_11010111 : OUT <= 0;  //86 / 215 = 0
    16'b01010110_11011000 : OUT <= 0;  //86 / 216 = 0
    16'b01010110_11011001 : OUT <= 0;  //86 / 217 = 0
    16'b01010110_11011010 : OUT <= 0;  //86 / 218 = 0
    16'b01010110_11011011 : OUT <= 0;  //86 / 219 = 0
    16'b01010110_11011100 : OUT <= 0;  //86 / 220 = 0
    16'b01010110_11011101 : OUT <= 0;  //86 / 221 = 0
    16'b01010110_11011110 : OUT <= 0;  //86 / 222 = 0
    16'b01010110_11011111 : OUT <= 0;  //86 / 223 = 0
    16'b01010110_11100000 : OUT <= 0;  //86 / 224 = 0
    16'b01010110_11100001 : OUT <= 0;  //86 / 225 = 0
    16'b01010110_11100010 : OUT <= 0;  //86 / 226 = 0
    16'b01010110_11100011 : OUT <= 0;  //86 / 227 = 0
    16'b01010110_11100100 : OUT <= 0;  //86 / 228 = 0
    16'b01010110_11100101 : OUT <= 0;  //86 / 229 = 0
    16'b01010110_11100110 : OUT <= 0;  //86 / 230 = 0
    16'b01010110_11100111 : OUT <= 0;  //86 / 231 = 0
    16'b01010110_11101000 : OUT <= 0;  //86 / 232 = 0
    16'b01010110_11101001 : OUT <= 0;  //86 / 233 = 0
    16'b01010110_11101010 : OUT <= 0;  //86 / 234 = 0
    16'b01010110_11101011 : OUT <= 0;  //86 / 235 = 0
    16'b01010110_11101100 : OUT <= 0;  //86 / 236 = 0
    16'b01010110_11101101 : OUT <= 0;  //86 / 237 = 0
    16'b01010110_11101110 : OUT <= 0;  //86 / 238 = 0
    16'b01010110_11101111 : OUT <= 0;  //86 / 239 = 0
    16'b01010110_11110000 : OUT <= 0;  //86 / 240 = 0
    16'b01010110_11110001 : OUT <= 0;  //86 / 241 = 0
    16'b01010110_11110010 : OUT <= 0;  //86 / 242 = 0
    16'b01010110_11110011 : OUT <= 0;  //86 / 243 = 0
    16'b01010110_11110100 : OUT <= 0;  //86 / 244 = 0
    16'b01010110_11110101 : OUT <= 0;  //86 / 245 = 0
    16'b01010110_11110110 : OUT <= 0;  //86 / 246 = 0
    16'b01010110_11110111 : OUT <= 0;  //86 / 247 = 0
    16'b01010110_11111000 : OUT <= 0;  //86 / 248 = 0
    16'b01010110_11111001 : OUT <= 0;  //86 / 249 = 0
    16'b01010110_11111010 : OUT <= 0;  //86 / 250 = 0
    16'b01010110_11111011 : OUT <= 0;  //86 / 251 = 0
    16'b01010110_11111100 : OUT <= 0;  //86 / 252 = 0
    16'b01010110_11111101 : OUT <= 0;  //86 / 253 = 0
    16'b01010110_11111110 : OUT <= 0;  //86 / 254 = 0
    16'b01010110_11111111 : OUT <= 0;  //86 / 255 = 0
    16'b01010111_00000000 : OUT <= 0;  //87 / 0 = 0
    16'b01010111_00000001 : OUT <= 87;  //87 / 1 = 87
    16'b01010111_00000010 : OUT <= 43;  //87 / 2 = 43
    16'b01010111_00000011 : OUT <= 29;  //87 / 3 = 29
    16'b01010111_00000100 : OUT <= 21;  //87 / 4 = 21
    16'b01010111_00000101 : OUT <= 17;  //87 / 5 = 17
    16'b01010111_00000110 : OUT <= 14;  //87 / 6 = 14
    16'b01010111_00000111 : OUT <= 12;  //87 / 7 = 12
    16'b01010111_00001000 : OUT <= 10;  //87 / 8 = 10
    16'b01010111_00001001 : OUT <= 9;  //87 / 9 = 9
    16'b01010111_00001010 : OUT <= 8;  //87 / 10 = 8
    16'b01010111_00001011 : OUT <= 7;  //87 / 11 = 7
    16'b01010111_00001100 : OUT <= 7;  //87 / 12 = 7
    16'b01010111_00001101 : OUT <= 6;  //87 / 13 = 6
    16'b01010111_00001110 : OUT <= 6;  //87 / 14 = 6
    16'b01010111_00001111 : OUT <= 5;  //87 / 15 = 5
    16'b01010111_00010000 : OUT <= 5;  //87 / 16 = 5
    16'b01010111_00010001 : OUT <= 5;  //87 / 17 = 5
    16'b01010111_00010010 : OUT <= 4;  //87 / 18 = 4
    16'b01010111_00010011 : OUT <= 4;  //87 / 19 = 4
    16'b01010111_00010100 : OUT <= 4;  //87 / 20 = 4
    16'b01010111_00010101 : OUT <= 4;  //87 / 21 = 4
    16'b01010111_00010110 : OUT <= 3;  //87 / 22 = 3
    16'b01010111_00010111 : OUT <= 3;  //87 / 23 = 3
    16'b01010111_00011000 : OUT <= 3;  //87 / 24 = 3
    16'b01010111_00011001 : OUT <= 3;  //87 / 25 = 3
    16'b01010111_00011010 : OUT <= 3;  //87 / 26 = 3
    16'b01010111_00011011 : OUT <= 3;  //87 / 27 = 3
    16'b01010111_00011100 : OUT <= 3;  //87 / 28 = 3
    16'b01010111_00011101 : OUT <= 3;  //87 / 29 = 3
    16'b01010111_00011110 : OUT <= 2;  //87 / 30 = 2
    16'b01010111_00011111 : OUT <= 2;  //87 / 31 = 2
    16'b01010111_00100000 : OUT <= 2;  //87 / 32 = 2
    16'b01010111_00100001 : OUT <= 2;  //87 / 33 = 2
    16'b01010111_00100010 : OUT <= 2;  //87 / 34 = 2
    16'b01010111_00100011 : OUT <= 2;  //87 / 35 = 2
    16'b01010111_00100100 : OUT <= 2;  //87 / 36 = 2
    16'b01010111_00100101 : OUT <= 2;  //87 / 37 = 2
    16'b01010111_00100110 : OUT <= 2;  //87 / 38 = 2
    16'b01010111_00100111 : OUT <= 2;  //87 / 39 = 2
    16'b01010111_00101000 : OUT <= 2;  //87 / 40 = 2
    16'b01010111_00101001 : OUT <= 2;  //87 / 41 = 2
    16'b01010111_00101010 : OUT <= 2;  //87 / 42 = 2
    16'b01010111_00101011 : OUT <= 2;  //87 / 43 = 2
    16'b01010111_00101100 : OUT <= 1;  //87 / 44 = 1
    16'b01010111_00101101 : OUT <= 1;  //87 / 45 = 1
    16'b01010111_00101110 : OUT <= 1;  //87 / 46 = 1
    16'b01010111_00101111 : OUT <= 1;  //87 / 47 = 1
    16'b01010111_00110000 : OUT <= 1;  //87 / 48 = 1
    16'b01010111_00110001 : OUT <= 1;  //87 / 49 = 1
    16'b01010111_00110010 : OUT <= 1;  //87 / 50 = 1
    16'b01010111_00110011 : OUT <= 1;  //87 / 51 = 1
    16'b01010111_00110100 : OUT <= 1;  //87 / 52 = 1
    16'b01010111_00110101 : OUT <= 1;  //87 / 53 = 1
    16'b01010111_00110110 : OUT <= 1;  //87 / 54 = 1
    16'b01010111_00110111 : OUT <= 1;  //87 / 55 = 1
    16'b01010111_00111000 : OUT <= 1;  //87 / 56 = 1
    16'b01010111_00111001 : OUT <= 1;  //87 / 57 = 1
    16'b01010111_00111010 : OUT <= 1;  //87 / 58 = 1
    16'b01010111_00111011 : OUT <= 1;  //87 / 59 = 1
    16'b01010111_00111100 : OUT <= 1;  //87 / 60 = 1
    16'b01010111_00111101 : OUT <= 1;  //87 / 61 = 1
    16'b01010111_00111110 : OUT <= 1;  //87 / 62 = 1
    16'b01010111_00111111 : OUT <= 1;  //87 / 63 = 1
    16'b01010111_01000000 : OUT <= 1;  //87 / 64 = 1
    16'b01010111_01000001 : OUT <= 1;  //87 / 65 = 1
    16'b01010111_01000010 : OUT <= 1;  //87 / 66 = 1
    16'b01010111_01000011 : OUT <= 1;  //87 / 67 = 1
    16'b01010111_01000100 : OUT <= 1;  //87 / 68 = 1
    16'b01010111_01000101 : OUT <= 1;  //87 / 69 = 1
    16'b01010111_01000110 : OUT <= 1;  //87 / 70 = 1
    16'b01010111_01000111 : OUT <= 1;  //87 / 71 = 1
    16'b01010111_01001000 : OUT <= 1;  //87 / 72 = 1
    16'b01010111_01001001 : OUT <= 1;  //87 / 73 = 1
    16'b01010111_01001010 : OUT <= 1;  //87 / 74 = 1
    16'b01010111_01001011 : OUT <= 1;  //87 / 75 = 1
    16'b01010111_01001100 : OUT <= 1;  //87 / 76 = 1
    16'b01010111_01001101 : OUT <= 1;  //87 / 77 = 1
    16'b01010111_01001110 : OUT <= 1;  //87 / 78 = 1
    16'b01010111_01001111 : OUT <= 1;  //87 / 79 = 1
    16'b01010111_01010000 : OUT <= 1;  //87 / 80 = 1
    16'b01010111_01010001 : OUT <= 1;  //87 / 81 = 1
    16'b01010111_01010010 : OUT <= 1;  //87 / 82 = 1
    16'b01010111_01010011 : OUT <= 1;  //87 / 83 = 1
    16'b01010111_01010100 : OUT <= 1;  //87 / 84 = 1
    16'b01010111_01010101 : OUT <= 1;  //87 / 85 = 1
    16'b01010111_01010110 : OUT <= 1;  //87 / 86 = 1
    16'b01010111_01010111 : OUT <= 1;  //87 / 87 = 1
    16'b01010111_01011000 : OUT <= 0;  //87 / 88 = 0
    16'b01010111_01011001 : OUT <= 0;  //87 / 89 = 0
    16'b01010111_01011010 : OUT <= 0;  //87 / 90 = 0
    16'b01010111_01011011 : OUT <= 0;  //87 / 91 = 0
    16'b01010111_01011100 : OUT <= 0;  //87 / 92 = 0
    16'b01010111_01011101 : OUT <= 0;  //87 / 93 = 0
    16'b01010111_01011110 : OUT <= 0;  //87 / 94 = 0
    16'b01010111_01011111 : OUT <= 0;  //87 / 95 = 0
    16'b01010111_01100000 : OUT <= 0;  //87 / 96 = 0
    16'b01010111_01100001 : OUT <= 0;  //87 / 97 = 0
    16'b01010111_01100010 : OUT <= 0;  //87 / 98 = 0
    16'b01010111_01100011 : OUT <= 0;  //87 / 99 = 0
    16'b01010111_01100100 : OUT <= 0;  //87 / 100 = 0
    16'b01010111_01100101 : OUT <= 0;  //87 / 101 = 0
    16'b01010111_01100110 : OUT <= 0;  //87 / 102 = 0
    16'b01010111_01100111 : OUT <= 0;  //87 / 103 = 0
    16'b01010111_01101000 : OUT <= 0;  //87 / 104 = 0
    16'b01010111_01101001 : OUT <= 0;  //87 / 105 = 0
    16'b01010111_01101010 : OUT <= 0;  //87 / 106 = 0
    16'b01010111_01101011 : OUT <= 0;  //87 / 107 = 0
    16'b01010111_01101100 : OUT <= 0;  //87 / 108 = 0
    16'b01010111_01101101 : OUT <= 0;  //87 / 109 = 0
    16'b01010111_01101110 : OUT <= 0;  //87 / 110 = 0
    16'b01010111_01101111 : OUT <= 0;  //87 / 111 = 0
    16'b01010111_01110000 : OUT <= 0;  //87 / 112 = 0
    16'b01010111_01110001 : OUT <= 0;  //87 / 113 = 0
    16'b01010111_01110010 : OUT <= 0;  //87 / 114 = 0
    16'b01010111_01110011 : OUT <= 0;  //87 / 115 = 0
    16'b01010111_01110100 : OUT <= 0;  //87 / 116 = 0
    16'b01010111_01110101 : OUT <= 0;  //87 / 117 = 0
    16'b01010111_01110110 : OUT <= 0;  //87 / 118 = 0
    16'b01010111_01110111 : OUT <= 0;  //87 / 119 = 0
    16'b01010111_01111000 : OUT <= 0;  //87 / 120 = 0
    16'b01010111_01111001 : OUT <= 0;  //87 / 121 = 0
    16'b01010111_01111010 : OUT <= 0;  //87 / 122 = 0
    16'b01010111_01111011 : OUT <= 0;  //87 / 123 = 0
    16'b01010111_01111100 : OUT <= 0;  //87 / 124 = 0
    16'b01010111_01111101 : OUT <= 0;  //87 / 125 = 0
    16'b01010111_01111110 : OUT <= 0;  //87 / 126 = 0
    16'b01010111_01111111 : OUT <= 0;  //87 / 127 = 0
    16'b01010111_10000000 : OUT <= 0;  //87 / 128 = 0
    16'b01010111_10000001 : OUT <= 0;  //87 / 129 = 0
    16'b01010111_10000010 : OUT <= 0;  //87 / 130 = 0
    16'b01010111_10000011 : OUT <= 0;  //87 / 131 = 0
    16'b01010111_10000100 : OUT <= 0;  //87 / 132 = 0
    16'b01010111_10000101 : OUT <= 0;  //87 / 133 = 0
    16'b01010111_10000110 : OUT <= 0;  //87 / 134 = 0
    16'b01010111_10000111 : OUT <= 0;  //87 / 135 = 0
    16'b01010111_10001000 : OUT <= 0;  //87 / 136 = 0
    16'b01010111_10001001 : OUT <= 0;  //87 / 137 = 0
    16'b01010111_10001010 : OUT <= 0;  //87 / 138 = 0
    16'b01010111_10001011 : OUT <= 0;  //87 / 139 = 0
    16'b01010111_10001100 : OUT <= 0;  //87 / 140 = 0
    16'b01010111_10001101 : OUT <= 0;  //87 / 141 = 0
    16'b01010111_10001110 : OUT <= 0;  //87 / 142 = 0
    16'b01010111_10001111 : OUT <= 0;  //87 / 143 = 0
    16'b01010111_10010000 : OUT <= 0;  //87 / 144 = 0
    16'b01010111_10010001 : OUT <= 0;  //87 / 145 = 0
    16'b01010111_10010010 : OUT <= 0;  //87 / 146 = 0
    16'b01010111_10010011 : OUT <= 0;  //87 / 147 = 0
    16'b01010111_10010100 : OUT <= 0;  //87 / 148 = 0
    16'b01010111_10010101 : OUT <= 0;  //87 / 149 = 0
    16'b01010111_10010110 : OUT <= 0;  //87 / 150 = 0
    16'b01010111_10010111 : OUT <= 0;  //87 / 151 = 0
    16'b01010111_10011000 : OUT <= 0;  //87 / 152 = 0
    16'b01010111_10011001 : OUT <= 0;  //87 / 153 = 0
    16'b01010111_10011010 : OUT <= 0;  //87 / 154 = 0
    16'b01010111_10011011 : OUT <= 0;  //87 / 155 = 0
    16'b01010111_10011100 : OUT <= 0;  //87 / 156 = 0
    16'b01010111_10011101 : OUT <= 0;  //87 / 157 = 0
    16'b01010111_10011110 : OUT <= 0;  //87 / 158 = 0
    16'b01010111_10011111 : OUT <= 0;  //87 / 159 = 0
    16'b01010111_10100000 : OUT <= 0;  //87 / 160 = 0
    16'b01010111_10100001 : OUT <= 0;  //87 / 161 = 0
    16'b01010111_10100010 : OUT <= 0;  //87 / 162 = 0
    16'b01010111_10100011 : OUT <= 0;  //87 / 163 = 0
    16'b01010111_10100100 : OUT <= 0;  //87 / 164 = 0
    16'b01010111_10100101 : OUT <= 0;  //87 / 165 = 0
    16'b01010111_10100110 : OUT <= 0;  //87 / 166 = 0
    16'b01010111_10100111 : OUT <= 0;  //87 / 167 = 0
    16'b01010111_10101000 : OUT <= 0;  //87 / 168 = 0
    16'b01010111_10101001 : OUT <= 0;  //87 / 169 = 0
    16'b01010111_10101010 : OUT <= 0;  //87 / 170 = 0
    16'b01010111_10101011 : OUT <= 0;  //87 / 171 = 0
    16'b01010111_10101100 : OUT <= 0;  //87 / 172 = 0
    16'b01010111_10101101 : OUT <= 0;  //87 / 173 = 0
    16'b01010111_10101110 : OUT <= 0;  //87 / 174 = 0
    16'b01010111_10101111 : OUT <= 0;  //87 / 175 = 0
    16'b01010111_10110000 : OUT <= 0;  //87 / 176 = 0
    16'b01010111_10110001 : OUT <= 0;  //87 / 177 = 0
    16'b01010111_10110010 : OUT <= 0;  //87 / 178 = 0
    16'b01010111_10110011 : OUT <= 0;  //87 / 179 = 0
    16'b01010111_10110100 : OUT <= 0;  //87 / 180 = 0
    16'b01010111_10110101 : OUT <= 0;  //87 / 181 = 0
    16'b01010111_10110110 : OUT <= 0;  //87 / 182 = 0
    16'b01010111_10110111 : OUT <= 0;  //87 / 183 = 0
    16'b01010111_10111000 : OUT <= 0;  //87 / 184 = 0
    16'b01010111_10111001 : OUT <= 0;  //87 / 185 = 0
    16'b01010111_10111010 : OUT <= 0;  //87 / 186 = 0
    16'b01010111_10111011 : OUT <= 0;  //87 / 187 = 0
    16'b01010111_10111100 : OUT <= 0;  //87 / 188 = 0
    16'b01010111_10111101 : OUT <= 0;  //87 / 189 = 0
    16'b01010111_10111110 : OUT <= 0;  //87 / 190 = 0
    16'b01010111_10111111 : OUT <= 0;  //87 / 191 = 0
    16'b01010111_11000000 : OUT <= 0;  //87 / 192 = 0
    16'b01010111_11000001 : OUT <= 0;  //87 / 193 = 0
    16'b01010111_11000010 : OUT <= 0;  //87 / 194 = 0
    16'b01010111_11000011 : OUT <= 0;  //87 / 195 = 0
    16'b01010111_11000100 : OUT <= 0;  //87 / 196 = 0
    16'b01010111_11000101 : OUT <= 0;  //87 / 197 = 0
    16'b01010111_11000110 : OUT <= 0;  //87 / 198 = 0
    16'b01010111_11000111 : OUT <= 0;  //87 / 199 = 0
    16'b01010111_11001000 : OUT <= 0;  //87 / 200 = 0
    16'b01010111_11001001 : OUT <= 0;  //87 / 201 = 0
    16'b01010111_11001010 : OUT <= 0;  //87 / 202 = 0
    16'b01010111_11001011 : OUT <= 0;  //87 / 203 = 0
    16'b01010111_11001100 : OUT <= 0;  //87 / 204 = 0
    16'b01010111_11001101 : OUT <= 0;  //87 / 205 = 0
    16'b01010111_11001110 : OUT <= 0;  //87 / 206 = 0
    16'b01010111_11001111 : OUT <= 0;  //87 / 207 = 0
    16'b01010111_11010000 : OUT <= 0;  //87 / 208 = 0
    16'b01010111_11010001 : OUT <= 0;  //87 / 209 = 0
    16'b01010111_11010010 : OUT <= 0;  //87 / 210 = 0
    16'b01010111_11010011 : OUT <= 0;  //87 / 211 = 0
    16'b01010111_11010100 : OUT <= 0;  //87 / 212 = 0
    16'b01010111_11010101 : OUT <= 0;  //87 / 213 = 0
    16'b01010111_11010110 : OUT <= 0;  //87 / 214 = 0
    16'b01010111_11010111 : OUT <= 0;  //87 / 215 = 0
    16'b01010111_11011000 : OUT <= 0;  //87 / 216 = 0
    16'b01010111_11011001 : OUT <= 0;  //87 / 217 = 0
    16'b01010111_11011010 : OUT <= 0;  //87 / 218 = 0
    16'b01010111_11011011 : OUT <= 0;  //87 / 219 = 0
    16'b01010111_11011100 : OUT <= 0;  //87 / 220 = 0
    16'b01010111_11011101 : OUT <= 0;  //87 / 221 = 0
    16'b01010111_11011110 : OUT <= 0;  //87 / 222 = 0
    16'b01010111_11011111 : OUT <= 0;  //87 / 223 = 0
    16'b01010111_11100000 : OUT <= 0;  //87 / 224 = 0
    16'b01010111_11100001 : OUT <= 0;  //87 / 225 = 0
    16'b01010111_11100010 : OUT <= 0;  //87 / 226 = 0
    16'b01010111_11100011 : OUT <= 0;  //87 / 227 = 0
    16'b01010111_11100100 : OUT <= 0;  //87 / 228 = 0
    16'b01010111_11100101 : OUT <= 0;  //87 / 229 = 0
    16'b01010111_11100110 : OUT <= 0;  //87 / 230 = 0
    16'b01010111_11100111 : OUT <= 0;  //87 / 231 = 0
    16'b01010111_11101000 : OUT <= 0;  //87 / 232 = 0
    16'b01010111_11101001 : OUT <= 0;  //87 / 233 = 0
    16'b01010111_11101010 : OUT <= 0;  //87 / 234 = 0
    16'b01010111_11101011 : OUT <= 0;  //87 / 235 = 0
    16'b01010111_11101100 : OUT <= 0;  //87 / 236 = 0
    16'b01010111_11101101 : OUT <= 0;  //87 / 237 = 0
    16'b01010111_11101110 : OUT <= 0;  //87 / 238 = 0
    16'b01010111_11101111 : OUT <= 0;  //87 / 239 = 0
    16'b01010111_11110000 : OUT <= 0;  //87 / 240 = 0
    16'b01010111_11110001 : OUT <= 0;  //87 / 241 = 0
    16'b01010111_11110010 : OUT <= 0;  //87 / 242 = 0
    16'b01010111_11110011 : OUT <= 0;  //87 / 243 = 0
    16'b01010111_11110100 : OUT <= 0;  //87 / 244 = 0
    16'b01010111_11110101 : OUT <= 0;  //87 / 245 = 0
    16'b01010111_11110110 : OUT <= 0;  //87 / 246 = 0
    16'b01010111_11110111 : OUT <= 0;  //87 / 247 = 0
    16'b01010111_11111000 : OUT <= 0;  //87 / 248 = 0
    16'b01010111_11111001 : OUT <= 0;  //87 / 249 = 0
    16'b01010111_11111010 : OUT <= 0;  //87 / 250 = 0
    16'b01010111_11111011 : OUT <= 0;  //87 / 251 = 0
    16'b01010111_11111100 : OUT <= 0;  //87 / 252 = 0
    16'b01010111_11111101 : OUT <= 0;  //87 / 253 = 0
    16'b01010111_11111110 : OUT <= 0;  //87 / 254 = 0
    16'b01010111_11111111 : OUT <= 0;  //87 / 255 = 0
    16'b01011000_00000000 : OUT <= 0;  //88 / 0 = 0
    16'b01011000_00000001 : OUT <= 88;  //88 / 1 = 88
    16'b01011000_00000010 : OUT <= 44;  //88 / 2 = 44
    16'b01011000_00000011 : OUT <= 29;  //88 / 3 = 29
    16'b01011000_00000100 : OUT <= 22;  //88 / 4 = 22
    16'b01011000_00000101 : OUT <= 17;  //88 / 5 = 17
    16'b01011000_00000110 : OUT <= 14;  //88 / 6 = 14
    16'b01011000_00000111 : OUT <= 12;  //88 / 7 = 12
    16'b01011000_00001000 : OUT <= 11;  //88 / 8 = 11
    16'b01011000_00001001 : OUT <= 9;  //88 / 9 = 9
    16'b01011000_00001010 : OUT <= 8;  //88 / 10 = 8
    16'b01011000_00001011 : OUT <= 8;  //88 / 11 = 8
    16'b01011000_00001100 : OUT <= 7;  //88 / 12 = 7
    16'b01011000_00001101 : OUT <= 6;  //88 / 13 = 6
    16'b01011000_00001110 : OUT <= 6;  //88 / 14 = 6
    16'b01011000_00001111 : OUT <= 5;  //88 / 15 = 5
    16'b01011000_00010000 : OUT <= 5;  //88 / 16 = 5
    16'b01011000_00010001 : OUT <= 5;  //88 / 17 = 5
    16'b01011000_00010010 : OUT <= 4;  //88 / 18 = 4
    16'b01011000_00010011 : OUT <= 4;  //88 / 19 = 4
    16'b01011000_00010100 : OUT <= 4;  //88 / 20 = 4
    16'b01011000_00010101 : OUT <= 4;  //88 / 21 = 4
    16'b01011000_00010110 : OUT <= 4;  //88 / 22 = 4
    16'b01011000_00010111 : OUT <= 3;  //88 / 23 = 3
    16'b01011000_00011000 : OUT <= 3;  //88 / 24 = 3
    16'b01011000_00011001 : OUT <= 3;  //88 / 25 = 3
    16'b01011000_00011010 : OUT <= 3;  //88 / 26 = 3
    16'b01011000_00011011 : OUT <= 3;  //88 / 27 = 3
    16'b01011000_00011100 : OUT <= 3;  //88 / 28 = 3
    16'b01011000_00011101 : OUT <= 3;  //88 / 29 = 3
    16'b01011000_00011110 : OUT <= 2;  //88 / 30 = 2
    16'b01011000_00011111 : OUT <= 2;  //88 / 31 = 2
    16'b01011000_00100000 : OUT <= 2;  //88 / 32 = 2
    16'b01011000_00100001 : OUT <= 2;  //88 / 33 = 2
    16'b01011000_00100010 : OUT <= 2;  //88 / 34 = 2
    16'b01011000_00100011 : OUT <= 2;  //88 / 35 = 2
    16'b01011000_00100100 : OUT <= 2;  //88 / 36 = 2
    16'b01011000_00100101 : OUT <= 2;  //88 / 37 = 2
    16'b01011000_00100110 : OUT <= 2;  //88 / 38 = 2
    16'b01011000_00100111 : OUT <= 2;  //88 / 39 = 2
    16'b01011000_00101000 : OUT <= 2;  //88 / 40 = 2
    16'b01011000_00101001 : OUT <= 2;  //88 / 41 = 2
    16'b01011000_00101010 : OUT <= 2;  //88 / 42 = 2
    16'b01011000_00101011 : OUT <= 2;  //88 / 43 = 2
    16'b01011000_00101100 : OUT <= 2;  //88 / 44 = 2
    16'b01011000_00101101 : OUT <= 1;  //88 / 45 = 1
    16'b01011000_00101110 : OUT <= 1;  //88 / 46 = 1
    16'b01011000_00101111 : OUT <= 1;  //88 / 47 = 1
    16'b01011000_00110000 : OUT <= 1;  //88 / 48 = 1
    16'b01011000_00110001 : OUT <= 1;  //88 / 49 = 1
    16'b01011000_00110010 : OUT <= 1;  //88 / 50 = 1
    16'b01011000_00110011 : OUT <= 1;  //88 / 51 = 1
    16'b01011000_00110100 : OUT <= 1;  //88 / 52 = 1
    16'b01011000_00110101 : OUT <= 1;  //88 / 53 = 1
    16'b01011000_00110110 : OUT <= 1;  //88 / 54 = 1
    16'b01011000_00110111 : OUT <= 1;  //88 / 55 = 1
    16'b01011000_00111000 : OUT <= 1;  //88 / 56 = 1
    16'b01011000_00111001 : OUT <= 1;  //88 / 57 = 1
    16'b01011000_00111010 : OUT <= 1;  //88 / 58 = 1
    16'b01011000_00111011 : OUT <= 1;  //88 / 59 = 1
    16'b01011000_00111100 : OUT <= 1;  //88 / 60 = 1
    16'b01011000_00111101 : OUT <= 1;  //88 / 61 = 1
    16'b01011000_00111110 : OUT <= 1;  //88 / 62 = 1
    16'b01011000_00111111 : OUT <= 1;  //88 / 63 = 1
    16'b01011000_01000000 : OUT <= 1;  //88 / 64 = 1
    16'b01011000_01000001 : OUT <= 1;  //88 / 65 = 1
    16'b01011000_01000010 : OUT <= 1;  //88 / 66 = 1
    16'b01011000_01000011 : OUT <= 1;  //88 / 67 = 1
    16'b01011000_01000100 : OUT <= 1;  //88 / 68 = 1
    16'b01011000_01000101 : OUT <= 1;  //88 / 69 = 1
    16'b01011000_01000110 : OUT <= 1;  //88 / 70 = 1
    16'b01011000_01000111 : OUT <= 1;  //88 / 71 = 1
    16'b01011000_01001000 : OUT <= 1;  //88 / 72 = 1
    16'b01011000_01001001 : OUT <= 1;  //88 / 73 = 1
    16'b01011000_01001010 : OUT <= 1;  //88 / 74 = 1
    16'b01011000_01001011 : OUT <= 1;  //88 / 75 = 1
    16'b01011000_01001100 : OUT <= 1;  //88 / 76 = 1
    16'b01011000_01001101 : OUT <= 1;  //88 / 77 = 1
    16'b01011000_01001110 : OUT <= 1;  //88 / 78 = 1
    16'b01011000_01001111 : OUT <= 1;  //88 / 79 = 1
    16'b01011000_01010000 : OUT <= 1;  //88 / 80 = 1
    16'b01011000_01010001 : OUT <= 1;  //88 / 81 = 1
    16'b01011000_01010010 : OUT <= 1;  //88 / 82 = 1
    16'b01011000_01010011 : OUT <= 1;  //88 / 83 = 1
    16'b01011000_01010100 : OUT <= 1;  //88 / 84 = 1
    16'b01011000_01010101 : OUT <= 1;  //88 / 85 = 1
    16'b01011000_01010110 : OUT <= 1;  //88 / 86 = 1
    16'b01011000_01010111 : OUT <= 1;  //88 / 87 = 1
    16'b01011000_01011000 : OUT <= 1;  //88 / 88 = 1
    16'b01011000_01011001 : OUT <= 0;  //88 / 89 = 0
    16'b01011000_01011010 : OUT <= 0;  //88 / 90 = 0
    16'b01011000_01011011 : OUT <= 0;  //88 / 91 = 0
    16'b01011000_01011100 : OUT <= 0;  //88 / 92 = 0
    16'b01011000_01011101 : OUT <= 0;  //88 / 93 = 0
    16'b01011000_01011110 : OUT <= 0;  //88 / 94 = 0
    16'b01011000_01011111 : OUT <= 0;  //88 / 95 = 0
    16'b01011000_01100000 : OUT <= 0;  //88 / 96 = 0
    16'b01011000_01100001 : OUT <= 0;  //88 / 97 = 0
    16'b01011000_01100010 : OUT <= 0;  //88 / 98 = 0
    16'b01011000_01100011 : OUT <= 0;  //88 / 99 = 0
    16'b01011000_01100100 : OUT <= 0;  //88 / 100 = 0
    16'b01011000_01100101 : OUT <= 0;  //88 / 101 = 0
    16'b01011000_01100110 : OUT <= 0;  //88 / 102 = 0
    16'b01011000_01100111 : OUT <= 0;  //88 / 103 = 0
    16'b01011000_01101000 : OUT <= 0;  //88 / 104 = 0
    16'b01011000_01101001 : OUT <= 0;  //88 / 105 = 0
    16'b01011000_01101010 : OUT <= 0;  //88 / 106 = 0
    16'b01011000_01101011 : OUT <= 0;  //88 / 107 = 0
    16'b01011000_01101100 : OUT <= 0;  //88 / 108 = 0
    16'b01011000_01101101 : OUT <= 0;  //88 / 109 = 0
    16'b01011000_01101110 : OUT <= 0;  //88 / 110 = 0
    16'b01011000_01101111 : OUT <= 0;  //88 / 111 = 0
    16'b01011000_01110000 : OUT <= 0;  //88 / 112 = 0
    16'b01011000_01110001 : OUT <= 0;  //88 / 113 = 0
    16'b01011000_01110010 : OUT <= 0;  //88 / 114 = 0
    16'b01011000_01110011 : OUT <= 0;  //88 / 115 = 0
    16'b01011000_01110100 : OUT <= 0;  //88 / 116 = 0
    16'b01011000_01110101 : OUT <= 0;  //88 / 117 = 0
    16'b01011000_01110110 : OUT <= 0;  //88 / 118 = 0
    16'b01011000_01110111 : OUT <= 0;  //88 / 119 = 0
    16'b01011000_01111000 : OUT <= 0;  //88 / 120 = 0
    16'b01011000_01111001 : OUT <= 0;  //88 / 121 = 0
    16'b01011000_01111010 : OUT <= 0;  //88 / 122 = 0
    16'b01011000_01111011 : OUT <= 0;  //88 / 123 = 0
    16'b01011000_01111100 : OUT <= 0;  //88 / 124 = 0
    16'b01011000_01111101 : OUT <= 0;  //88 / 125 = 0
    16'b01011000_01111110 : OUT <= 0;  //88 / 126 = 0
    16'b01011000_01111111 : OUT <= 0;  //88 / 127 = 0
    16'b01011000_10000000 : OUT <= 0;  //88 / 128 = 0
    16'b01011000_10000001 : OUT <= 0;  //88 / 129 = 0
    16'b01011000_10000010 : OUT <= 0;  //88 / 130 = 0
    16'b01011000_10000011 : OUT <= 0;  //88 / 131 = 0
    16'b01011000_10000100 : OUT <= 0;  //88 / 132 = 0
    16'b01011000_10000101 : OUT <= 0;  //88 / 133 = 0
    16'b01011000_10000110 : OUT <= 0;  //88 / 134 = 0
    16'b01011000_10000111 : OUT <= 0;  //88 / 135 = 0
    16'b01011000_10001000 : OUT <= 0;  //88 / 136 = 0
    16'b01011000_10001001 : OUT <= 0;  //88 / 137 = 0
    16'b01011000_10001010 : OUT <= 0;  //88 / 138 = 0
    16'b01011000_10001011 : OUT <= 0;  //88 / 139 = 0
    16'b01011000_10001100 : OUT <= 0;  //88 / 140 = 0
    16'b01011000_10001101 : OUT <= 0;  //88 / 141 = 0
    16'b01011000_10001110 : OUT <= 0;  //88 / 142 = 0
    16'b01011000_10001111 : OUT <= 0;  //88 / 143 = 0
    16'b01011000_10010000 : OUT <= 0;  //88 / 144 = 0
    16'b01011000_10010001 : OUT <= 0;  //88 / 145 = 0
    16'b01011000_10010010 : OUT <= 0;  //88 / 146 = 0
    16'b01011000_10010011 : OUT <= 0;  //88 / 147 = 0
    16'b01011000_10010100 : OUT <= 0;  //88 / 148 = 0
    16'b01011000_10010101 : OUT <= 0;  //88 / 149 = 0
    16'b01011000_10010110 : OUT <= 0;  //88 / 150 = 0
    16'b01011000_10010111 : OUT <= 0;  //88 / 151 = 0
    16'b01011000_10011000 : OUT <= 0;  //88 / 152 = 0
    16'b01011000_10011001 : OUT <= 0;  //88 / 153 = 0
    16'b01011000_10011010 : OUT <= 0;  //88 / 154 = 0
    16'b01011000_10011011 : OUT <= 0;  //88 / 155 = 0
    16'b01011000_10011100 : OUT <= 0;  //88 / 156 = 0
    16'b01011000_10011101 : OUT <= 0;  //88 / 157 = 0
    16'b01011000_10011110 : OUT <= 0;  //88 / 158 = 0
    16'b01011000_10011111 : OUT <= 0;  //88 / 159 = 0
    16'b01011000_10100000 : OUT <= 0;  //88 / 160 = 0
    16'b01011000_10100001 : OUT <= 0;  //88 / 161 = 0
    16'b01011000_10100010 : OUT <= 0;  //88 / 162 = 0
    16'b01011000_10100011 : OUT <= 0;  //88 / 163 = 0
    16'b01011000_10100100 : OUT <= 0;  //88 / 164 = 0
    16'b01011000_10100101 : OUT <= 0;  //88 / 165 = 0
    16'b01011000_10100110 : OUT <= 0;  //88 / 166 = 0
    16'b01011000_10100111 : OUT <= 0;  //88 / 167 = 0
    16'b01011000_10101000 : OUT <= 0;  //88 / 168 = 0
    16'b01011000_10101001 : OUT <= 0;  //88 / 169 = 0
    16'b01011000_10101010 : OUT <= 0;  //88 / 170 = 0
    16'b01011000_10101011 : OUT <= 0;  //88 / 171 = 0
    16'b01011000_10101100 : OUT <= 0;  //88 / 172 = 0
    16'b01011000_10101101 : OUT <= 0;  //88 / 173 = 0
    16'b01011000_10101110 : OUT <= 0;  //88 / 174 = 0
    16'b01011000_10101111 : OUT <= 0;  //88 / 175 = 0
    16'b01011000_10110000 : OUT <= 0;  //88 / 176 = 0
    16'b01011000_10110001 : OUT <= 0;  //88 / 177 = 0
    16'b01011000_10110010 : OUT <= 0;  //88 / 178 = 0
    16'b01011000_10110011 : OUT <= 0;  //88 / 179 = 0
    16'b01011000_10110100 : OUT <= 0;  //88 / 180 = 0
    16'b01011000_10110101 : OUT <= 0;  //88 / 181 = 0
    16'b01011000_10110110 : OUT <= 0;  //88 / 182 = 0
    16'b01011000_10110111 : OUT <= 0;  //88 / 183 = 0
    16'b01011000_10111000 : OUT <= 0;  //88 / 184 = 0
    16'b01011000_10111001 : OUT <= 0;  //88 / 185 = 0
    16'b01011000_10111010 : OUT <= 0;  //88 / 186 = 0
    16'b01011000_10111011 : OUT <= 0;  //88 / 187 = 0
    16'b01011000_10111100 : OUT <= 0;  //88 / 188 = 0
    16'b01011000_10111101 : OUT <= 0;  //88 / 189 = 0
    16'b01011000_10111110 : OUT <= 0;  //88 / 190 = 0
    16'b01011000_10111111 : OUT <= 0;  //88 / 191 = 0
    16'b01011000_11000000 : OUT <= 0;  //88 / 192 = 0
    16'b01011000_11000001 : OUT <= 0;  //88 / 193 = 0
    16'b01011000_11000010 : OUT <= 0;  //88 / 194 = 0
    16'b01011000_11000011 : OUT <= 0;  //88 / 195 = 0
    16'b01011000_11000100 : OUT <= 0;  //88 / 196 = 0
    16'b01011000_11000101 : OUT <= 0;  //88 / 197 = 0
    16'b01011000_11000110 : OUT <= 0;  //88 / 198 = 0
    16'b01011000_11000111 : OUT <= 0;  //88 / 199 = 0
    16'b01011000_11001000 : OUT <= 0;  //88 / 200 = 0
    16'b01011000_11001001 : OUT <= 0;  //88 / 201 = 0
    16'b01011000_11001010 : OUT <= 0;  //88 / 202 = 0
    16'b01011000_11001011 : OUT <= 0;  //88 / 203 = 0
    16'b01011000_11001100 : OUT <= 0;  //88 / 204 = 0
    16'b01011000_11001101 : OUT <= 0;  //88 / 205 = 0
    16'b01011000_11001110 : OUT <= 0;  //88 / 206 = 0
    16'b01011000_11001111 : OUT <= 0;  //88 / 207 = 0
    16'b01011000_11010000 : OUT <= 0;  //88 / 208 = 0
    16'b01011000_11010001 : OUT <= 0;  //88 / 209 = 0
    16'b01011000_11010010 : OUT <= 0;  //88 / 210 = 0
    16'b01011000_11010011 : OUT <= 0;  //88 / 211 = 0
    16'b01011000_11010100 : OUT <= 0;  //88 / 212 = 0
    16'b01011000_11010101 : OUT <= 0;  //88 / 213 = 0
    16'b01011000_11010110 : OUT <= 0;  //88 / 214 = 0
    16'b01011000_11010111 : OUT <= 0;  //88 / 215 = 0
    16'b01011000_11011000 : OUT <= 0;  //88 / 216 = 0
    16'b01011000_11011001 : OUT <= 0;  //88 / 217 = 0
    16'b01011000_11011010 : OUT <= 0;  //88 / 218 = 0
    16'b01011000_11011011 : OUT <= 0;  //88 / 219 = 0
    16'b01011000_11011100 : OUT <= 0;  //88 / 220 = 0
    16'b01011000_11011101 : OUT <= 0;  //88 / 221 = 0
    16'b01011000_11011110 : OUT <= 0;  //88 / 222 = 0
    16'b01011000_11011111 : OUT <= 0;  //88 / 223 = 0
    16'b01011000_11100000 : OUT <= 0;  //88 / 224 = 0
    16'b01011000_11100001 : OUT <= 0;  //88 / 225 = 0
    16'b01011000_11100010 : OUT <= 0;  //88 / 226 = 0
    16'b01011000_11100011 : OUT <= 0;  //88 / 227 = 0
    16'b01011000_11100100 : OUT <= 0;  //88 / 228 = 0
    16'b01011000_11100101 : OUT <= 0;  //88 / 229 = 0
    16'b01011000_11100110 : OUT <= 0;  //88 / 230 = 0
    16'b01011000_11100111 : OUT <= 0;  //88 / 231 = 0
    16'b01011000_11101000 : OUT <= 0;  //88 / 232 = 0
    16'b01011000_11101001 : OUT <= 0;  //88 / 233 = 0
    16'b01011000_11101010 : OUT <= 0;  //88 / 234 = 0
    16'b01011000_11101011 : OUT <= 0;  //88 / 235 = 0
    16'b01011000_11101100 : OUT <= 0;  //88 / 236 = 0
    16'b01011000_11101101 : OUT <= 0;  //88 / 237 = 0
    16'b01011000_11101110 : OUT <= 0;  //88 / 238 = 0
    16'b01011000_11101111 : OUT <= 0;  //88 / 239 = 0
    16'b01011000_11110000 : OUT <= 0;  //88 / 240 = 0
    16'b01011000_11110001 : OUT <= 0;  //88 / 241 = 0
    16'b01011000_11110010 : OUT <= 0;  //88 / 242 = 0
    16'b01011000_11110011 : OUT <= 0;  //88 / 243 = 0
    16'b01011000_11110100 : OUT <= 0;  //88 / 244 = 0
    16'b01011000_11110101 : OUT <= 0;  //88 / 245 = 0
    16'b01011000_11110110 : OUT <= 0;  //88 / 246 = 0
    16'b01011000_11110111 : OUT <= 0;  //88 / 247 = 0
    16'b01011000_11111000 : OUT <= 0;  //88 / 248 = 0
    16'b01011000_11111001 : OUT <= 0;  //88 / 249 = 0
    16'b01011000_11111010 : OUT <= 0;  //88 / 250 = 0
    16'b01011000_11111011 : OUT <= 0;  //88 / 251 = 0
    16'b01011000_11111100 : OUT <= 0;  //88 / 252 = 0
    16'b01011000_11111101 : OUT <= 0;  //88 / 253 = 0
    16'b01011000_11111110 : OUT <= 0;  //88 / 254 = 0
    16'b01011000_11111111 : OUT <= 0;  //88 / 255 = 0
    16'b01011001_00000000 : OUT <= 0;  //89 / 0 = 0
    16'b01011001_00000001 : OUT <= 89;  //89 / 1 = 89
    16'b01011001_00000010 : OUT <= 44;  //89 / 2 = 44
    16'b01011001_00000011 : OUT <= 29;  //89 / 3 = 29
    16'b01011001_00000100 : OUT <= 22;  //89 / 4 = 22
    16'b01011001_00000101 : OUT <= 17;  //89 / 5 = 17
    16'b01011001_00000110 : OUT <= 14;  //89 / 6 = 14
    16'b01011001_00000111 : OUT <= 12;  //89 / 7 = 12
    16'b01011001_00001000 : OUT <= 11;  //89 / 8 = 11
    16'b01011001_00001001 : OUT <= 9;  //89 / 9 = 9
    16'b01011001_00001010 : OUT <= 8;  //89 / 10 = 8
    16'b01011001_00001011 : OUT <= 8;  //89 / 11 = 8
    16'b01011001_00001100 : OUT <= 7;  //89 / 12 = 7
    16'b01011001_00001101 : OUT <= 6;  //89 / 13 = 6
    16'b01011001_00001110 : OUT <= 6;  //89 / 14 = 6
    16'b01011001_00001111 : OUT <= 5;  //89 / 15 = 5
    16'b01011001_00010000 : OUT <= 5;  //89 / 16 = 5
    16'b01011001_00010001 : OUT <= 5;  //89 / 17 = 5
    16'b01011001_00010010 : OUT <= 4;  //89 / 18 = 4
    16'b01011001_00010011 : OUT <= 4;  //89 / 19 = 4
    16'b01011001_00010100 : OUT <= 4;  //89 / 20 = 4
    16'b01011001_00010101 : OUT <= 4;  //89 / 21 = 4
    16'b01011001_00010110 : OUT <= 4;  //89 / 22 = 4
    16'b01011001_00010111 : OUT <= 3;  //89 / 23 = 3
    16'b01011001_00011000 : OUT <= 3;  //89 / 24 = 3
    16'b01011001_00011001 : OUT <= 3;  //89 / 25 = 3
    16'b01011001_00011010 : OUT <= 3;  //89 / 26 = 3
    16'b01011001_00011011 : OUT <= 3;  //89 / 27 = 3
    16'b01011001_00011100 : OUT <= 3;  //89 / 28 = 3
    16'b01011001_00011101 : OUT <= 3;  //89 / 29 = 3
    16'b01011001_00011110 : OUT <= 2;  //89 / 30 = 2
    16'b01011001_00011111 : OUT <= 2;  //89 / 31 = 2
    16'b01011001_00100000 : OUT <= 2;  //89 / 32 = 2
    16'b01011001_00100001 : OUT <= 2;  //89 / 33 = 2
    16'b01011001_00100010 : OUT <= 2;  //89 / 34 = 2
    16'b01011001_00100011 : OUT <= 2;  //89 / 35 = 2
    16'b01011001_00100100 : OUT <= 2;  //89 / 36 = 2
    16'b01011001_00100101 : OUT <= 2;  //89 / 37 = 2
    16'b01011001_00100110 : OUT <= 2;  //89 / 38 = 2
    16'b01011001_00100111 : OUT <= 2;  //89 / 39 = 2
    16'b01011001_00101000 : OUT <= 2;  //89 / 40 = 2
    16'b01011001_00101001 : OUT <= 2;  //89 / 41 = 2
    16'b01011001_00101010 : OUT <= 2;  //89 / 42 = 2
    16'b01011001_00101011 : OUT <= 2;  //89 / 43 = 2
    16'b01011001_00101100 : OUT <= 2;  //89 / 44 = 2
    16'b01011001_00101101 : OUT <= 1;  //89 / 45 = 1
    16'b01011001_00101110 : OUT <= 1;  //89 / 46 = 1
    16'b01011001_00101111 : OUT <= 1;  //89 / 47 = 1
    16'b01011001_00110000 : OUT <= 1;  //89 / 48 = 1
    16'b01011001_00110001 : OUT <= 1;  //89 / 49 = 1
    16'b01011001_00110010 : OUT <= 1;  //89 / 50 = 1
    16'b01011001_00110011 : OUT <= 1;  //89 / 51 = 1
    16'b01011001_00110100 : OUT <= 1;  //89 / 52 = 1
    16'b01011001_00110101 : OUT <= 1;  //89 / 53 = 1
    16'b01011001_00110110 : OUT <= 1;  //89 / 54 = 1
    16'b01011001_00110111 : OUT <= 1;  //89 / 55 = 1
    16'b01011001_00111000 : OUT <= 1;  //89 / 56 = 1
    16'b01011001_00111001 : OUT <= 1;  //89 / 57 = 1
    16'b01011001_00111010 : OUT <= 1;  //89 / 58 = 1
    16'b01011001_00111011 : OUT <= 1;  //89 / 59 = 1
    16'b01011001_00111100 : OUT <= 1;  //89 / 60 = 1
    16'b01011001_00111101 : OUT <= 1;  //89 / 61 = 1
    16'b01011001_00111110 : OUT <= 1;  //89 / 62 = 1
    16'b01011001_00111111 : OUT <= 1;  //89 / 63 = 1
    16'b01011001_01000000 : OUT <= 1;  //89 / 64 = 1
    16'b01011001_01000001 : OUT <= 1;  //89 / 65 = 1
    16'b01011001_01000010 : OUT <= 1;  //89 / 66 = 1
    16'b01011001_01000011 : OUT <= 1;  //89 / 67 = 1
    16'b01011001_01000100 : OUT <= 1;  //89 / 68 = 1
    16'b01011001_01000101 : OUT <= 1;  //89 / 69 = 1
    16'b01011001_01000110 : OUT <= 1;  //89 / 70 = 1
    16'b01011001_01000111 : OUT <= 1;  //89 / 71 = 1
    16'b01011001_01001000 : OUT <= 1;  //89 / 72 = 1
    16'b01011001_01001001 : OUT <= 1;  //89 / 73 = 1
    16'b01011001_01001010 : OUT <= 1;  //89 / 74 = 1
    16'b01011001_01001011 : OUT <= 1;  //89 / 75 = 1
    16'b01011001_01001100 : OUT <= 1;  //89 / 76 = 1
    16'b01011001_01001101 : OUT <= 1;  //89 / 77 = 1
    16'b01011001_01001110 : OUT <= 1;  //89 / 78 = 1
    16'b01011001_01001111 : OUT <= 1;  //89 / 79 = 1
    16'b01011001_01010000 : OUT <= 1;  //89 / 80 = 1
    16'b01011001_01010001 : OUT <= 1;  //89 / 81 = 1
    16'b01011001_01010010 : OUT <= 1;  //89 / 82 = 1
    16'b01011001_01010011 : OUT <= 1;  //89 / 83 = 1
    16'b01011001_01010100 : OUT <= 1;  //89 / 84 = 1
    16'b01011001_01010101 : OUT <= 1;  //89 / 85 = 1
    16'b01011001_01010110 : OUT <= 1;  //89 / 86 = 1
    16'b01011001_01010111 : OUT <= 1;  //89 / 87 = 1
    16'b01011001_01011000 : OUT <= 1;  //89 / 88 = 1
    16'b01011001_01011001 : OUT <= 1;  //89 / 89 = 1
    16'b01011001_01011010 : OUT <= 0;  //89 / 90 = 0
    16'b01011001_01011011 : OUT <= 0;  //89 / 91 = 0
    16'b01011001_01011100 : OUT <= 0;  //89 / 92 = 0
    16'b01011001_01011101 : OUT <= 0;  //89 / 93 = 0
    16'b01011001_01011110 : OUT <= 0;  //89 / 94 = 0
    16'b01011001_01011111 : OUT <= 0;  //89 / 95 = 0
    16'b01011001_01100000 : OUT <= 0;  //89 / 96 = 0
    16'b01011001_01100001 : OUT <= 0;  //89 / 97 = 0
    16'b01011001_01100010 : OUT <= 0;  //89 / 98 = 0
    16'b01011001_01100011 : OUT <= 0;  //89 / 99 = 0
    16'b01011001_01100100 : OUT <= 0;  //89 / 100 = 0
    16'b01011001_01100101 : OUT <= 0;  //89 / 101 = 0
    16'b01011001_01100110 : OUT <= 0;  //89 / 102 = 0
    16'b01011001_01100111 : OUT <= 0;  //89 / 103 = 0
    16'b01011001_01101000 : OUT <= 0;  //89 / 104 = 0
    16'b01011001_01101001 : OUT <= 0;  //89 / 105 = 0
    16'b01011001_01101010 : OUT <= 0;  //89 / 106 = 0
    16'b01011001_01101011 : OUT <= 0;  //89 / 107 = 0
    16'b01011001_01101100 : OUT <= 0;  //89 / 108 = 0
    16'b01011001_01101101 : OUT <= 0;  //89 / 109 = 0
    16'b01011001_01101110 : OUT <= 0;  //89 / 110 = 0
    16'b01011001_01101111 : OUT <= 0;  //89 / 111 = 0
    16'b01011001_01110000 : OUT <= 0;  //89 / 112 = 0
    16'b01011001_01110001 : OUT <= 0;  //89 / 113 = 0
    16'b01011001_01110010 : OUT <= 0;  //89 / 114 = 0
    16'b01011001_01110011 : OUT <= 0;  //89 / 115 = 0
    16'b01011001_01110100 : OUT <= 0;  //89 / 116 = 0
    16'b01011001_01110101 : OUT <= 0;  //89 / 117 = 0
    16'b01011001_01110110 : OUT <= 0;  //89 / 118 = 0
    16'b01011001_01110111 : OUT <= 0;  //89 / 119 = 0
    16'b01011001_01111000 : OUT <= 0;  //89 / 120 = 0
    16'b01011001_01111001 : OUT <= 0;  //89 / 121 = 0
    16'b01011001_01111010 : OUT <= 0;  //89 / 122 = 0
    16'b01011001_01111011 : OUT <= 0;  //89 / 123 = 0
    16'b01011001_01111100 : OUT <= 0;  //89 / 124 = 0
    16'b01011001_01111101 : OUT <= 0;  //89 / 125 = 0
    16'b01011001_01111110 : OUT <= 0;  //89 / 126 = 0
    16'b01011001_01111111 : OUT <= 0;  //89 / 127 = 0
    16'b01011001_10000000 : OUT <= 0;  //89 / 128 = 0
    16'b01011001_10000001 : OUT <= 0;  //89 / 129 = 0
    16'b01011001_10000010 : OUT <= 0;  //89 / 130 = 0
    16'b01011001_10000011 : OUT <= 0;  //89 / 131 = 0
    16'b01011001_10000100 : OUT <= 0;  //89 / 132 = 0
    16'b01011001_10000101 : OUT <= 0;  //89 / 133 = 0
    16'b01011001_10000110 : OUT <= 0;  //89 / 134 = 0
    16'b01011001_10000111 : OUT <= 0;  //89 / 135 = 0
    16'b01011001_10001000 : OUT <= 0;  //89 / 136 = 0
    16'b01011001_10001001 : OUT <= 0;  //89 / 137 = 0
    16'b01011001_10001010 : OUT <= 0;  //89 / 138 = 0
    16'b01011001_10001011 : OUT <= 0;  //89 / 139 = 0
    16'b01011001_10001100 : OUT <= 0;  //89 / 140 = 0
    16'b01011001_10001101 : OUT <= 0;  //89 / 141 = 0
    16'b01011001_10001110 : OUT <= 0;  //89 / 142 = 0
    16'b01011001_10001111 : OUT <= 0;  //89 / 143 = 0
    16'b01011001_10010000 : OUT <= 0;  //89 / 144 = 0
    16'b01011001_10010001 : OUT <= 0;  //89 / 145 = 0
    16'b01011001_10010010 : OUT <= 0;  //89 / 146 = 0
    16'b01011001_10010011 : OUT <= 0;  //89 / 147 = 0
    16'b01011001_10010100 : OUT <= 0;  //89 / 148 = 0
    16'b01011001_10010101 : OUT <= 0;  //89 / 149 = 0
    16'b01011001_10010110 : OUT <= 0;  //89 / 150 = 0
    16'b01011001_10010111 : OUT <= 0;  //89 / 151 = 0
    16'b01011001_10011000 : OUT <= 0;  //89 / 152 = 0
    16'b01011001_10011001 : OUT <= 0;  //89 / 153 = 0
    16'b01011001_10011010 : OUT <= 0;  //89 / 154 = 0
    16'b01011001_10011011 : OUT <= 0;  //89 / 155 = 0
    16'b01011001_10011100 : OUT <= 0;  //89 / 156 = 0
    16'b01011001_10011101 : OUT <= 0;  //89 / 157 = 0
    16'b01011001_10011110 : OUT <= 0;  //89 / 158 = 0
    16'b01011001_10011111 : OUT <= 0;  //89 / 159 = 0
    16'b01011001_10100000 : OUT <= 0;  //89 / 160 = 0
    16'b01011001_10100001 : OUT <= 0;  //89 / 161 = 0
    16'b01011001_10100010 : OUT <= 0;  //89 / 162 = 0
    16'b01011001_10100011 : OUT <= 0;  //89 / 163 = 0
    16'b01011001_10100100 : OUT <= 0;  //89 / 164 = 0
    16'b01011001_10100101 : OUT <= 0;  //89 / 165 = 0
    16'b01011001_10100110 : OUT <= 0;  //89 / 166 = 0
    16'b01011001_10100111 : OUT <= 0;  //89 / 167 = 0
    16'b01011001_10101000 : OUT <= 0;  //89 / 168 = 0
    16'b01011001_10101001 : OUT <= 0;  //89 / 169 = 0
    16'b01011001_10101010 : OUT <= 0;  //89 / 170 = 0
    16'b01011001_10101011 : OUT <= 0;  //89 / 171 = 0
    16'b01011001_10101100 : OUT <= 0;  //89 / 172 = 0
    16'b01011001_10101101 : OUT <= 0;  //89 / 173 = 0
    16'b01011001_10101110 : OUT <= 0;  //89 / 174 = 0
    16'b01011001_10101111 : OUT <= 0;  //89 / 175 = 0
    16'b01011001_10110000 : OUT <= 0;  //89 / 176 = 0
    16'b01011001_10110001 : OUT <= 0;  //89 / 177 = 0
    16'b01011001_10110010 : OUT <= 0;  //89 / 178 = 0
    16'b01011001_10110011 : OUT <= 0;  //89 / 179 = 0
    16'b01011001_10110100 : OUT <= 0;  //89 / 180 = 0
    16'b01011001_10110101 : OUT <= 0;  //89 / 181 = 0
    16'b01011001_10110110 : OUT <= 0;  //89 / 182 = 0
    16'b01011001_10110111 : OUT <= 0;  //89 / 183 = 0
    16'b01011001_10111000 : OUT <= 0;  //89 / 184 = 0
    16'b01011001_10111001 : OUT <= 0;  //89 / 185 = 0
    16'b01011001_10111010 : OUT <= 0;  //89 / 186 = 0
    16'b01011001_10111011 : OUT <= 0;  //89 / 187 = 0
    16'b01011001_10111100 : OUT <= 0;  //89 / 188 = 0
    16'b01011001_10111101 : OUT <= 0;  //89 / 189 = 0
    16'b01011001_10111110 : OUT <= 0;  //89 / 190 = 0
    16'b01011001_10111111 : OUT <= 0;  //89 / 191 = 0
    16'b01011001_11000000 : OUT <= 0;  //89 / 192 = 0
    16'b01011001_11000001 : OUT <= 0;  //89 / 193 = 0
    16'b01011001_11000010 : OUT <= 0;  //89 / 194 = 0
    16'b01011001_11000011 : OUT <= 0;  //89 / 195 = 0
    16'b01011001_11000100 : OUT <= 0;  //89 / 196 = 0
    16'b01011001_11000101 : OUT <= 0;  //89 / 197 = 0
    16'b01011001_11000110 : OUT <= 0;  //89 / 198 = 0
    16'b01011001_11000111 : OUT <= 0;  //89 / 199 = 0
    16'b01011001_11001000 : OUT <= 0;  //89 / 200 = 0
    16'b01011001_11001001 : OUT <= 0;  //89 / 201 = 0
    16'b01011001_11001010 : OUT <= 0;  //89 / 202 = 0
    16'b01011001_11001011 : OUT <= 0;  //89 / 203 = 0
    16'b01011001_11001100 : OUT <= 0;  //89 / 204 = 0
    16'b01011001_11001101 : OUT <= 0;  //89 / 205 = 0
    16'b01011001_11001110 : OUT <= 0;  //89 / 206 = 0
    16'b01011001_11001111 : OUT <= 0;  //89 / 207 = 0
    16'b01011001_11010000 : OUT <= 0;  //89 / 208 = 0
    16'b01011001_11010001 : OUT <= 0;  //89 / 209 = 0
    16'b01011001_11010010 : OUT <= 0;  //89 / 210 = 0
    16'b01011001_11010011 : OUT <= 0;  //89 / 211 = 0
    16'b01011001_11010100 : OUT <= 0;  //89 / 212 = 0
    16'b01011001_11010101 : OUT <= 0;  //89 / 213 = 0
    16'b01011001_11010110 : OUT <= 0;  //89 / 214 = 0
    16'b01011001_11010111 : OUT <= 0;  //89 / 215 = 0
    16'b01011001_11011000 : OUT <= 0;  //89 / 216 = 0
    16'b01011001_11011001 : OUT <= 0;  //89 / 217 = 0
    16'b01011001_11011010 : OUT <= 0;  //89 / 218 = 0
    16'b01011001_11011011 : OUT <= 0;  //89 / 219 = 0
    16'b01011001_11011100 : OUT <= 0;  //89 / 220 = 0
    16'b01011001_11011101 : OUT <= 0;  //89 / 221 = 0
    16'b01011001_11011110 : OUT <= 0;  //89 / 222 = 0
    16'b01011001_11011111 : OUT <= 0;  //89 / 223 = 0
    16'b01011001_11100000 : OUT <= 0;  //89 / 224 = 0
    16'b01011001_11100001 : OUT <= 0;  //89 / 225 = 0
    16'b01011001_11100010 : OUT <= 0;  //89 / 226 = 0
    16'b01011001_11100011 : OUT <= 0;  //89 / 227 = 0
    16'b01011001_11100100 : OUT <= 0;  //89 / 228 = 0
    16'b01011001_11100101 : OUT <= 0;  //89 / 229 = 0
    16'b01011001_11100110 : OUT <= 0;  //89 / 230 = 0
    16'b01011001_11100111 : OUT <= 0;  //89 / 231 = 0
    16'b01011001_11101000 : OUT <= 0;  //89 / 232 = 0
    16'b01011001_11101001 : OUT <= 0;  //89 / 233 = 0
    16'b01011001_11101010 : OUT <= 0;  //89 / 234 = 0
    16'b01011001_11101011 : OUT <= 0;  //89 / 235 = 0
    16'b01011001_11101100 : OUT <= 0;  //89 / 236 = 0
    16'b01011001_11101101 : OUT <= 0;  //89 / 237 = 0
    16'b01011001_11101110 : OUT <= 0;  //89 / 238 = 0
    16'b01011001_11101111 : OUT <= 0;  //89 / 239 = 0
    16'b01011001_11110000 : OUT <= 0;  //89 / 240 = 0
    16'b01011001_11110001 : OUT <= 0;  //89 / 241 = 0
    16'b01011001_11110010 : OUT <= 0;  //89 / 242 = 0
    16'b01011001_11110011 : OUT <= 0;  //89 / 243 = 0
    16'b01011001_11110100 : OUT <= 0;  //89 / 244 = 0
    16'b01011001_11110101 : OUT <= 0;  //89 / 245 = 0
    16'b01011001_11110110 : OUT <= 0;  //89 / 246 = 0
    16'b01011001_11110111 : OUT <= 0;  //89 / 247 = 0
    16'b01011001_11111000 : OUT <= 0;  //89 / 248 = 0
    16'b01011001_11111001 : OUT <= 0;  //89 / 249 = 0
    16'b01011001_11111010 : OUT <= 0;  //89 / 250 = 0
    16'b01011001_11111011 : OUT <= 0;  //89 / 251 = 0
    16'b01011001_11111100 : OUT <= 0;  //89 / 252 = 0
    16'b01011001_11111101 : OUT <= 0;  //89 / 253 = 0
    16'b01011001_11111110 : OUT <= 0;  //89 / 254 = 0
    16'b01011001_11111111 : OUT <= 0;  //89 / 255 = 0
    16'b01011010_00000000 : OUT <= 0;  //90 / 0 = 0
    16'b01011010_00000001 : OUT <= 90;  //90 / 1 = 90
    16'b01011010_00000010 : OUT <= 45;  //90 / 2 = 45
    16'b01011010_00000011 : OUT <= 30;  //90 / 3 = 30
    16'b01011010_00000100 : OUT <= 22;  //90 / 4 = 22
    16'b01011010_00000101 : OUT <= 18;  //90 / 5 = 18
    16'b01011010_00000110 : OUT <= 15;  //90 / 6 = 15
    16'b01011010_00000111 : OUT <= 12;  //90 / 7 = 12
    16'b01011010_00001000 : OUT <= 11;  //90 / 8 = 11
    16'b01011010_00001001 : OUT <= 10;  //90 / 9 = 10
    16'b01011010_00001010 : OUT <= 9;  //90 / 10 = 9
    16'b01011010_00001011 : OUT <= 8;  //90 / 11 = 8
    16'b01011010_00001100 : OUT <= 7;  //90 / 12 = 7
    16'b01011010_00001101 : OUT <= 6;  //90 / 13 = 6
    16'b01011010_00001110 : OUT <= 6;  //90 / 14 = 6
    16'b01011010_00001111 : OUT <= 6;  //90 / 15 = 6
    16'b01011010_00010000 : OUT <= 5;  //90 / 16 = 5
    16'b01011010_00010001 : OUT <= 5;  //90 / 17 = 5
    16'b01011010_00010010 : OUT <= 5;  //90 / 18 = 5
    16'b01011010_00010011 : OUT <= 4;  //90 / 19 = 4
    16'b01011010_00010100 : OUT <= 4;  //90 / 20 = 4
    16'b01011010_00010101 : OUT <= 4;  //90 / 21 = 4
    16'b01011010_00010110 : OUT <= 4;  //90 / 22 = 4
    16'b01011010_00010111 : OUT <= 3;  //90 / 23 = 3
    16'b01011010_00011000 : OUT <= 3;  //90 / 24 = 3
    16'b01011010_00011001 : OUT <= 3;  //90 / 25 = 3
    16'b01011010_00011010 : OUT <= 3;  //90 / 26 = 3
    16'b01011010_00011011 : OUT <= 3;  //90 / 27 = 3
    16'b01011010_00011100 : OUT <= 3;  //90 / 28 = 3
    16'b01011010_00011101 : OUT <= 3;  //90 / 29 = 3
    16'b01011010_00011110 : OUT <= 3;  //90 / 30 = 3
    16'b01011010_00011111 : OUT <= 2;  //90 / 31 = 2
    16'b01011010_00100000 : OUT <= 2;  //90 / 32 = 2
    16'b01011010_00100001 : OUT <= 2;  //90 / 33 = 2
    16'b01011010_00100010 : OUT <= 2;  //90 / 34 = 2
    16'b01011010_00100011 : OUT <= 2;  //90 / 35 = 2
    16'b01011010_00100100 : OUT <= 2;  //90 / 36 = 2
    16'b01011010_00100101 : OUT <= 2;  //90 / 37 = 2
    16'b01011010_00100110 : OUT <= 2;  //90 / 38 = 2
    16'b01011010_00100111 : OUT <= 2;  //90 / 39 = 2
    16'b01011010_00101000 : OUT <= 2;  //90 / 40 = 2
    16'b01011010_00101001 : OUT <= 2;  //90 / 41 = 2
    16'b01011010_00101010 : OUT <= 2;  //90 / 42 = 2
    16'b01011010_00101011 : OUT <= 2;  //90 / 43 = 2
    16'b01011010_00101100 : OUT <= 2;  //90 / 44 = 2
    16'b01011010_00101101 : OUT <= 2;  //90 / 45 = 2
    16'b01011010_00101110 : OUT <= 1;  //90 / 46 = 1
    16'b01011010_00101111 : OUT <= 1;  //90 / 47 = 1
    16'b01011010_00110000 : OUT <= 1;  //90 / 48 = 1
    16'b01011010_00110001 : OUT <= 1;  //90 / 49 = 1
    16'b01011010_00110010 : OUT <= 1;  //90 / 50 = 1
    16'b01011010_00110011 : OUT <= 1;  //90 / 51 = 1
    16'b01011010_00110100 : OUT <= 1;  //90 / 52 = 1
    16'b01011010_00110101 : OUT <= 1;  //90 / 53 = 1
    16'b01011010_00110110 : OUT <= 1;  //90 / 54 = 1
    16'b01011010_00110111 : OUT <= 1;  //90 / 55 = 1
    16'b01011010_00111000 : OUT <= 1;  //90 / 56 = 1
    16'b01011010_00111001 : OUT <= 1;  //90 / 57 = 1
    16'b01011010_00111010 : OUT <= 1;  //90 / 58 = 1
    16'b01011010_00111011 : OUT <= 1;  //90 / 59 = 1
    16'b01011010_00111100 : OUT <= 1;  //90 / 60 = 1
    16'b01011010_00111101 : OUT <= 1;  //90 / 61 = 1
    16'b01011010_00111110 : OUT <= 1;  //90 / 62 = 1
    16'b01011010_00111111 : OUT <= 1;  //90 / 63 = 1
    16'b01011010_01000000 : OUT <= 1;  //90 / 64 = 1
    16'b01011010_01000001 : OUT <= 1;  //90 / 65 = 1
    16'b01011010_01000010 : OUT <= 1;  //90 / 66 = 1
    16'b01011010_01000011 : OUT <= 1;  //90 / 67 = 1
    16'b01011010_01000100 : OUT <= 1;  //90 / 68 = 1
    16'b01011010_01000101 : OUT <= 1;  //90 / 69 = 1
    16'b01011010_01000110 : OUT <= 1;  //90 / 70 = 1
    16'b01011010_01000111 : OUT <= 1;  //90 / 71 = 1
    16'b01011010_01001000 : OUT <= 1;  //90 / 72 = 1
    16'b01011010_01001001 : OUT <= 1;  //90 / 73 = 1
    16'b01011010_01001010 : OUT <= 1;  //90 / 74 = 1
    16'b01011010_01001011 : OUT <= 1;  //90 / 75 = 1
    16'b01011010_01001100 : OUT <= 1;  //90 / 76 = 1
    16'b01011010_01001101 : OUT <= 1;  //90 / 77 = 1
    16'b01011010_01001110 : OUT <= 1;  //90 / 78 = 1
    16'b01011010_01001111 : OUT <= 1;  //90 / 79 = 1
    16'b01011010_01010000 : OUT <= 1;  //90 / 80 = 1
    16'b01011010_01010001 : OUT <= 1;  //90 / 81 = 1
    16'b01011010_01010010 : OUT <= 1;  //90 / 82 = 1
    16'b01011010_01010011 : OUT <= 1;  //90 / 83 = 1
    16'b01011010_01010100 : OUT <= 1;  //90 / 84 = 1
    16'b01011010_01010101 : OUT <= 1;  //90 / 85 = 1
    16'b01011010_01010110 : OUT <= 1;  //90 / 86 = 1
    16'b01011010_01010111 : OUT <= 1;  //90 / 87 = 1
    16'b01011010_01011000 : OUT <= 1;  //90 / 88 = 1
    16'b01011010_01011001 : OUT <= 1;  //90 / 89 = 1
    16'b01011010_01011010 : OUT <= 1;  //90 / 90 = 1
    16'b01011010_01011011 : OUT <= 0;  //90 / 91 = 0
    16'b01011010_01011100 : OUT <= 0;  //90 / 92 = 0
    16'b01011010_01011101 : OUT <= 0;  //90 / 93 = 0
    16'b01011010_01011110 : OUT <= 0;  //90 / 94 = 0
    16'b01011010_01011111 : OUT <= 0;  //90 / 95 = 0
    16'b01011010_01100000 : OUT <= 0;  //90 / 96 = 0
    16'b01011010_01100001 : OUT <= 0;  //90 / 97 = 0
    16'b01011010_01100010 : OUT <= 0;  //90 / 98 = 0
    16'b01011010_01100011 : OUT <= 0;  //90 / 99 = 0
    16'b01011010_01100100 : OUT <= 0;  //90 / 100 = 0
    16'b01011010_01100101 : OUT <= 0;  //90 / 101 = 0
    16'b01011010_01100110 : OUT <= 0;  //90 / 102 = 0
    16'b01011010_01100111 : OUT <= 0;  //90 / 103 = 0
    16'b01011010_01101000 : OUT <= 0;  //90 / 104 = 0
    16'b01011010_01101001 : OUT <= 0;  //90 / 105 = 0
    16'b01011010_01101010 : OUT <= 0;  //90 / 106 = 0
    16'b01011010_01101011 : OUT <= 0;  //90 / 107 = 0
    16'b01011010_01101100 : OUT <= 0;  //90 / 108 = 0
    16'b01011010_01101101 : OUT <= 0;  //90 / 109 = 0
    16'b01011010_01101110 : OUT <= 0;  //90 / 110 = 0
    16'b01011010_01101111 : OUT <= 0;  //90 / 111 = 0
    16'b01011010_01110000 : OUT <= 0;  //90 / 112 = 0
    16'b01011010_01110001 : OUT <= 0;  //90 / 113 = 0
    16'b01011010_01110010 : OUT <= 0;  //90 / 114 = 0
    16'b01011010_01110011 : OUT <= 0;  //90 / 115 = 0
    16'b01011010_01110100 : OUT <= 0;  //90 / 116 = 0
    16'b01011010_01110101 : OUT <= 0;  //90 / 117 = 0
    16'b01011010_01110110 : OUT <= 0;  //90 / 118 = 0
    16'b01011010_01110111 : OUT <= 0;  //90 / 119 = 0
    16'b01011010_01111000 : OUT <= 0;  //90 / 120 = 0
    16'b01011010_01111001 : OUT <= 0;  //90 / 121 = 0
    16'b01011010_01111010 : OUT <= 0;  //90 / 122 = 0
    16'b01011010_01111011 : OUT <= 0;  //90 / 123 = 0
    16'b01011010_01111100 : OUT <= 0;  //90 / 124 = 0
    16'b01011010_01111101 : OUT <= 0;  //90 / 125 = 0
    16'b01011010_01111110 : OUT <= 0;  //90 / 126 = 0
    16'b01011010_01111111 : OUT <= 0;  //90 / 127 = 0
    16'b01011010_10000000 : OUT <= 0;  //90 / 128 = 0
    16'b01011010_10000001 : OUT <= 0;  //90 / 129 = 0
    16'b01011010_10000010 : OUT <= 0;  //90 / 130 = 0
    16'b01011010_10000011 : OUT <= 0;  //90 / 131 = 0
    16'b01011010_10000100 : OUT <= 0;  //90 / 132 = 0
    16'b01011010_10000101 : OUT <= 0;  //90 / 133 = 0
    16'b01011010_10000110 : OUT <= 0;  //90 / 134 = 0
    16'b01011010_10000111 : OUT <= 0;  //90 / 135 = 0
    16'b01011010_10001000 : OUT <= 0;  //90 / 136 = 0
    16'b01011010_10001001 : OUT <= 0;  //90 / 137 = 0
    16'b01011010_10001010 : OUT <= 0;  //90 / 138 = 0
    16'b01011010_10001011 : OUT <= 0;  //90 / 139 = 0
    16'b01011010_10001100 : OUT <= 0;  //90 / 140 = 0
    16'b01011010_10001101 : OUT <= 0;  //90 / 141 = 0
    16'b01011010_10001110 : OUT <= 0;  //90 / 142 = 0
    16'b01011010_10001111 : OUT <= 0;  //90 / 143 = 0
    16'b01011010_10010000 : OUT <= 0;  //90 / 144 = 0
    16'b01011010_10010001 : OUT <= 0;  //90 / 145 = 0
    16'b01011010_10010010 : OUT <= 0;  //90 / 146 = 0
    16'b01011010_10010011 : OUT <= 0;  //90 / 147 = 0
    16'b01011010_10010100 : OUT <= 0;  //90 / 148 = 0
    16'b01011010_10010101 : OUT <= 0;  //90 / 149 = 0
    16'b01011010_10010110 : OUT <= 0;  //90 / 150 = 0
    16'b01011010_10010111 : OUT <= 0;  //90 / 151 = 0
    16'b01011010_10011000 : OUT <= 0;  //90 / 152 = 0
    16'b01011010_10011001 : OUT <= 0;  //90 / 153 = 0
    16'b01011010_10011010 : OUT <= 0;  //90 / 154 = 0
    16'b01011010_10011011 : OUT <= 0;  //90 / 155 = 0
    16'b01011010_10011100 : OUT <= 0;  //90 / 156 = 0
    16'b01011010_10011101 : OUT <= 0;  //90 / 157 = 0
    16'b01011010_10011110 : OUT <= 0;  //90 / 158 = 0
    16'b01011010_10011111 : OUT <= 0;  //90 / 159 = 0
    16'b01011010_10100000 : OUT <= 0;  //90 / 160 = 0
    16'b01011010_10100001 : OUT <= 0;  //90 / 161 = 0
    16'b01011010_10100010 : OUT <= 0;  //90 / 162 = 0
    16'b01011010_10100011 : OUT <= 0;  //90 / 163 = 0
    16'b01011010_10100100 : OUT <= 0;  //90 / 164 = 0
    16'b01011010_10100101 : OUT <= 0;  //90 / 165 = 0
    16'b01011010_10100110 : OUT <= 0;  //90 / 166 = 0
    16'b01011010_10100111 : OUT <= 0;  //90 / 167 = 0
    16'b01011010_10101000 : OUT <= 0;  //90 / 168 = 0
    16'b01011010_10101001 : OUT <= 0;  //90 / 169 = 0
    16'b01011010_10101010 : OUT <= 0;  //90 / 170 = 0
    16'b01011010_10101011 : OUT <= 0;  //90 / 171 = 0
    16'b01011010_10101100 : OUT <= 0;  //90 / 172 = 0
    16'b01011010_10101101 : OUT <= 0;  //90 / 173 = 0
    16'b01011010_10101110 : OUT <= 0;  //90 / 174 = 0
    16'b01011010_10101111 : OUT <= 0;  //90 / 175 = 0
    16'b01011010_10110000 : OUT <= 0;  //90 / 176 = 0
    16'b01011010_10110001 : OUT <= 0;  //90 / 177 = 0
    16'b01011010_10110010 : OUT <= 0;  //90 / 178 = 0
    16'b01011010_10110011 : OUT <= 0;  //90 / 179 = 0
    16'b01011010_10110100 : OUT <= 0;  //90 / 180 = 0
    16'b01011010_10110101 : OUT <= 0;  //90 / 181 = 0
    16'b01011010_10110110 : OUT <= 0;  //90 / 182 = 0
    16'b01011010_10110111 : OUT <= 0;  //90 / 183 = 0
    16'b01011010_10111000 : OUT <= 0;  //90 / 184 = 0
    16'b01011010_10111001 : OUT <= 0;  //90 / 185 = 0
    16'b01011010_10111010 : OUT <= 0;  //90 / 186 = 0
    16'b01011010_10111011 : OUT <= 0;  //90 / 187 = 0
    16'b01011010_10111100 : OUT <= 0;  //90 / 188 = 0
    16'b01011010_10111101 : OUT <= 0;  //90 / 189 = 0
    16'b01011010_10111110 : OUT <= 0;  //90 / 190 = 0
    16'b01011010_10111111 : OUT <= 0;  //90 / 191 = 0
    16'b01011010_11000000 : OUT <= 0;  //90 / 192 = 0
    16'b01011010_11000001 : OUT <= 0;  //90 / 193 = 0
    16'b01011010_11000010 : OUT <= 0;  //90 / 194 = 0
    16'b01011010_11000011 : OUT <= 0;  //90 / 195 = 0
    16'b01011010_11000100 : OUT <= 0;  //90 / 196 = 0
    16'b01011010_11000101 : OUT <= 0;  //90 / 197 = 0
    16'b01011010_11000110 : OUT <= 0;  //90 / 198 = 0
    16'b01011010_11000111 : OUT <= 0;  //90 / 199 = 0
    16'b01011010_11001000 : OUT <= 0;  //90 / 200 = 0
    16'b01011010_11001001 : OUT <= 0;  //90 / 201 = 0
    16'b01011010_11001010 : OUT <= 0;  //90 / 202 = 0
    16'b01011010_11001011 : OUT <= 0;  //90 / 203 = 0
    16'b01011010_11001100 : OUT <= 0;  //90 / 204 = 0
    16'b01011010_11001101 : OUT <= 0;  //90 / 205 = 0
    16'b01011010_11001110 : OUT <= 0;  //90 / 206 = 0
    16'b01011010_11001111 : OUT <= 0;  //90 / 207 = 0
    16'b01011010_11010000 : OUT <= 0;  //90 / 208 = 0
    16'b01011010_11010001 : OUT <= 0;  //90 / 209 = 0
    16'b01011010_11010010 : OUT <= 0;  //90 / 210 = 0
    16'b01011010_11010011 : OUT <= 0;  //90 / 211 = 0
    16'b01011010_11010100 : OUT <= 0;  //90 / 212 = 0
    16'b01011010_11010101 : OUT <= 0;  //90 / 213 = 0
    16'b01011010_11010110 : OUT <= 0;  //90 / 214 = 0
    16'b01011010_11010111 : OUT <= 0;  //90 / 215 = 0
    16'b01011010_11011000 : OUT <= 0;  //90 / 216 = 0
    16'b01011010_11011001 : OUT <= 0;  //90 / 217 = 0
    16'b01011010_11011010 : OUT <= 0;  //90 / 218 = 0
    16'b01011010_11011011 : OUT <= 0;  //90 / 219 = 0
    16'b01011010_11011100 : OUT <= 0;  //90 / 220 = 0
    16'b01011010_11011101 : OUT <= 0;  //90 / 221 = 0
    16'b01011010_11011110 : OUT <= 0;  //90 / 222 = 0
    16'b01011010_11011111 : OUT <= 0;  //90 / 223 = 0
    16'b01011010_11100000 : OUT <= 0;  //90 / 224 = 0
    16'b01011010_11100001 : OUT <= 0;  //90 / 225 = 0
    16'b01011010_11100010 : OUT <= 0;  //90 / 226 = 0
    16'b01011010_11100011 : OUT <= 0;  //90 / 227 = 0
    16'b01011010_11100100 : OUT <= 0;  //90 / 228 = 0
    16'b01011010_11100101 : OUT <= 0;  //90 / 229 = 0
    16'b01011010_11100110 : OUT <= 0;  //90 / 230 = 0
    16'b01011010_11100111 : OUT <= 0;  //90 / 231 = 0
    16'b01011010_11101000 : OUT <= 0;  //90 / 232 = 0
    16'b01011010_11101001 : OUT <= 0;  //90 / 233 = 0
    16'b01011010_11101010 : OUT <= 0;  //90 / 234 = 0
    16'b01011010_11101011 : OUT <= 0;  //90 / 235 = 0
    16'b01011010_11101100 : OUT <= 0;  //90 / 236 = 0
    16'b01011010_11101101 : OUT <= 0;  //90 / 237 = 0
    16'b01011010_11101110 : OUT <= 0;  //90 / 238 = 0
    16'b01011010_11101111 : OUT <= 0;  //90 / 239 = 0
    16'b01011010_11110000 : OUT <= 0;  //90 / 240 = 0
    16'b01011010_11110001 : OUT <= 0;  //90 / 241 = 0
    16'b01011010_11110010 : OUT <= 0;  //90 / 242 = 0
    16'b01011010_11110011 : OUT <= 0;  //90 / 243 = 0
    16'b01011010_11110100 : OUT <= 0;  //90 / 244 = 0
    16'b01011010_11110101 : OUT <= 0;  //90 / 245 = 0
    16'b01011010_11110110 : OUT <= 0;  //90 / 246 = 0
    16'b01011010_11110111 : OUT <= 0;  //90 / 247 = 0
    16'b01011010_11111000 : OUT <= 0;  //90 / 248 = 0
    16'b01011010_11111001 : OUT <= 0;  //90 / 249 = 0
    16'b01011010_11111010 : OUT <= 0;  //90 / 250 = 0
    16'b01011010_11111011 : OUT <= 0;  //90 / 251 = 0
    16'b01011010_11111100 : OUT <= 0;  //90 / 252 = 0
    16'b01011010_11111101 : OUT <= 0;  //90 / 253 = 0
    16'b01011010_11111110 : OUT <= 0;  //90 / 254 = 0
    16'b01011010_11111111 : OUT <= 0;  //90 / 255 = 0
    16'b01011011_00000000 : OUT <= 0;  //91 / 0 = 0
    16'b01011011_00000001 : OUT <= 91;  //91 / 1 = 91
    16'b01011011_00000010 : OUT <= 45;  //91 / 2 = 45
    16'b01011011_00000011 : OUT <= 30;  //91 / 3 = 30
    16'b01011011_00000100 : OUT <= 22;  //91 / 4 = 22
    16'b01011011_00000101 : OUT <= 18;  //91 / 5 = 18
    16'b01011011_00000110 : OUT <= 15;  //91 / 6 = 15
    16'b01011011_00000111 : OUT <= 13;  //91 / 7 = 13
    16'b01011011_00001000 : OUT <= 11;  //91 / 8 = 11
    16'b01011011_00001001 : OUT <= 10;  //91 / 9 = 10
    16'b01011011_00001010 : OUT <= 9;  //91 / 10 = 9
    16'b01011011_00001011 : OUT <= 8;  //91 / 11 = 8
    16'b01011011_00001100 : OUT <= 7;  //91 / 12 = 7
    16'b01011011_00001101 : OUT <= 7;  //91 / 13 = 7
    16'b01011011_00001110 : OUT <= 6;  //91 / 14 = 6
    16'b01011011_00001111 : OUT <= 6;  //91 / 15 = 6
    16'b01011011_00010000 : OUT <= 5;  //91 / 16 = 5
    16'b01011011_00010001 : OUT <= 5;  //91 / 17 = 5
    16'b01011011_00010010 : OUT <= 5;  //91 / 18 = 5
    16'b01011011_00010011 : OUT <= 4;  //91 / 19 = 4
    16'b01011011_00010100 : OUT <= 4;  //91 / 20 = 4
    16'b01011011_00010101 : OUT <= 4;  //91 / 21 = 4
    16'b01011011_00010110 : OUT <= 4;  //91 / 22 = 4
    16'b01011011_00010111 : OUT <= 3;  //91 / 23 = 3
    16'b01011011_00011000 : OUT <= 3;  //91 / 24 = 3
    16'b01011011_00011001 : OUT <= 3;  //91 / 25 = 3
    16'b01011011_00011010 : OUT <= 3;  //91 / 26 = 3
    16'b01011011_00011011 : OUT <= 3;  //91 / 27 = 3
    16'b01011011_00011100 : OUT <= 3;  //91 / 28 = 3
    16'b01011011_00011101 : OUT <= 3;  //91 / 29 = 3
    16'b01011011_00011110 : OUT <= 3;  //91 / 30 = 3
    16'b01011011_00011111 : OUT <= 2;  //91 / 31 = 2
    16'b01011011_00100000 : OUT <= 2;  //91 / 32 = 2
    16'b01011011_00100001 : OUT <= 2;  //91 / 33 = 2
    16'b01011011_00100010 : OUT <= 2;  //91 / 34 = 2
    16'b01011011_00100011 : OUT <= 2;  //91 / 35 = 2
    16'b01011011_00100100 : OUT <= 2;  //91 / 36 = 2
    16'b01011011_00100101 : OUT <= 2;  //91 / 37 = 2
    16'b01011011_00100110 : OUT <= 2;  //91 / 38 = 2
    16'b01011011_00100111 : OUT <= 2;  //91 / 39 = 2
    16'b01011011_00101000 : OUT <= 2;  //91 / 40 = 2
    16'b01011011_00101001 : OUT <= 2;  //91 / 41 = 2
    16'b01011011_00101010 : OUT <= 2;  //91 / 42 = 2
    16'b01011011_00101011 : OUT <= 2;  //91 / 43 = 2
    16'b01011011_00101100 : OUT <= 2;  //91 / 44 = 2
    16'b01011011_00101101 : OUT <= 2;  //91 / 45 = 2
    16'b01011011_00101110 : OUT <= 1;  //91 / 46 = 1
    16'b01011011_00101111 : OUT <= 1;  //91 / 47 = 1
    16'b01011011_00110000 : OUT <= 1;  //91 / 48 = 1
    16'b01011011_00110001 : OUT <= 1;  //91 / 49 = 1
    16'b01011011_00110010 : OUT <= 1;  //91 / 50 = 1
    16'b01011011_00110011 : OUT <= 1;  //91 / 51 = 1
    16'b01011011_00110100 : OUT <= 1;  //91 / 52 = 1
    16'b01011011_00110101 : OUT <= 1;  //91 / 53 = 1
    16'b01011011_00110110 : OUT <= 1;  //91 / 54 = 1
    16'b01011011_00110111 : OUT <= 1;  //91 / 55 = 1
    16'b01011011_00111000 : OUT <= 1;  //91 / 56 = 1
    16'b01011011_00111001 : OUT <= 1;  //91 / 57 = 1
    16'b01011011_00111010 : OUT <= 1;  //91 / 58 = 1
    16'b01011011_00111011 : OUT <= 1;  //91 / 59 = 1
    16'b01011011_00111100 : OUT <= 1;  //91 / 60 = 1
    16'b01011011_00111101 : OUT <= 1;  //91 / 61 = 1
    16'b01011011_00111110 : OUT <= 1;  //91 / 62 = 1
    16'b01011011_00111111 : OUT <= 1;  //91 / 63 = 1
    16'b01011011_01000000 : OUT <= 1;  //91 / 64 = 1
    16'b01011011_01000001 : OUT <= 1;  //91 / 65 = 1
    16'b01011011_01000010 : OUT <= 1;  //91 / 66 = 1
    16'b01011011_01000011 : OUT <= 1;  //91 / 67 = 1
    16'b01011011_01000100 : OUT <= 1;  //91 / 68 = 1
    16'b01011011_01000101 : OUT <= 1;  //91 / 69 = 1
    16'b01011011_01000110 : OUT <= 1;  //91 / 70 = 1
    16'b01011011_01000111 : OUT <= 1;  //91 / 71 = 1
    16'b01011011_01001000 : OUT <= 1;  //91 / 72 = 1
    16'b01011011_01001001 : OUT <= 1;  //91 / 73 = 1
    16'b01011011_01001010 : OUT <= 1;  //91 / 74 = 1
    16'b01011011_01001011 : OUT <= 1;  //91 / 75 = 1
    16'b01011011_01001100 : OUT <= 1;  //91 / 76 = 1
    16'b01011011_01001101 : OUT <= 1;  //91 / 77 = 1
    16'b01011011_01001110 : OUT <= 1;  //91 / 78 = 1
    16'b01011011_01001111 : OUT <= 1;  //91 / 79 = 1
    16'b01011011_01010000 : OUT <= 1;  //91 / 80 = 1
    16'b01011011_01010001 : OUT <= 1;  //91 / 81 = 1
    16'b01011011_01010010 : OUT <= 1;  //91 / 82 = 1
    16'b01011011_01010011 : OUT <= 1;  //91 / 83 = 1
    16'b01011011_01010100 : OUT <= 1;  //91 / 84 = 1
    16'b01011011_01010101 : OUT <= 1;  //91 / 85 = 1
    16'b01011011_01010110 : OUT <= 1;  //91 / 86 = 1
    16'b01011011_01010111 : OUT <= 1;  //91 / 87 = 1
    16'b01011011_01011000 : OUT <= 1;  //91 / 88 = 1
    16'b01011011_01011001 : OUT <= 1;  //91 / 89 = 1
    16'b01011011_01011010 : OUT <= 1;  //91 / 90 = 1
    16'b01011011_01011011 : OUT <= 1;  //91 / 91 = 1
    16'b01011011_01011100 : OUT <= 0;  //91 / 92 = 0
    16'b01011011_01011101 : OUT <= 0;  //91 / 93 = 0
    16'b01011011_01011110 : OUT <= 0;  //91 / 94 = 0
    16'b01011011_01011111 : OUT <= 0;  //91 / 95 = 0
    16'b01011011_01100000 : OUT <= 0;  //91 / 96 = 0
    16'b01011011_01100001 : OUT <= 0;  //91 / 97 = 0
    16'b01011011_01100010 : OUT <= 0;  //91 / 98 = 0
    16'b01011011_01100011 : OUT <= 0;  //91 / 99 = 0
    16'b01011011_01100100 : OUT <= 0;  //91 / 100 = 0
    16'b01011011_01100101 : OUT <= 0;  //91 / 101 = 0
    16'b01011011_01100110 : OUT <= 0;  //91 / 102 = 0
    16'b01011011_01100111 : OUT <= 0;  //91 / 103 = 0
    16'b01011011_01101000 : OUT <= 0;  //91 / 104 = 0
    16'b01011011_01101001 : OUT <= 0;  //91 / 105 = 0
    16'b01011011_01101010 : OUT <= 0;  //91 / 106 = 0
    16'b01011011_01101011 : OUT <= 0;  //91 / 107 = 0
    16'b01011011_01101100 : OUT <= 0;  //91 / 108 = 0
    16'b01011011_01101101 : OUT <= 0;  //91 / 109 = 0
    16'b01011011_01101110 : OUT <= 0;  //91 / 110 = 0
    16'b01011011_01101111 : OUT <= 0;  //91 / 111 = 0
    16'b01011011_01110000 : OUT <= 0;  //91 / 112 = 0
    16'b01011011_01110001 : OUT <= 0;  //91 / 113 = 0
    16'b01011011_01110010 : OUT <= 0;  //91 / 114 = 0
    16'b01011011_01110011 : OUT <= 0;  //91 / 115 = 0
    16'b01011011_01110100 : OUT <= 0;  //91 / 116 = 0
    16'b01011011_01110101 : OUT <= 0;  //91 / 117 = 0
    16'b01011011_01110110 : OUT <= 0;  //91 / 118 = 0
    16'b01011011_01110111 : OUT <= 0;  //91 / 119 = 0
    16'b01011011_01111000 : OUT <= 0;  //91 / 120 = 0
    16'b01011011_01111001 : OUT <= 0;  //91 / 121 = 0
    16'b01011011_01111010 : OUT <= 0;  //91 / 122 = 0
    16'b01011011_01111011 : OUT <= 0;  //91 / 123 = 0
    16'b01011011_01111100 : OUT <= 0;  //91 / 124 = 0
    16'b01011011_01111101 : OUT <= 0;  //91 / 125 = 0
    16'b01011011_01111110 : OUT <= 0;  //91 / 126 = 0
    16'b01011011_01111111 : OUT <= 0;  //91 / 127 = 0
    16'b01011011_10000000 : OUT <= 0;  //91 / 128 = 0
    16'b01011011_10000001 : OUT <= 0;  //91 / 129 = 0
    16'b01011011_10000010 : OUT <= 0;  //91 / 130 = 0
    16'b01011011_10000011 : OUT <= 0;  //91 / 131 = 0
    16'b01011011_10000100 : OUT <= 0;  //91 / 132 = 0
    16'b01011011_10000101 : OUT <= 0;  //91 / 133 = 0
    16'b01011011_10000110 : OUT <= 0;  //91 / 134 = 0
    16'b01011011_10000111 : OUT <= 0;  //91 / 135 = 0
    16'b01011011_10001000 : OUT <= 0;  //91 / 136 = 0
    16'b01011011_10001001 : OUT <= 0;  //91 / 137 = 0
    16'b01011011_10001010 : OUT <= 0;  //91 / 138 = 0
    16'b01011011_10001011 : OUT <= 0;  //91 / 139 = 0
    16'b01011011_10001100 : OUT <= 0;  //91 / 140 = 0
    16'b01011011_10001101 : OUT <= 0;  //91 / 141 = 0
    16'b01011011_10001110 : OUT <= 0;  //91 / 142 = 0
    16'b01011011_10001111 : OUT <= 0;  //91 / 143 = 0
    16'b01011011_10010000 : OUT <= 0;  //91 / 144 = 0
    16'b01011011_10010001 : OUT <= 0;  //91 / 145 = 0
    16'b01011011_10010010 : OUT <= 0;  //91 / 146 = 0
    16'b01011011_10010011 : OUT <= 0;  //91 / 147 = 0
    16'b01011011_10010100 : OUT <= 0;  //91 / 148 = 0
    16'b01011011_10010101 : OUT <= 0;  //91 / 149 = 0
    16'b01011011_10010110 : OUT <= 0;  //91 / 150 = 0
    16'b01011011_10010111 : OUT <= 0;  //91 / 151 = 0
    16'b01011011_10011000 : OUT <= 0;  //91 / 152 = 0
    16'b01011011_10011001 : OUT <= 0;  //91 / 153 = 0
    16'b01011011_10011010 : OUT <= 0;  //91 / 154 = 0
    16'b01011011_10011011 : OUT <= 0;  //91 / 155 = 0
    16'b01011011_10011100 : OUT <= 0;  //91 / 156 = 0
    16'b01011011_10011101 : OUT <= 0;  //91 / 157 = 0
    16'b01011011_10011110 : OUT <= 0;  //91 / 158 = 0
    16'b01011011_10011111 : OUT <= 0;  //91 / 159 = 0
    16'b01011011_10100000 : OUT <= 0;  //91 / 160 = 0
    16'b01011011_10100001 : OUT <= 0;  //91 / 161 = 0
    16'b01011011_10100010 : OUT <= 0;  //91 / 162 = 0
    16'b01011011_10100011 : OUT <= 0;  //91 / 163 = 0
    16'b01011011_10100100 : OUT <= 0;  //91 / 164 = 0
    16'b01011011_10100101 : OUT <= 0;  //91 / 165 = 0
    16'b01011011_10100110 : OUT <= 0;  //91 / 166 = 0
    16'b01011011_10100111 : OUT <= 0;  //91 / 167 = 0
    16'b01011011_10101000 : OUT <= 0;  //91 / 168 = 0
    16'b01011011_10101001 : OUT <= 0;  //91 / 169 = 0
    16'b01011011_10101010 : OUT <= 0;  //91 / 170 = 0
    16'b01011011_10101011 : OUT <= 0;  //91 / 171 = 0
    16'b01011011_10101100 : OUT <= 0;  //91 / 172 = 0
    16'b01011011_10101101 : OUT <= 0;  //91 / 173 = 0
    16'b01011011_10101110 : OUT <= 0;  //91 / 174 = 0
    16'b01011011_10101111 : OUT <= 0;  //91 / 175 = 0
    16'b01011011_10110000 : OUT <= 0;  //91 / 176 = 0
    16'b01011011_10110001 : OUT <= 0;  //91 / 177 = 0
    16'b01011011_10110010 : OUT <= 0;  //91 / 178 = 0
    16'b01011011_10110011 : OUT <= 0;  //91 / 179 = 0
    16'b01011011_10110100 : OUT <= 0;  //91 / 180 = 0
    16'b01011011_10110101 : OUT <= 0;  //91 / 181 = 0
    16'b01011011_10110110 : OUT <= 0;  //91 / 182 = 0
    16'b01011011_10110111 : OUT <= 0;  //91 / 183 = 0
    16'b01011011_10111000 : OUT <= 0;  //91 / 184 = 0
    16'b01011011_10111001 : OUT <= 0;  //91 / 185 = 0
    16'b01011011_10111010 : OUT <= 0;  //91 / 186 = 0
    16'b01011011_10111011 : OUT <= 0;  //91 / 187 = 0
    16'b01011011_10111100 : OUT <= 0;  //91 / 188 = 0
    16'b01011011_10111101 : OUT <= 0;  //91 / 189 = 0
    16'b01011011_10111110 : OUT <= 0;  //91 / 190 = 0
    16'b01011011_10111111 : OUT <= 0;  //91 / 191 = 0
    16'b01011011_11000000 : OUT <= 0;  //91 / 192 = 0
    16'b01011011_11000001 : OUT <= 0;  //91 / 193 = 0
    16'b01011011_11000010 : OUT <= 0;  //91 / 194 = 0
    16'b01011011_11000011 : OUT <= 0;  //91 / 195 = 0
    16'b01011011_11000100 : OUT <= 0;  //91 / 196 = 0
    16'b01011011_11000101 : OUT <= 0;  //91 / 197 = 0
    16'b01011011_11000110 : OUT <= 0;  //91 / 198 = 0
    16'b01011011_11000111 : OUT <= 0;  //91 / 199 = 0
    16'b01011011_11001000 : OUT <= 0;  //91 / 200 = 0
    16'b01011011_11001001 : OUT <= 0;  //91 / 201 = 0
    16'b01011011_11001010 : OUT <= 0;  //91 / 202 = 0
    16'b01011011_11001011 : OUT <= 0;  //91 / 203 = 0
    16'b01011011_11001100 : OUT <= 0;  //91 / 204 = 0
    16'b01011011_11001101 : OUT <= 0;  //91 / 205 = 0
    16'b01011011_11001110 : OUT <= 0;  //91 / 206 = 0
    16'b01011011_11001111 : OUT <= 0;  //91 / 207 = 0
    16'b01011011_11010000 : OUT <= 0;  //91 / 208 = 0
    16'b01011011_11010001 : OUT <= 0;  //91 / 209 = 0
    16'b01011011_11010010 : OUT <= 0;  //91 / 210 = 0
    16'b01011011_11010011 : OUT <= 0;  //91 / 211 = 0
    16'b01011011_11010100 : OUT <= 0;  //91 / 212 = 0
    16'b01011011_11010101 : OUT <= 0;  //91 / 213 = 0
    16'b01011011_11010110 : OUT <= 0;  //91 / 214 = 0
    16'b01011011_11010111 : OUT <= 0;  //91 / 215 = 0
    16'b01011011_11011000 : OUT <= 0;  //91 / 216 = 0
    16'b01011011_11011001 : OUT <= 0;  //91 / 217 = 0
    16'b01011011_11011010 : OUT <= 0;  //91 / 218 = 0
    16'b01011011_11011011 : OUT <= 0;  //91 / 219 = 0
    16'b01011011_11011100 : OUT <= 0;  //91 / 220 = 0
    16'b01011011_11011101 : OUT <= 0;  //91 / 221 = 0
    16'b01011011_11011110 : OUT <= 0;  //91 / 222 = 0
    16'b01011011_11011111 : OUT <= 0;  //91 / 223 = 0
    16'b01011011_11100000 : OUT <= 0;  //91 / 224 = 0
    16'b01011011_11100001 : OUT <= 0;  //91 / 225 = 0
    16'b01011011_11100010 : OUT <= 0;  //91 / 226 = 0
    16'b01011011_11100011 : OUT <= 0;  //91 / 227 = 0
    16'b01011011_11100100 : OUT <= 0;  //91 / 228 = 0
    16'b01011011_11100101 : OUT <= 0;  //91 / 229 = 0
    16'b01011011_11100110 : OUT <= 0;  //91 / 230 = 0
    16'b01011011_11100111 : OUT <= 0;  //91 / 231 = 0
    16'b01011011_11101000 : OUT <= 0;  //91 / 232 = 0
    16'b01011011_11101001 : OUT <= 0;  //91 / 233 = 0
    16'b01011011_11101010 : OUT <= 0;  //91 / 234 = 0
    16'b01011011_11101011 : OUT <= 0;  //91 / 235 = 0
    16'b01011011_11101100 : OUT <= 0;  //91 / 236 = 0
    16'b01011011_11101101 : OUT <= 0;  //91 / 237 = 0
    16'b01011011_11101110 : OUT <= 0;  //91 / 238 = 0
    16'b01011011_11101111 : OUT <= 0;  //91 / 239 = 0
    16'b01011011_11110000 : OUT <= 0;  //91 / 240 = 0
    16'b01011011_11110001 : OUT <= 0;  //91 / 241 = 0
    16'b01011011_11110010 : OUT <= 0;  //91 / 242 = 0
    16'b01011011_11110011 : OUT <= 0;  //91 / 243 = 0
    16'b01011011_11110100 : OUT <= 0;  //91 / 244 = 0
    16'b01011011_11110101 : OUT <= 0;  //91 / 245 = 0
    16'b01011011_11110110 : OUT <= 0;  //91 / 246 = 0
    16'b01011011_11110111 : OUT <= 0;  //91 / 247 = 0
    16'b01011011_11111000 : OUT <= 0;  //91 / 248 = 0
    16'b01011011_11111001 : OUT <= 0;  //91 / 249 = 0
    16'b01011011_11111010 : OUT <= 0;  //91 / 250 = 0
    16'b01011011_11111011 : OUT <= 0;  //91 / 251 = 0
    16'b01011011_11111100 : OUT <= 0;  //91 / 252 = 0
    16'b01011011_11111101 : OUT <= 0;  //91 / 253 = 0
    16'b01011011_11111110 : OUT <= 0;  //91 / 254 = 0
    16'b01011011_11111111 : OUT <= 0;  //91 / 255 = 0
    16'b01011100_00000000 : OUT <= 0;  //92 / 0 = 0
    16'b01011100_00000001 : OUT <= 92;  //92 / 1 = 92
    16'b01011100_00000010 : OUT <= 46;  //92 / 2 = 46
    16'b01011100_00000011 : OUT <= 30;  //92 / 3 = 30
    16'b01011100_00000100 : OUT <= 23;  //92 / 4 = 23
    16'b01011100_00000101 : OUT <= 18;  //92 / 5 = 18
    16'b01011100_00000110 : OUT <= 15;  //92 / 6 = 15
    16'b01011100_00000111 : OUT <= 13;  //92 / 7 = 13
    16'b01011100_00001000 : OUT <= 11;  //92 / 8 = 11
    16'b01011100_00001001 : OUT <= 10;  //92 / 9 = 10
    16'b01011100_00001010 : OUT <= 9;  //92 / 10 = 9
    16'b01011100_00001011 : OUT <= 8;  //92 / 11 = 8
    16'b01011100_00001100 : OUT <= 7;  //92 / 12 = 7
    16'b01011100_00001101 : OUT <= 7;  //92 / 13 = 7
    16'b01011100_00001110 : OUT <= 6;  //92 / 14 = 6
    16'b01011100_00001111 : OUT <= 6;  //92 / 15 = 6
    16'b01011100_00010000 : OUT <= 5;  //92 / 16 = 5
    16'b01011100_00010001 : OUT <= 5;  //92 / 17 = 5
    16'b01011100_00010010 : OUT <= 5;  //92 / 18 = 5
    16'b01011100_00010011 : OUT <= 4;  //92 / 19 = 4
    16'b01011100_00010100 : OUT <= 4;  //92 / 20 = 4
    16'b01011100_00010101 : OUT <= 4;  //92 / 21 = 4
    16'b01011100_00010110 : OUT <= 4;  //92 / 22 = 4
    16'b01011100_00010111 : OUT <= 4;  //92 / 23 = 4
    16'b01011100_00011000 : OUT <= 3;  //92 / 24 = 3
    16'b01011100_00011001 : OUT <= 3;  //92 / 25 = 3
    16'b01011100_00011010 : OUT <= 3;  //92 / 26 = 3
    16'b01011100_00011011 : OUT <= 3;  //92 / 27 = 3
    16'b01011100_00011100 : OUT <= 3;  //92 / 28 = 3
    16'b01011100_00011101 : OUT <= 3;  //92 / 29 = 3
    16'b01011100_00011110 : OUT <= 3;  //92 / 30 = 3
    16'b01011100_00011111 : OUT <= 2;  //92 / 31 = 2
    16'b01011100_00100000 : OUT <= 2;  //92 / 32 = 2
    16'b01011100_00100001 : OUT <= 2;  //92 / 33 = 2
    16'b01011100_00100010 : OUT <= 2;  //92 / 34 = 2
    16'b01011100_00100011 : OUT <= 2;  //92 / 35 = 2
    16'b01011100_00100100 : OUT <= 2;  //92 / 36 = 2
    16'b01011100_00100101 : OUT <= 2;  //92 / 37 = 2
    16'b01011100_00100110 : OUT <= 2;  //92 / 38 = 2
    16'b01011100_00100111 : OUT <= 2;  //92 / 39 = 2
    16'b01011100_00101000 : OUT <= 2;  //92 / 40 = 2
    16'b01011100_00101001 : OUT <= 2;  //92 / 41 = 2
    16'b01011100_00101010 : OUT <= 2;  //92 / 42 = 2
    16'b01011100_00101011 : OUT <= 2;  //92 / 43 = 2
    16'b01011100_00101100 : OUT <= 2;  //92 / 44 = 2
    16'b01011100_00101101 : OUT <= 2;  //92 / 45 = 2
    16'b01011100_00101110 : OUT <= 2;  //92 / 46 = 2
    16'b01011100_00101111 : OUT <= 1;  //92 / 47 = 1
    16'b01011100_00110000 : OUT <= 1;  //92 / 48 = 1
    16'b01011100_00110001 : OUT <= 1;  //92 / 49 = 1
    16'b01011100_00110010 : OUT <= 1;  //92 / 50 = 1
    16'b01011100_00110011 : OUT <= 1;  //92 / 51 = 1
    16'b01011100_00110100 : OUT <= 1;  //92 / 52 = 1
    16'b01011100_00110101 : OUT <= 1;  //92 / 53 = 1
    16'b01011100_00110110 : OUT <= 1;  //92 / 54 = 1
    16'b01011100_00110111 : OUT <= 1;  //92 / 55 = 1
    16'b01011100_00111000 : OUT <= 1;  //92 / 56 = 1
    16'b01011100_00111001 : OUT <= 1;  //92 / 57 = 1
    16'b01011100_00111010 : OUT <= 1;  //92 / 58 = 1
    16'b01011100_00111011 : OUT <= 1;  //92 / 59 = 1
    16'b01011100_00111100 : OUT <= 1;  //92 / 60 = 1
    16'b01011100_00111101 : OUT <= 1;  //92 / 61 = 1
    16'b01011100_00111110 : OUT <= 1;  //92 / 62 = 1
    16'b01011100_00111111 : OUT <= 1;  //92 / 63 = 1
    16'b01011100_01000000 : OUT <= 1;  //92 / 64 = 1
    16'b01011100_01000001 : OUT <= 1;  //92 / 65 = 1
    16'b01011100_01000010 : OUT <= 1;  //92 / 66 = 1
    16'b01011100_01000011 : OUT <= 1;  //92 / 67 = 1
    16'b01011100_01000100 : OUT <= 1;  //92 / 68 = 1
    16'b01011100_01000101 : OUT <= 1;  //92 / 69 = 1
    16'b01011100_01000110 : OUT <= 1;  //92 / 70 = 1
    16'b01011100_01000111 : OUT <= 1;  //92 / 71 = 1
    16'b01011100_01001000 : OUT <= 1;  //92 / 72 = 1
    16'b01011100_01001001 : OUT <= 1;  //92 / 73 = 1
    16'b01011100_01001010 : OUT <= 1;  //92 / 74 = 1
    16'b01011100_01001011 : OUT <= 1;  //92 / 75 = 1
    16'b01011100_01001100 : OUT <= 1;  //92 / 76 = 1
    16'b01011100_01001101 : OUT <= 1;  //92 / 77 = 1
    16'b01011100_01001110 : OUT <= 1;  //92 / 78 = 1
    16'b01011100_01001111 : OUT <= 1;  //92 / 79 = 1
    16'b01011100_01010000 : OUT <= 1;  //92 / 80 = 1
    16'b01011100_01010001 : OUT <= 1;  //92 / 81 = 1
    16'b01011100_01010010 : OUT <= 1;  //92 / 82 = 1
    16'b01011100_01010011 : OUT <= 1;  //92 / 83 = 1
    16'b01011100_01010100 : OUT <= 1;  //92 / 84 = 1
    16'b01011100_01010101 : OUT <= 1;  //92 / 85 = 1
    16'b01011100_01010110 : OUT <= 1;  //92 / 86 = 1
    16'b01011100_01010111 : OUT <= 1;  //92 / 87 = 1
    16'b01011100_01011000 : OUT <= 1;  //92 / 88 = 1
    16'b01011100_01011001 : OUT <= 1;  //92 / 89 = 1
    16'b01011100_01011010 : OUT <= 1;  //92 / 90 = 1
    16'b01011100_01011011 : OUT <= 1;  //92 / 91 = 1
    16'b01011100_01011100 : OUT <= 1;  //92 / 92 = 1
    16'b01011100_01011101 : OUT <= 0;  //92 / 93 = 0
    16'b01011100_01011110 : OUT <= 0;  //92 / 94 = 0
    16'b01011100_01011111 : OUT <= 0;  //92 / 95 = 0
    16'b01011100_01100000 : OUT <= 0;  //92 / 96 = 0
    16'b01011100_01100001 : OUT <= 0;  //92 / 97 = 0
    16'b01011100_01100010 : OUT <= 0;  //92 / 98 = 0
    16'b01011100_01100011 : OUT <= 0;  //92 / 99 = 0
    16'b01011100_01100100 : OUT <= 0;  //92 / 100 = 0
    16'b01011100_01100101 : OUT <= 0;  //92 / 101 = 0
    16'b01011100_01100110 : OUT <= 0;  //92 / 102 = 0
    16'b01011100_01100111 : OUT <= 0;  //92 / 103 = 0
    16'b01011100_01101000 : OUT <= 0;  //92 / 104 = 0
    16'b01011100_01101001 : OUT <= 0;  //92 / 105 = 0
    16'b01011100_01101010 : OUT <= 0;  //92 / 106 = 0
    16'b01011100_01101011 : OUT <= 0;  //92 / 107 = 0
    16'b01011100_01101100 : OUT <= 0;  //92 / 108 = 0
    16'b01011100_01101101 : OUT <= 0;  //92 / 109 = 0
    16'b01011100_01101110 : OUT <= 0;  //92 / 110 = 0
    16'b01011100_01101111 : OUT <= 0;  //92 / 111 = 0
    16'b01011100_01110000 : OUT <= 0;  //92 / 112 = 0
    16'b01011100_01110001 : OUT <= 0;  //92 / 113 = 0
    16'b01011100_01110010 : OUT <= 0;  //92 / 114 = 0
    16'b01011100_01110011 : OUT <= 0;  //92 / 115 = 0
    16'b01011100_01110100 : OUT <= 0;  //92 / 116 = 0
    16'b01011100_01110101 : OUT <= 0;  //92 / 117 = 0
    16'b01011100_01110110 : OUT <= 0;  //92 / 118 = 0
    16'b01011100_01110111 : OUT <= 0;  //92 / 119 = 0
    16'b01011100_01111000 : OUT <= 0;  //92 / 120 = 0
    16'b01011100_01111001 : OUT <= 0;  //92 / 121 = 0
    16'b01011100_01111010 : OUT <= 0;  //92 / 122 = 0
    16'b01011100_01111011 : OUT <= 0;  //92 / 123 = 0
    16'b01011100_01111100 : OUT <= 0;  //92 / 124 = 0
    16'b01011100_01111101 : OUT <= 0;  //92 / 125 = 0
    16'b01011100_01111110 : OUT <= 0;  //92 / 126 = 0
    16'b01011100_01111111 : OUT <= 0;  //92 / 127 = 0
    16'b01011100_10000000 : OUT <= 0;  //92 / 128 = 0
    16'b01011100_10000001 : OUT <= 0;  //92 / 129 = 0
    16'b01011100_10000010 : OUT <= 0;  //92 / 130 = 0
    16'b01011100_10000011 : OUT <= 0;  //92 / 131 = 0
    16'b01011100_10000100 : OUT <= 0;  //92 / 132 = 0
    16'b01011100_10000101 : OUT <= 0;  //92 / 133 = 0
    16'b01011100_10000110 : OUT <= 0;  //92 / 134 = 0
    16'b01011100_10000111 : OUT <= 0;  //92 / 135 = 0
    16'b01011100_10001000 : OUT <= 0;  //92 / 136 = 0
    16'b01011100_10001001 : OUT <= 0;  //92 / 137 = 0
    16'b01011100_10001010 : OUT <= 0;  //92 / 138 = 0
    16'b01011100_10001011 : OUT <= 0;  //92 / 139 = 0
    16'b01011100_10001100 : OUT <= 0;  //92 / 140 = 0
    16'b01011100_10001101 : OUT <= 0;  //92 / 141 = 0
    16'b01011100_10001110 : OUT <= 0;  //92 / 142 = 0
    16'b01011100_10001111 : OUT <= 0;  //92 / 143 = 0
    16'b01011100_10010000 : OUT <= 0;  //92 / 144 = 0
    16'b01011100_10010001 : OUT <= 0;  //92 / 145 = 0
    16'b01011100_10010010 : OUT <= 0;  //92 / 146 = 0
    16'b01011100_10010011 : OUT <= 0;  //92 / 147 = 0
    16'b01011100_10010100 : OUT <= 0;  //92 / 148 = 0
    16'b01011100_10010101 : OUT <= 0;  //92 / 149 = 0
    16'b01011100_10010110 : OUT <= 0;  //92 / 150 = 0
    16'b01011100_10010111 : OUT <= 0;  //92 / 151 = 0
    16'b01011100_10011000 : OUT <= 0;  //92 / 152 = 0
    16'b01011100_10011001 : OUT <= 0;  //92 / 153 = 0
    16'b01011100_10011010 : OUT <= 0;  //92 / 154 = 0
    16'b01011100_10011011 : OUT <= 0;  //92 / 155 = 0
    16'b01011100_10011100 : OUT <= 0;  //92 / 156 = 0
    16'b01011100_10011101 : OUT <= 0;  //92 / 157 = 0
    16'b01011100_10011110 : OUT <= 0;  //92 / 158 = 0
    16'b01011100_10011111 : OUT <= 0;  //92 / 159 = 0
    16'b01011100_10100000 : OUT <= 0;  //92 / 160 = 0
    16'b01011100_10100001 : OUT <= 0;  //92 / 161 = 0
    16'b01011100_10100010 : OUT <= 0;  //92 / 162 = 0
    16'b01011100_10100011 : OUT <= 0;  //92 / 163 = 0
    16'b01011100_10100100 : OUT <= 0;  //92 / 164 = 0
    16'b01011100_10100101 : OUT <= 0;  //92 / 165 = 0
    16'b01011100_10100110 : OUT <= 0;  //92 / 166 = 0
    16'b01011100_10100111 : OUT <= 0;  //92 / 167 = 0
    16'b01011100_10101000 : OUT <= 0;  //92 / 168 = 0
    16'b01011100_10101001 : OUT <= 0;  //92 / 169 = 0
    16'b01011100_10101010 : OUT <= 0;  //92 / 170 = 0
    16'b01011100_10101011 : OUT <= 0;  //92 / 171 = 0
    16'b01011100_10101100 : OUT <= 0;  //92 / 172 = 0
    16'b01011100_10101101 : OUT <= 0;  //92 / 173 = 0
    16'b01011100_10101110 : OUT <= 0;  //92 / 174 = 0
    16'b01011100_10101111 : OUT <= 0;  //92 / 175 = 0
    16'b01011100_10110000 : OUT <= 0;  //92 / 176 = 0
    16'b01011100_10110001 : OUT <= 0;  //92 / 177 = 0
    16'b01011100_10110010 : OUT <= 0;  //92 / 178 = 0
    16'b01011100_10110011 : OUT <= 0;  //92 / 179 = 0
    16'b01011100_10110100 : OUT <= 0;  //92 / 180 = 0
    16'b01011100_10110101 : OUT <= 0;  //92 / 181 = 0
    16'b01011100_10110110 : OUT <= 0;  //92 / 182 = 0
    16'b01011100_10110111 : OUT <= 0;  //92 / 183 = 0
    16'b01011100_10111000 : OUT <= 0;  //92 / 184 = 0
    16'b01011100_10111001 : OUT <= 0;  //92 / 185 = 0
    16'b01011100_10111010 : OUT <= 0;  //92 / 186 = 0
    16'b01011100_10111011 : OUT <= 0;  //92 / 187 = 0
    16'b01011100_10111100 : OUT <= 0;  //92 / 188 = 0
    16'b01011100_10111101 : OUT <= 0;  //92 / 189 = 0
    16'b01011100_10111110 : OUT <= 0;  //92 / 190 = 0
    16'b01011100_10111111 : OUT <= 0;  //92 / 191 = 0
    16'b01011100_11000000 : OUT <= 0;  //92 / 192 = 0
    16'b01011100_11000001 : OUT <= 0;  //92 / 193 = 0
    16'b01011100_11000010 : OUT <= 0;  //92 / 194 = 0
    16'b01011100_11000011 : OUT <= 0;  //92 / 195 = 0
    16'b01011100_11000100 : OUT <= 0;  //92 / 196 = 0
    16'b01011100_11000101 : OUT <= 0;  //92 / 197 = 0
    16'b01011100_11000110 : OUT <= 0;  //92 / 198 = 0
    16'b01011100_11000111 : OUT <= 0;  //92 / 199 = 0
    16'b01011100_11001000 : OUT <= 0;  //92 / 200 = 0
    16'b01011100_11001001 : OUT <= 0;  //92 / 201 = 0
    16'b01011100_11001010 : OUT <= 0;  //92 / 202 = 0
    16'b01011100_11001011 : OUT <= 0;  //92 / 203 = 0
    16'b01011100_11001100 : OUT <= 0;  //92 / 204 = 0
    16'b01011100_11001101 : OUT <= 0;  //92 / 205 = 0
    16'b01011100_11001110 : OUT <= 0;  //92 / 206 = 0
    16'b01011100_11001111 : OUT <= 0;  //92 / 207 = 0
    16'b01011100_11010000 : OUT <= 0;  //92 / 208 = 0
    16'b01011100_11010001 : OUT <= 0;  //92 / 209 = 0
    16'b01011100_11010010 : OUT <= 0;  //92 / 210 = 0
    16'b01011100_11010011 : OUT <= 0;  //92 / 211 = 0
    16'b01011100_11010100 : OUT <= 0;  //92 / 212 = 0
    16'b01011100_11010101 : OUT <= 0;  //92 / 213 = 0
    16'b01011100_11010110 : OUT <= 0;  //92 / 214 = 0
    16'b01011100_11010111 : OUT <= 0;  //92 / 215 = 0
    16'b01011100_11011000 : OUT <= 0;  //92 / 216 = 0
    16'b01011100_11011001 : OUT <= 0;  //92 / 217 = 0
    16'b01011100_11011010 : OUT <= 0;  //92 / 218 = 0
    16'b01011100_11011011 : OUT <= 0;  //92 / 219 = 0
    16'b01011100_11011100 : OUT <= 0;  //92 / 220 = 0
    16'b01011100_11011101 : OUT <= 0;  //92 / 221 = 0
    16'b01011100_11011110 : OUT <= 0;  //92 / 222 = 0
    16'b01011100_11011111 : OUT <= 0;  //92 / 223 = 0
    16'b01011100_11100000 : OUT <= 0;  //92 / 224 = 0
    16'b01011100_11100001 : OUT <= 0;  //92 / 225 = 0
    16'b01011100_11100010 : OUT <= 0;  //92 / 226 = 0
    16'b01011100_11100011 : OUT <= 0;  //92 / 227 = 0
    16'b01011100_11100100 : OUT <= 0;  //92 / 228 = 0
    16'b01011100_11100101 : OUT <= 0;  //92 / 229 = 0
    16'b01011100_11100110 : OUT <= 0;  //92 / 230 = 0
    16'b01011100_11100111 : OUT <= 0;  //92 / 231 = 0
    16'b01011100_11101000 : OUT <= 0;  //92 / 232 = 0
    16'b01011100_11101001 : OUT <= 0;  //92 / 233 = 0
    16'b01011100_11101010 : OUT <= 0;  //92 / 234 = 0
    16'b01011100_11101011 : OUT <= 0;  //92 / 235 = 0
    16'b01011100_11101100 : OUT <= 0;  //92 / 236 = 0
    16'b01011100_11101101 : OUT <= 0;  //92 / 237 = 0
    16'b01011100_11101110 : OUT <= 0;  //92 / 238 = 0
    16'b01011100_11101111 : OUT <= 0;  //92 / 239 = 0
    16'b01011100_11110000 : OUT <= 0;  //92 / 240 = 0
    16'b01011100_11110001 : OUT <= 0;  //92 / 241 = 0
    16'b01011100_11110010 : OUT <= 0;  //92 / 242 = 0
    16'b01011100_11110011 : OUT <= 0;  //92 / 243 = 0
    16'b01011100_11110100 : OUT <= 0;  //92 / 244 = 0
    16'b01011100_11110101 : OUT <= 0;  //92 / 245 = 0
    16'b01011100_11110110 : OUT <= 0;  //92 / 246 = 0
    16'b01011100_11110111 : OUT <= 0;  //92 / 247 = 0
    16'b01011100_11111000 : OUT <= 0;  //92 / 248 = 0
    16'b01011100_11111001 : OUT <= 0;  //92 / 249 = 0
    16'b01011100_11111010 : OUT <= 0;  //92 / 250 = 0
    16'b01011100_11111011 : OUT <= 0;  //92 / 251 = 0
    16'b01011100_11111100 : OUT <= 0;  //92 / 252 = 0
    16'b01011100_11111101 : OUT <= 0;  //92 / 253 = 0
    16'b01011100_11111110 : OUT <= 0;  //92 / 254 = 0
    16'b01011100_11111111 : OUT <= 0;  //92 / 255 = 0
    16'b01011101_00000000 : OUT <= 0;  //93 / 0 = 0
    16'b01011101_00000001 : OUT <= 93;  //93 / 1 = 93
    16'b01011101_00000010 : OUT <= 46;  //93 / 2 = 46
    16'b01011101_00000011 : OUT <= 31;  //93 / 3 = 31
    16'b01011101_00000100 : OUT <= 23;  //93 / 4 = 23
    16'b01011101_00000101 : OUT <= 18;  //93 / 5 = 18
    16'b01011101_00000110 : OUT <= 15;  //93 / 6 = 15
    16'b01011101_00000111 : OUT <= 13;  //93 / 7 = 13
    16'b01011101_00001000 : OUT <= 11;  //93 / 8 = 11
    16'b01011101_00001001 : OUT <= 10;  //93 / 9 = 10
    16'b01011101_00001010 : OUT <= 9;  //93 / 10 = 9
    16'b01011101_00001011 : OUT <= 8;  //93 / 11 = 8
    16'b01011101_00001100 : OUT <= 7;  //93 / 12 = 7
    16'b01011101_00001101 : OUT <= 7;  //93 / 13 = 7
    16'b01011101_00001110 : OUT <= 6;  //93 / 14 = 6
    16'b01011101_00001111 : OUT <= 6;  //93 / 15 = 6
    16'b01011101_00010000 : OUT <= 5;  //93 / 16 = 5
    16'b01011101_00010001 : OUT <= 5;  //93 / 17 = 5
    16'b01011101_00010010 : OUT <= 5;  //93 / 18 = 5
    16'b01011101_00010011 : OUT <= 4;  //93 / 19 = 4
    16'b01011101_00010100 : OUT <= 4;  //93 / 20 = 4
    16'b01011101_00010101 : OUT <= 4;  //93 / 21 = 4
    16'b01011101_00010110 : OUT <= 4;  //93 / 22 = 4
    16'b01011101_00010111 : OUT <= 4;  //93 / 23 = 4
    16'b01011101_00011000 : OUT <= 3;  //93 / 24 = 3
    16'b01011101_00011001 : OUT <= 3;  //93 / 25 = 3
    16'b01011101_00011010 : OUT <= 3;  //93 / 26 = 3
    16'b01011101_00011011 : OUT <= 3;  //93 / 27 = 3
    16'b01011101_00011100 : OUT <= 3;  //93 / 28 = 3
    16'b01011101_00011101 : OUT <= 3;  //93 / 29 = 3
    16'b01011101_00011110 : OUT <= 3;  //93 / 30 = 3
    16'b01011101_00011111 : OUT <= 3;  //93 / 31 = 3
    16'b01011101_00100000 : OUT <= 2;  //93 / 32 = 2
    16'b01011101_00100001 : OUT <= 2;  //93 / 33 = 2
    16'b01011101_00100010 : OUT <= 2;  //93 / 34 = 2
    16'b01011101_00100011 : OUT <= 2;  //93 / 35 = 2
    16'b01011101_00100100 : OUT <= 2;  //93 / 36 = 2
    16'b01011101_00100101 : OUT <= 2;  //93 / 37 = 2
    16'b01011101_00100110 : OUT <= 2;  //93 / 38 = 2
    16'b01011101_00100111 : OUT <= 2;  //93 / 39 = 2
    16'b01011101_00101000 : OUT <= 2;  //93 / 40 = 2
    16'b01011101_00101001 : OUT <= 2;  //93 / 41 = 2
    16'b01011101_00101010 : OUT <= 2;  //93 / 42 = 2
    16'b01011101_00101011 : OUT <= 2;  //93 / 43 = 2
    16'b01011101_00101100 : OUT <= 2;  //93 / 44 = 2
    16'b01011101_00101101 : OUT <= 2;  //93 / 45 = 2
    16'b01011101_00101110 : OUT <= 2;  //93 / 46 = 2
    16'b01011101_00101111 : OUT <= 1;  //93 / 47 = 1
    16'b01011101_00110000 : OUT <= 1;  //93 / 48 = 1
    16'b01011101_00110001 : OUT <= 1;  //93 / 49 = 1
    16'b01011101_00110010 : OUT <= 1;  //93 / 50 = 1
    16'b01011101_00110011 : OUT <= 1;  //93 / 51 = 1
    16'b01011101_00110100 : OUT <= 1;  //93 / 52 = 1
    16'b01011101_00110101 : OUT <= 1;  //93 / 53 = 1
    16'b01011101_00110110 : OUT <= 1;  //93 / 54 = 1
    16'b01011101_00110111 : OUT <= 1;  //93 / 55 = 1
    16'b01011101_00111000 : OUT <= 1;  //93 / 56 = 1
    16'b01011101_00111001 : OUT <= 1;  //93 / 57 = 1
    16'b01011101_00111010 : OUT <= 1;  //93 / 58 = 1
    16'b01011101_00111011 : OUT <= 1;  //93 / 59 = 1
    16'b01011101_00111100 : OUT <= 1;  //93 / 60 = 1
    16'b01011101_00111101 : OUT <= 1;  //93 / 61 = 1
    16'b01011101_00111110 : OUT <= 1;  //93 / 62 = 1
    16'b01011101_00111111 : OUT <= 1;  //93 / 63 = 1
    16'b01011101_01000000 : OUT <= 1;  //93 / 64 = 1
    16'b01011101_01000001 : OUT <= 1;  //93 / 65 = 1
    16'b01011101_01000010 : OUT <= 1;  //93 / 66 = 1
    16'b01011101_01000011 : OUT <= 1;  //93 / 67 = 1
    16'b01011101_01000100 : OUT <= 1;  //93 / 68 = 1
    16'b01011101_01000101 : OUT <= 1;  //93 / 69 = 1
    16'b01011101_01000110 : OUT <= 1;  //93 / 70 = 1
    16'b01011101_01000111 : OUT <= 1;  //93 / 71 = 1
    16'b01011101_01001000 : OUT <= 1;  //93 / 72 = 1
    16'b01011101_01001001 : OUT <= 1;  //93 / 73 = 1
    16'b01011101_01001010 : OUT <= 1;  //93 / 74 = 1
    16'b01011101_01001011 : OUT <= 1;  //93 / 75 = 1
    16'b01011101_01001100 : OUT <= 1;  //93 / 76 = 1
    16'b01011101_01001101 : OUT <= 1;  //93 / 77 = 1
    16'b01011101_01001110 : OUT <= 1;  //93 / 78 = 1
    16'b01011101_01001111 : OUT <= 1;  //93 / 79 = 1
    16'b01011101_01010000 : OUT <= 1;  //93 / 80 = 1
    16'b01011101_01010001 : OUT <= 1;  //93 / 81 = 1
    16'b01011101_01010010 : OUT <= 1;  //93 / 82 = 1
    16'b01011101_01010011 : OUT <= 1;  //93 / 83 = 1
    16'b01011101_01010100 : OUT <= 1;  //93 / 84 = 1
    16'b01011101_01010101 : OUT <= 1;  //93 / 85 = 1
    16'b01011101_01010110 : OUT <= 1;  //93 / 86 = 1
    16'b01011101_01010111 : OUT <= 1;  //93 / 87 = 1
    16'b01011101_01011000 : OUT <= 1;  //93 / 88 = 1
    16'b01011101_01011001 : OUT <= 1;  //93 / 89 = 1
    16'b01011101_01011010 : OUT <= 1;  //93 / 90 = 1
    16'b01011101_01011011 : OUT <= 1;  //93 / 91 = 1
    16'b01011101_01011100 : OUT <= 1;  //93 / 92 = 1
    16'b01011101_01011101 : OUT <= 1;  //93 / 93 = 1
    16'b01011101_01011110 : OUT <= 0;  //93 / 94 = 0
    16'b01011101_01011111 : OUT <= 0;  //93 / 95 = 0
    16'b01011101_01100000 : OUT <= 0;  //93 / 96 = 0
    16'b01011101_01100001 : OUT <= 0;  //93 / 97 = 0
    16'b01011101_01100010 : OUT <= 0;  //93 / 98 = 0
    16'b01011101_01100011 : OUT <= 0;  //93 / 99 = 0
    16'b01011101_01100100 : OUT <= 0;  //93 / 100 = 0
    16'b01011101_01100101 : OUT <= 0;  //93 / 101 = 0
    16'b01011101_01100110 : OUT <= 0;  //93 / 102 = 0
    16'b01011101_01100111 : OUT <= 0;  //93 / 103 = 0
    16'b01011101_01101000 : OUT <= 0;  //93 / 104 = 0
    16'b01011101_01101001 : OUT <= 0;  //93 / 105 = 0
    16'b01011101_01101010 : OUT <= 0;  //93 / 106 = 0
    16'b01011101_01101011 : OUT <= 0;  //93 / 107 = 0
    16'b01011101_01101100 : OUT <= 0;  //93 / 108 = 0
    16'b01011101_01101101 : OUT <= 0;  //93 / 109 = 0
    16'b01011101_01101110 : OUT <= 0;  //93 / 110 = 0
    16'b01011101_01101111 : OUT <= 0;  //93 / 111 = 0
    16'b01011101_01110000 : OUT <= 0;  //93 / 112 = 0
    16'b01011101_01110001 : OUT <= 0;  //93 / 113 = 0
    16'b01011101_01110010 : OUT <= 0;  //93 / 114 = 0
    16'b01011101_01110011 : OUT <= 0;  //93 / 115 = 0
    16'b01011101_01110100 : OUT <= 0;  //93 / 116 = 0
    16'b01011101_01110101 : OUT <= 0;  //93 / 117 = 0
    16'b01011101_01110110 : OUT <= 0;  //93 / 118 = 0
    16'b01011101_01110111 : OUT <= 0;  //93 / 119 = 0
    16'b01011101_01111000 : OUT <= 0;  //93 / 120 = 0
    16'b01011101_01111001 : OUT <= 0;  //93 / 121 = 0
    16'b01011101_01111010 : OUT <= 0;  //93 / 122 = 0
    16'b01011101_01111011 : OUT <= 0;  //93 / 123 = 0
    16'b01011101_01111100 : OUT <= 0;  //93 / 124 = 0
    16'b01011101_01111101 : OUT <= 0;  //93 / 125 = 0
    16'b01011101_01111110 : OUT <= 0;  //93 / 126 = 0
    16'b01011101_01111111 : OUT <= 0;  //93 / 127 = 0
    16'b01011101_10000000 : OUT <= 0;  //93 / 128 = 0
    16'b01011101_10000001 : OUT <= 0;  //93 / 129 = 0
    16'b01011101_10000010 : OUT <= 0;  //93 / 130 = 0
    16'b01011101_10000011 : OUT <= 0;  //93 / 131 = 0
    16'b01011101_10000100 : OUT <= 0;  //93 / 132 = 0
    16'b01011101_10000101 : OUT <= 0;  //93 / 133 = 0
    16'b01011101_10000110 : OUT <= 0;  //93 / 134 = 0
    16'b01011101_10000111 : OUT <= 0;  //93 / 135 = 0
    16'b01011101_10001000 : OUT <= 0;  //93 / 136 = 0
    16'b01011101_10001001 : OUT <= 0;  //93 / 137 = 0
    16'b01011101_10001010 : OUT <= 0;  //93 / 138 = 0
    16'b01011101_10001011 : OUT <= 0;  //93 / 139 = 0
    16'b01011101_10001100 : OUT <= 0;  //93 / 140 = 0
    16'b01011101_10001101 : OUT <= 0;  //93 / 141 = 0
    16'b01011101_10001110 : OUT <= 0;  //93 / 142 = 0
    16'b01011101_10001111 : OUT <= 0;  //93 / 143 = 0
    16'b01011101_10010000 : OUT <= 0;  //93 / 144 = 0
    16'b01011101_10010001 : OUT <= 0;  //93 / 145 = 0
    16'b01011101_10010010 : OUT <= 0;  //93 / 146 = 0
    16'b01011101_10010011 : OUT <= 0;  //93 / 147 = 0
    16'b01011101_10010100 : OUT <= 0;  //93 / 148 = 0
    16'b01011101_10010101 : OUT <= 0;  //93 / 149 = 0
    16'b01011101_10010110 : OUT <= 0;  //93 / 150 = 0
    16'b01011101_10010111 : OUT <= 0;  //93 / 151 = 0
    16'b01011101_10011000 : OUT <= 0;  //93 / 152 = 0
    16'b01011101_10011001 : OUT <= 0;  //93 / 153 = 0
    16'b01011101_10011010 : OUT <= 0;  //93 / 154 = 0
    16'b01011101_10011011 : OUT <= 0;  //93 / 155 = 0
    16'b01011101_10011100 : OUT <= 0;  //93 / 156 = 0
    16'b01011101_10011101 : OUT <= 0;  //93 / 157 = 0
    16'b01011101_10011110 : OUT <= 0;  //93 / 158 = 0
    16'b01011101_10011111 : OUT <= 0;  //93 / 159 = 0
    16'b01011101_10100000 : OUT <= 0;  //93 / 160 = 0
    16'b01011101_10100001 : OUT <= 0;  //93 / 161 = 0
    16'b01011101_10100010 : OUT <= 0;  //93 / 162 = 0
    16'b01011101_10100011 : OUT <= 0;  //93 / 163 = 0
    16'b01011101_10100100 : OUT <= 0;  //93 / 164 = 0
    16'b01011101_10100101 : OUT <= 0;  //93 / 165 = 0
    16'b01011101_10100110 : OUT <= 0;  //93 / 166 = 0
    16'b01011101_10100111 : OUT <= 0;  //93 / 167 = 0
    16'b01011101_10101000 : OUT <= 0;  //93 / 168 = 0
    16'b01011101_10101001 : OUT <= 0;  //93 / 169 = 0
    16'b01011101_10101010 : OUT <= 0;  //93 / 170 = 0
    16'b01011101_10101011 : OUT <= 0;  //93 / 171 = 0
    16'b01011101_10101100 : OUT <= 0;  //93 / 172 = 0
    16'b01011101_10101101 : OUT <= 0;  //93 / 173 = 0
    16'b01011101_10101110 : OUT <= 0;  //93 / 174 = 0
    16'b01011101_10101111 : OUT <= 0;  //93 / 175 = 0
    16'b01011101_10110000 : OUT <= 0;  //93 / 176 = 0
    16'b01011101_10110001 : OUT <= 0;  //93 / 177 = 0
    16'b01011101_10110010 : OUT <= 0;  //93 / 178 = 0
    16'b01011101_10110011 : OUT <= 0;  //93 / 179 = 0
    16'b01011101_10110100 : OUT <= 0;  //93 / 180 = 0
    16'b01011101_10110101 : OUT <= 0;  //93 / 181 = 0
    16'b01011101_10110110 : OUT <= 0;  //93 / 182 = 0
    16'b01011101_10110111 : OUT <= 0;  //93 / 183 = 0
    16'b01011101_10111000 : OUT <= 0;  //93 / 184 = 0
    16'b01011101_10111001 : OUT <= 0;  //93 / 185 = 0
    16'b01011101_10111010 : OUT <= 0;  //93 / 186 = 0
    16'b01011101_10111011 : OUT <= 0;  //93 / 187 = 0
    16'b01011101_10111100 : OUT <= 0;  //93 / 188 = 0
    16'b01011101_10111101 : OUT <= 0;  //93 / 189 = 0
    16'b01011101_10111110 : OUT <= 0;  //93 / 190 = 0
    16'b01011101_10111111 : OUT <= 0;  //93 / 191 = 0
    16'b01011101_11000000 : OUT <= 0;  //93 / 192 = 0
    16'b01011101_11000001 : OUT <= 0;  //93 / 193 = 0
    16'b01011101_11000010 : OUT <= 0;  //93 / 194 = 0
    16'b01011101_11000011 : OUT <= 0;  //93 / 195 = 0
    16'b01011101_11000100 : OUT <= 0;  //93 / 196 = 0
    16'b01011101_11000101 : OUT <= 0;  //93 / 197 = 0
    16'b01011101_11000110 : OUT <= 0;  //93 / 198 = 0
    16'b01011101_11000111 : OUT <= 0;  //93 / 199 = 0
    16'b01011101_11001000 : OUT <= 0;  //93 / 200 = 0
    16'b01011101_11001001 : OUT <= 0;  //93 / 201 = 0
    16'b01011101_11001010 : OUT <= 0;  //93 / 202 = 0
    16'b01011101_11001011 : OUT <= 0;  //93 / 203 = 0
    16'b01011101_11001100 : OUT <= 0;  //93 / 204 = 0
    16'b01011101_11001101 : OUT <= 0;  //93 / 205 = 0
    16'b01011101_11001110 : OUT <= 0;  //93 / 206 = 0
    16'b01011101_11001111 : OUT <= 0;  //93 / 207 = 0
    16'b01011101_11010000 : OUT <= 0;  //93 / 208 = 0
    16'b01011101_11010001 : OUT <= 0;  //93 / 209 = 0
    16'b01011101_11010010 : OUT <= 0;  //93 / 210 = 0
    16'b01011101_11010011 : OUT <= 0;  //93 / 211 = 0
    16'b01011101_11010100 : OUT <= 0;  //93 / 212 = 0
    16'b01011101_11010101 : OUT <= 0;  //93 / 213 = 0
    16'b01011101_11010110 : OUT <= 0;  //93 / 214 = 0
    16'b01011101_11010111 : OUT <= 0;  //93 / 215 = 0
    16'b01011101_11011000 : OUT <= 0;  //93 / 216 = 0
    16'b01011101_11011001 : OUT <= 0;  //93 / 217 = 0
    16'b01011101_11011010 : OUT <= 0;  //93 / 218 = 0
    16'b01011101_11011011 : OUT <= 0;  //93 / 219 = 0
    16'b01011101_11011100 : OUT <= 0;  //93 / 220 = 0
    16'b01011101_11011101 : OUT <= 0;  //93 / 221 = 0
    16'b01011101_11011110 : OUT <= 0;  //93 / 222 = 0
    16'b01011101_11011111 : OUT <= 0;  //93 / 223 = 0
    16'b01011101_11100000 : OUT <= 0;  //93 / 224 = 0
    16'b01011101_11100001 : OUT <= 0;  //93 / 225 = 0
    16'b01011101_11100010 : OUT <= 0;  //93 / 226 = 0
    16'b01011101_11100011 : OUT <= 0;  //93 / 227 = 0
    16'b01011101_11100100 : OUT <= 0;  //93 / 228 = 0
    16'b01011101_11100101 : OUT <= 0;  //93 / 229 = 0
    16'b01011101_11100110 : OUT <= 0;  //93 / 230 = 0
    16'b01011101_11100111 : OUT <= 0;  //93 / 231 = 0
    16'b01011101_11101000 : OUT <= 0;  //93 / 232 = 0
    16'b01011101_11101001 : OUT <= 0;  //93 / 233 = 0
    16'b01011101_11101010 : OUT <= 0;  //93 / 234 = 0
    16'b01011101_11101011 : OUT <= 0;  //93 / 235 = 0
    16'b01011101_11101100 : OUT <= 0;  //93 / 236 = 0
    16'b01011101_11101101 : OUT <= 0;  //93 / 237 = 0
    16'b01011101_11101110 : OUT <= 0;  //93 / 238 = 0
    16'b01011101_11101111 : OUT <= 0;  //93 / 239 = 0
    16'b01011101_11110000 : OUT <= 0;  //93 / 240 = 0
    16'b01011101_11110001 : OUT <= 0;  //93 / 241 = 0
    16'b01011101_11110010 : OUT <= 0;  //93 / 242 = 0
    16'b01011101_11110011 : OUT <= 0;  //93 / 243 = 0
    16'b01011101_11110100 : OUT <= 0;  //93 / 244 = 0
    16'b01011101_11110101 : OUT <= 0;  //93 / 245 = 0
    16'b01011101_11110110 : OUT <= 0;  //93 / 246 = 0
    16'b01011101_11110111 : OUT <= 0;  //93 / 247 = 0
    16'b01011101_11111000 : OUT <= 0;  //93 / 248 = 0
    16'b01011101_11111001 : OUT <= 0;  //93 / 249 = 0
    16'b01011101_11111010 : OUT <= 0;  //93 / 250 = 0
    16'b01011101_11111011 : OUT <= 0;  //93 / 251 = 0
    16'b01011101_11111100 : OUT <= 0;  //93 / 252 = 0
    16'b01011101_11111101 : OUT <= 0;  //93 / 253 = 0
    16'b01011101_11111110 : OUT <= 0;  //93 / 254 = 0
    16'b01011101_11111111 : OUT <= 0;  //93 / 255 = 0
    16'b01011110_00000000 : OUT <= 0;  //94 / 0 = 0
    16'b01011110_00000001 : OUT <= 94;  //94 / 1 = 94
    16'b01011110_00000010 : OUT <= 47;  //94 / 2 = 47
    16'b01011110_00000011 : OUT <= 31;  //94 / 3 = 31
    16'b01011110_00000100 : OUT <= 23;  //94 / 4 = 23
    16'b01011110_00000101 : OUT <= 18;  //94 / 5 = 18
    16'b01011110_00000110 : OUT <= 15;  //94 / 6 = 15
    16'b01011110_00000111 : OUT <= 13;  //94 / 7 = 13
    16'b01011110_00001000 : OUT <= 11;  //94 / 8 = 11
    16'b01011110_00001001 : OUT <= 10;  //94 / 9 = 10
    16'b01011110_00001010 : OUT <= 9;  //94 / 10 = 9
    16'b01011110_00001011 : OUT <= 8;  //94 / 11 = 8
    16'b01011110_00001100 : OUT <= 7;  //94 / 12 = 7
    16'b01011110_00001101 : OUT <= 7;  //94 / 13 = 7
    16'b01011110_00001110 : OUT <= 6;  //94 / 14 = 6
    16'b01011110_00001111 : OUT <= 6;  //94 / 15 = 6
    16'b01011110_00010000 : OUT <= 5;  //94 / 16 = 5
    16'b01011110_00010001 : OUT <= 5;  //94 / 17 = 5
    16'b01011110_00010010 : OUT <= 5;  //94 / 18 = 5
    16'b01011110_00010011 : OUT <= 4;  //94 / 19 = 4
    16'b01011110_00010100 : OUT <= 4;  //94 / 20 = 4
    16'b01011110_00010101 : OUT <= 4;  //94 / 21 = 4
    16'b01011110_00010110 : OUT <= 4;  //94 / 22 = 4
    16'b01011110_00010111 : OUT <= 4;  //94 / 23 = 4
    16'b01011110_00011000 : OUT <= 3;  //94 / 24 = 3
    16'b01011110_00011001 : OUT <= 3;  //94 / 25 = 3
    16'b01011110_00011010 : OUT <= 3;  //94 / 26 = 3
    16'b01011110_00011011 : OUT <= 3;  //94 / 27 = 3
    16'b01011110_00011100 : OUT <= 3;  //94 / 28 = 3
    16'b01011110_00011101 : OUT <= 3;  //94 / 29 = 3
    16'b01011110_00011110 : OUT <= 3;  //94 / 30 = 3
    16'b01011110_00011111 : OUT <= 3;  //94 / 31 = 3
    16'b01011110_00100000 : OUT <= 2;  //94 / 32 = 2
    16'b01011110_00100001 : OUT <= 2;  //94 / 33 = 2
    16'b01011110_00100010 : OUT <= 2;  //94 / 34 = 2
    16'b01011110_00100011 : OUT <= 2;  //94 / 35 = 2
    16'b01011110_00100100 : OUT <= 2;  //94 / 36 = 2
    16'b01011110_00100101 : OUT <= 2;  //94 / 37 = 2
    16'b01011110_00100110 : OUT <= 2;  //94 / 38 = 2
    16'b01011110_00100111 : OUT <= 2;  //94 / 39 = 2
    16'b01011110_00101000 : OUT <= 2;  //94 / 40 = 2
    16'b01011110_00101001 : OUT <= 2;  //94 / 41 = 2
    16'b01011110_00101010 : OUT <= 2;  //94 / 42 = 2
    16'b01011110_00101011 : OUT <= 2;  //94 / 43 = 2
    16'b01011110_00101100 : OUT <= 2;  //94 / 44 = 2
    16'b01011110_00101101 : OUT <= 2;  //94 / 45 = 2
    16'b01011110_00101110 : OUT <= 2;  //94 / 46 = 2
    16'b01011110_00101111 : OUT <= 2;  //94 / 47 = 2
    16'b01011110_00110000 : OUT <= 1;  //94 / 48 = 1
    16'b01011110_00110001 : OUT <= 1;  //94 / 49 = 1
    16'b01011110_00110010 : OUT <= 1;  //94 / 50 = 1
    16'b01011110_00110011 : OUT <= 1;  //94 / 51 = 1
    16'b01011110_00110100 : OUT <= 1;  //94 / 52 = 1
    16'b01011110_00110101 : OUT <= 1;  //94 / 53 = 1
    16'b01011110_00110110 : OUT <= 1;  //94 / 54 = 1
    16'b01011110_00110111 : OUT <= 1;  //94 / 55 = 1
    16'b01011110_00111000 : OUT <= 1;  //94 / 56 = 1
    16'b01011110_00111001 : OUT <= 1;  //94 / 57 = 1
    16'b01011110_00111010 : OUT <= 1;  //94 / 58 = 1
    16'b01011110_00111011 : OUT <= 1;  //94 / 59 = 1
    16'b01011110_00111100 : OUT <= 1;  //94 / 60 = 1
    16'b01011110_00111101 : OUT <= 1;  //94 / 61 = 1
    16'b01011110_00111110 : OUT <= 1;  //94 / 62 = 1
    16'b01011110_00111111 : OUT <= 1;  //94 / 63 = 1
    16'b01011110_01000000 : OUT <= 1;  //94 / 64 = 1
    16'b01011110_01000001 : OUT <= 1;  //94 / 65 = 1
    16'b01011110_01000010 : OUT <= 1;  //94 / 66 = 1
    16'b01011110_01000011 : OUT <= 1;  //94 / 67 = 1
    16'b01011110_01000100 : OUT <= 1;  //94 / 68 = 1
    16'b01011110_01000101 : OUT <= 1;  //94 / 69 = 1
    16'b01011110_01000110 : OUT <= 1;  //94 / 70 = 1
    16'b01011110_01000111 : OUT <= 1;  //94 / 71 = 1
    16'b01011110_01001000 : OUT <= 1;  //94 / 72 = 1
    16'b01011110_01001001 : OUT <= 1;  //94 / 73 = 1
    16'b01011110_01001010 : OUT <= 1;  //94 / 74 = 1
    16'b01011110_01001011 : OUT <= 1;  //94 / 75 = 1
    16'b01011110_01001100 : OUT <= 1;  //94 / 76 = 1
    16'b01011110_01001101 : OUT <= 1;  //94 / 77 = 1
    16'b01011110_01001110 : OUT <= 1;  //94 / 78 = 1
    16'b01011110_01001111 : OUT <= 1;  //94 / 79 = 1
    16'b01011110_01010000 : OUT <= 1;  //94 / 80 = 1
    16'b01011110_01010001 : OUT <= 1;  //94 / 81 = 1
    16'b01011110_01010010 : OUT <= 1;  //94 / 82 = 1
    16'b01011110_01010011 : OUT <= 1;  //94 / 83 = 1
    16'b01011110_01010100 : OUT <= 1;  //94 / 84 = 1
    16'b01011110_01010101 : OUT <= 1;  //94 / 85 = 1
    16'b01011110_01010110 : OUT <= 1;  //94 / 86 = 1
    16'b01011110_01010111 : OUT <= 1;  //94 / 87 = 1
    16'b01011110_01011000 : OUT <= 1;  //94 / 88 = 1
    16'b01011110_01011001 : OUT <= 1;  //94 / 89 = 1
    16'b01011110_01011010 : OUT <= 1;  //94 / 90 = 1
    16'b01011110_01011011 : OUT <= 1;  //94 / 91 = 1
    16'b01011110_01011100 : OUT <= 1;  //94 / 92 = 1
    16'b01011110_01011101 : OUT <= 1;  //94 / 93 = 1
    16'b01011110_01011110 : OUT <= 1;  //94 / 94 = 1
    16'b01011110_01011111 : OUT <= 0;  //94 / 95 = 0
    16'b01011110_01100000 : OUT <= 0;  //94 / 96 = 0
    16'b01011110_01100001 : OUT <= 0;  //94 / 97 = 0
    16'b01011110_01100010 : OUT <= 0;  //94 / 98 = 0
    16'b01011110_01100011 : OUT <= 0;  //94 / 99 = 0
    16'b01011110_01100100 : OUT <= 0;  //94 / 100 = 0
    16'b01011110_01100101 : OUT <= 0;  //94 / 101 = 0
    16'b01011110_01100110 : OUT <= 0;  //94 / 102 = 0
    16'b01011110_01100111 : OUT <= 0;  //94 / 103 = 0
    16'b01011110_01101000 : OUT <= 0;  //94 / 104 = 0
    16'b01011110_01101001 : OUT <= 0;  //94 / 105 = 0
    16'b01011110_01101010 : OUT <= 0;  //94 / 106 = 0
    16'b01011110_01101011 : OUT <= 0;  //94 / 107 = 0
    16'b01011110_01101100 : OUT <= 0;  //94 / 108 = 0
    16'b01011110_01101101 : OUT <= 0;  //94 / 109 = 0
    16'b01011110_01101110 : OUT <= 0;  //94 / 110 = 0
    16'b01011110_01101111 : OUT <= 0;  //94 / 111 = 0
    16'b01011110_01110000 : OUT <= 0;  //94 / 112 = 0
    16'b01011110_01110001 : OUT <= 0;  //94 / 113 = 0
    16'b01011110_01110010 : OUT <= 0;  //94 / 114 = 0
    16'b01011110_01110011 : OUT <= 0;  //94 / 115 = 0
    16'b01011110_01110100 : OUT <= 0;  //94 / 116 = 0
    16'b01011110_01110101 : OUT <= 0;  //94 / 117 = 0
    16'b01011110_01110110 : OUT <= 0;  //94 / 118 = 0
    16'b01011110_01110111 : OUT <= 0;  //94 / 119 = 0
    16'b01011110_01111000 : OUT <= 0;  //94 / 120 = 0
    16'b01011110_01111001 : OUT <= 0;  //94 / 121 = 0
    16'b01011110_01111010 : OUT <= 0;  //94 / 122 = 0
    16'b01011110_01111011 : OUT <= 0;  //94 / 123 = 0
    16'b01011110_01111100 : OUT <= 0;  //94 / 124 = 0
    16'b01011110_01111101 : OUT <= 0;  //94 / 125 = 0
    16'b01011110_01111110 : OUT <= 0;  //94 / 126 = 0
    16'b01011110_01111111 : OUT <= 0;  //94 / 127 = 0
    16'b01011110_10000000 : OUT <= 0;  //94 / 128 = 0
    16'b01011110_10000001 : OUT <= 0;  //94 / 129 = 0
    16'b01011110_10000010 : OUT <= 0;  //94 / 130 = 0
    16'b01011110_10000011 : OUT <= 0;  //94 / 131 = 0
    16'b01011110_10000100 : OUT <= 0;  //94 / 132 = 0
    16'b01011110_10000101 : OUT <= 0;  //94 / 133 = 0
    16'b01011110_10000110 : OUT <= 0;  //94 / 134 = 0
    16'b01011110_10000111 : OUT <= 0;  //94 / 135 = 0
    16'b01011110_10001000 : OUT <= 0;  //94 / 136 = 0
    16'b01011110_10001001 : OUT <= 0;  //94 / 137 = 0
    16'b01011110_10001010 : OUT <= 0;  //94 / 138 = 0
    16'b01011110_10001011 : OUT <= 0;  //94 / 139 = 0
    16'b01011110_10001100 : OUT <= 0;  //94 / 140 = 0
    16'b01011110_10001101 : OUT <= 0;  //94 / 141 = 0
    16'b01011110_10001110 : OUT <= 0;  //94 / 142 = 0
    16'b01011110_10001111 : OUT <= 0;  //94 / 143 = 0
    16'b01011110_10010000 : OUT <= 0;  //94 / 144 = 0
    16'b01011110_10010001 : OUT <= 0;  //94 / 145 = 0
    16'b01011110_10010010 : OUT <= 0;  //94 / 146 = 0
    16'b01011110_10010011 : OUT <= 0;  //94 / 147 = 0
    16'b01011110_10010100 : OUT <= 0;  //94 / 148 = 0
    16'b01011110_10010101 : OUT <= 0;  //94 / 149 = 0
    16'b01011110_10010110 : OUT <= 0;  //94 / 150 = 0
    16'b01011110_10010111 : OUT <= 0;  //94 / 151 = 0
    16'b01011110_10011000 : OUT <= 0;  //94 / 152 = 0
    16'b01011110_10011001 : OUT <= 0;  //94 / 153 = 0
    16'b01011110_10011010 : OUT <= 0;  //94 / 154 = 0
    16'b01011110_10011011 : OUT <= 0;  //94 / 155 = 0
    16'b01011110_10011100 : OUT <= 0;  //94 / 156 = 0
    16'b01011110_10011101 : OUT <= 0;  //94 / 157 = 0
    16'b01011110_10011110 : OUT <= 0;  //94 / 158 = 0
    16'b01011110_10011111 : OUT <= 0;  //94 / 159 = 0
    16'b01011110_10100000 : OUT <= 0;  //94 / 160 = 0
    16'b01011110_10100001 : OUT <= 0;  //94 / 161 = 0
    16'b01011110_10100010 : OUT <= 0;  //94 / 162 = 0
    16'b01011110_10100011 : OUT <= 0;  //94 / 163 = 0
    16'b01011110_10100100 : OUT <= 0;  //94 / 164 = 0
    16'b01011110_10100101 : OUT <= 0;  //94 / 165 = 0
    16'b01011110_10100110 : OUT <= 0;  //94 / 166 = 0
    16'b01011110_10100111 : OUT <= 0;  //94 / 167 = 0
    16'b01011110_10101000 : OUT <= 0;  //94 / 168 = 0
    16'b01011110_10101001 : OUT <= 0;  //94 / 169 = 0
    16'b01011110_10101010 : OUT <= 0;  //94 / 170 = 0
    16'b01011110_10101011 : OUT <= 0;  //94 / 171 = 0
    16'b01011110_10101100 : OUT <= 0;  //94 / 172 = 0
    16'b01011110_10101101 : OUT <= 0;  //94 / 173 = 0
    16'b01011110_10101110 : OUT <= 0;  //94 / 174 = 0
    16'b01011110_10101111 : OUT <= 0;  //94 / 175 = 0
    16'b01011110_10110000 : OUT <= 0;  //94 / 176 = 0
    16'b01011110_10110001 : OUT <= 0;  //94 / 177 = 0
    16'b01011110_10110010 : OUT <= 0;  //94 / 178 = 0
    16'b01011110_10110011 : OUT <= 0;  //94 / 179 = 0
    16'b01011110_10110100 : OUT <= 0;  //94 / 180 = 0
    16'b01011110_10110101 : OUT <= 0;  //94 / 181 = 0
    16'b01011110_10110110 : OUT <= 0;  //94 / 182 = 0
    16'b01011110_10110111 : OUT <= 0;  //94 / 183 = 0
    16'b01011110_10111000 : OUT <= 0;  //94 / 184 = 0
    16'b01011110_10111001 : OUT <= 0;  //94 / 185 = 0
    16'b01011110_10111010 : OUT <= 0;  //94 / 186 = 0
    16'b01011110_10111011 : OUT <= 0;  //94 / 187 = 0
    16'b01011110_10111100 : OUT <= 0;  //94 / 188 = 0
    16'b01011110_10111101 : OUT <= 0;  //94 / 189 = 0
    16'b01011110_10111110 : OUT <= 0;  //94 / 190 = 0
    16'b01011110_10111111 : OUT <= 0;  //94 / 191 = 0
    16'b01011110_11000000 : OUT <= 0;  //94 / 192 = 0
    16'b01011110_11000001 : OUT <= 0;  //94 / 193 = 0
    16'b01011110_11000010 : OUT <= 0;  //94 / 194 = 0
    16'b01011110_11000011 : OUT <= 0;  //94 / 195 = 0
    16'b01011110_11000100 : OUT <= 0;  //94 / 196 = 0
    16'b01011110_11000101 : OUT <= 0;  //94 / 197 = 0
    16'b01011110_11000110 : OUT <= 0;  //94 / 198 = 0
    16'b01011110_11000111 : OUT <= 0;  //94 / 199 = 0
    16'b01011110_11001000 : OUT <= 0;  //94 / 200 = 0
    16'b01011110_11001001 : OUT <= 0;  //94 / 201 = 0
    16'b01011110_11001010 : OUT <= 0;  //94 / 202 = 0
    16'b01011110_11001011 : OUT <= 0;  //94 / 203 = 0
    16'b01011110_11001100 : OUT <= 0;  //94 / 204 = 0
    16'b01011110_11001101 : OUT <= 0;  //94 / 205 = 0
    16'b01011110_11001110 : OUT <= 0;  //94 / 206 = 0
    16'b01011110_11001111 : OUT <= 0;  //94 / 207 = 0
    16'b01011110_11010000 : OUT <= 0;  //94 / 208 = 0
    16'b01011110_11010001 : OUT <= 0;  //94 / 209 = 0
    16'b01011110_11010010 : OUT <= 0;  //94 / 210 = 0
    16'b01011110_11010011 : OUT <= 0;  //94 / 211 = 0
    16'b01011110_11010100 : OUT <= 0;  //94 / 212 = 0
    16'b01011110_11010101 : OUT <= 0;  //94 / 213 = 0
    16'b01011110_11010110 : OUT <= 0;  //94 / 214 = 0
    16'b01011110_11010111 : OUT <= 0;  //94 / 215 = 0
    16'b01011110_11011000 : OUT <= 0;  //94 / 216 = 0
    16'b01011110_11011001 : OUT <= 0;  //94 / 217 = 0
    16'b01011110_11011010 : OUT <= 0;  //94 / 218 = 0
    16'b01011110_11011011 : OUT <= 0;  //94 / 219 = 0
    16'b01011110_11011100 : OUT <= 0;  //94 / 220 = 0
    16'b01011110_11011101 : OUT <= 0;  //94 / 221 = 0
    16'b01011110_11011110 : OUT <= 0;  //94 / 222 = 0
    16'b01011110_11011111 : OUT <= 0;  //94 / 223 = 0
    16'b01011110_11100000 : OUT <= 0;  //94 / 224 = 0
    16'b01011110_11100001 : OUT <= 0;  //94 / 225 = 0
    16'b01011110_11100010 : OUT <= 0;  //94 / 226 = 0
    16'b01011110_11100011 : OUT <= 0;  //94 / 227 = 0
    16'b01011110_11100100 : OUT <= 0;  //94 / 228 = 0
    16'b01011110_11100101 : OUT <= 0;  //94 / 229 = 0
    16'b01011110_11100110 : OUT <= 0;  //94 / 230 = 0
    16'b01011110_11100111 : OUT <= 0;  //94 / 231 = 0
    16'b01011110_11101000 : OUT <= 0;  //94 / 232 = 0
    16'b01011110_11101001 : OUT <= 0;  //94 / 233 = 0
    16'b01011110_11101010 : OUT <= 0;  //94 / 234 = 0
    16'b01011110_11101011 : OUT <= 0;  //94 / 235 = 0
    16'b01011110_11101100 : OUT <= 0;  //94 / 236 = 0
    16'b01011110_11101101 : OUT <= 0;  //94 / 237 = 0
    16'b01011110_11101110 : OUT <= 0;  //94 / 238 = 0
    16'b01011110_11101111 : OUT <= 0;  //94 / 239 = 0
    16'b01011110_11110000 : OUT <= 0;  //94 / 240 = 0
    16'b01011110_11110001 : OUT <= 0;  //94 / 241 = 0
    16'b01011110_11110010 : OUT <= 0;  //94 / 242 = 0
    16'b01011110_11110011 : OUT <= 0;  //94 / 243 = 0
    16'b01011110_11110100 : OUT <= 0;  //94 / 244 = 0
    16'b01011110_11110101 : OUT <= 0;  //94 / 245 = 0
    16'b01011110_11110110 : OUT <= 0;  //94 / 246 = 0
    16'b01011110_11110111 : OUT <= 0;  //94 / 247 = 0
    16'b01011110_11111000 : OUT <= 0;  //94 / 248 = 0
    16'b01011110_11111001 : OUT <= 0;  //94 / 249 = 0
    16'b01011110_11111010 : OUT <= 0;  //94 / 250 = 0
    16'b01011110_11111011 : OUT <= 0;  //94 / 251 = 0
    16'b01011110_11111100 : OUT <= 0;  //94 / 252 = 0
    16'b01011110_11111101 : OUT <= 0;  //94 / 253 = 0
    16'b01011110_11111110 : OUT <= 0;  //94 / 254 = 0
    16'b01011110_11111111 : OUT <= 0;  //94 / 255 = 0
    16'b01011111_00000000 : OUT <= 0;  //95 / 0 = 0
    16'b01011111_00000001 : OUT <= 95;  //95 / 1 = 95
    16'b01011111_00000010 : OUT <= 47;  //95 / 2 = 47
    16'b01011111_00000011 : OUT <= 31;  //95 / 3 = 31
    16'b01011111_00000100 : OUT <= 23;  //95 / 4 = 23
    16'b01011111_00000101 : OUT <= 19;  //95 / 5 = 19
    16'b01011111_00000110 : OUT <= 15;  //95 / 6 = 15
    16'b01011111_00000111 : OUT <= 13;  //95 / 7 = 13
    16'b01011111_00001000 : OUT <= 11;  //95 / 8 = 11
    16'b01011111_00001001 : OUT <= 10;  //95 / 9 = 10
    16'b01011111_00001010 : OUT <= 9;  //95 / 10 = 9
    16'b01011111_00001011 : OUT <= 8;  //95 / 11 = 8
    16'b01011111_00001100 : OUT <= 7;  //95 / 12 = 7
    16'b01011111_00001101 : OUT <= 7;  //95 / 13 = 7
    16'b01011111_00001110 : OUT <= 6;  //95 / 14 = 6
    16'b01011111_00001111 : OUT <= 6;  //95 / 15 = 6
    16'b01011111_00010000 : OUT <= 5;  //95 / 16 = 5
    16'b01011111_00010001 : OUT <= 5;  //95 / 17 = 5
    16'b01011111_00010010 : OUT <= 5;  //95 / 18 = 5
    16'b01011111_00010011 : OUT <= 5;  //95 / 19 = 5
    16'b01011111_00010100 : OUT <= 4;  //95 / 20 = 4
    16'b01011111_00010101 : OUT <= 4;  //95 / 21 = 4
    16'b01011111_00010110 : OUT <= 4;  //95 / 22 = 4
    16'b01011111_00010111 : OUT <= 4;  //95 / 23 = 4
    16'b01011111_00011000 : OUT <= 3;  //95 / 24 = 3
    16'b01011111_00011001 : OUT <= 3;  //95 / 25 = 3
    16'b01011111_00011010 : OUT <= 3;  //95 / 26 = 3
    16'b01011111_00011011 : OUT <= 3;  //95 / 27 = 3
    16'b01011111_00011100 : OUT <= 3;  //95 / 28 = 3
    16'b01011111_00011101 : OUT <= 3;  //95 / 29 = 3
    16'b01011111_00011110 : OUT <= 3;  //95 / 30 = 3
    16'b01011111_00011111 : OUT <= 3;  //95 / 31 = 3
    16'b01011111_00100000 : OUT <= 2;  //95 / 32 = 2
    16'b01011111_00100001 : OUT <= 2;  //95 / 33 = 2
    16'b01011111_00100010 : OUT <= 2;  //95 / 34 = 2
    16'b01011111_00100011 : OUT <= 2;  //95 / 35 = 2
    16'b01011111_00100100 : OUT <= 2;  //95 / 36 = 2
    16'b01011111_00100101 : OUT <= 2;  //95 / 37 = 2
    16'b01011111_00100110 : OUT <= 2;  //95 / 38 = 2
    16'b01011111_00100111 : OUT <= 2;  //95 / 39 = 2
    16'b01011111_00101000 : OUT <= 2;  //95 / 40 = 2
    16'b01011111_00101001 : OUT <= 2;  //95 / 41 = 2
    16'b01011111_00101010 : OUT <= 2;  //95 / 42 = 2
    16'b01011111_00101011 : OUT <= 2;  //95 / 43 = 2
    16'b01011111_00101100 : OUT <= 2;  //95 / 44 = 2
    16'b01011111_00101101 : OUT <= 2;  //95 / 45 = 2
    16'b01011111_00101110 : OUT <= 2;  //95 / 46 = 2
    16'b01011111_00101111 : OUT <= 2;  //95 / 47 = 2
    16'b01011111_00110000 : OUT <= 1;  //95 / 48 = 1
    16'b01011111_00110001 : OUT <= 1;  //95 / 49 = 1
    16'b01011111_00110010 : OUT <= 1;  //95 / 50 = 1
    16'b01011111_00110011 : OUT <= 1;  //95 / 51 = 1
    16'b01011111_00110100 : OUT <= 1;  //95 / 52 = 1
    16'b01011111_00110101 : OUT <= 1;  //95 / 53 = 1
    16'b01011111_00110110 : OUT <= 1;  //95 / 54 = 1
    16'b01011111_00110111 : OUT <= 1;  //95 / 55 = 1
    16'b01011111_00111000 : OUT <= 1;  //95 / 56 = 1
    16'b01011111_00111001 : OUT <= 1;  //95 / 57 = 1
    16'b01011111_00111010 : OUT <= 1;  //95 / 58 = 1
    16'b01011111_00111011 : OUT <= 1;  //95 / 59 = 1
    16'b01011111_00111100 : OUT <= 1;  //95 / 60 = 1
    16'b01011111_00111101 : OUT <= 1;  //95 / 61 = 1
    16'b01011111_00111110 : OUT <= 1;  //95 / 62 = 1
    16'b01011111_00111111 : OUT <= 1;  //95 / 63 = 1
    16'b01011111_01000000 : OUT <= 1;  //95 / 64 = 1
    16'b01011111_01000001 : OUT <= 1;  //95 / 65 = 1
    16'b01011111_01000010 : OUT <= 1;  //95 / 66 = 1
    16'b01011111_01000011 : OUT <= 1;  //95 / 67 = 1
    16'b01011111_01000100 : OUT <= 1;  //95 / 68 = 1
    16'b01011111_01000101 : OUT <= 1;  //95 / 69 = 1
    16'b01011111_01000110 : OUT <= 1;  //95 / 70 = 1
    16'b01011111_01000111 : OUT <= 1;  //95 / 71 = 1
    16'b01011111_01001000 : OUT <= 1;  //95 / 72 = 1
    16'b01011111_01001001 : OUT <= 1;  //95 / 73 = 1
    16'b01011111_01001010 : OUT <= 1;  //95 / 74 = 1
    16'b01011111_01001011 : OUT <= 1;  //95 / 75 = 1
    16'b01011111_01001100 : OUT <= 1;  //95 / 76 = 1
    16'b01011111_01001101 : OUT <= 1;  //95 / 77 = 1
    16'b01011111_01001110 : OUT <= 1;  //95 / 78 = 1
    16'b01011111_01001111 : OUT <= 1;  //95 / 79 = 1
    16'b01011111_01010000 : OUT <= 1;  //95 / 80 = 1
    16'b01011111_01010001 : OUT <= 1;  //95 / 81 = 1
    16'b01011111_01010010 : OUT <= 1;  //95 / 82 = 1
    16'b01011111_01010011 : OUT <= 1;  //95 / 83 = 1
    16'b01011111_01010100 : OUT <= 1;  //95 / 84 = 1
    16'b01011111_01010101 : OUT <= 1;  //95 / 85 = 1
    16'b01011111_01010110 : OUT <= 1;  //95 / 86 = 1
    16'b01011111_01010111 : OUT <= 1;  //95 / 87 = 1
    16'b01011111_01011000 : OUT <= 1;  //95 / 88 = 1
    16'b01011111_01011001 : OUT <= 1;  //95 / 89 = 1
    16'b01011111_01011010 : OUT <= 1;  //95 / 90 = 1
    16'b01011111_01011011 : OUT <= 1;  //95 / 91 = 1
    16'b01011111_01011100 : OUT <= 1;  //95 / 92 = 1
    16'b01011111_01011101 : OUT <= 1;  //95 / 93 = 1
    16'b01011111_01011110 : OUT <= 1;  //95 / 94 = 1
    16'b01011111_01011111 : OUT <= 1;  //95 / 95 = 1
    16'b01011111_01100000 : OUT <= 0;  //95 / 96 = 0
    16'b01011111_01100001 : OUT <= 0;  //95 / 97 = 0
    16'b01011111_01100010 : OUT <= 0;  //95 / 98 = 0
    16'b01011111_01100011 : OUT <= 0;  //95 / 99 = 0
    16'b01011111_01100100 : OUT <= 0;  //95 / 100 = 0
    16'b01011111_01100101 : OUT <= 0;  //95 / 101 = 0
    16'b01011111_01100110 : OUT <= 0;  //95 / 102 = 0
    16'b01011111_01100111 : OUT <= 0;  //95 / 103 = 0
    16'b01011111_01101000 : OUT <= 0;  //95 / 104 = 0
    16'b01011111_01101001 : OUT <= 0;  //95 / 105 = 0
    16'b01011111_01101010 : OUT <= 0;  //95 / 106 = 0
    16'b01011111_01101011 : OUT <= 0;  //95 / 107 = 0
    16'b01011111_01101100 : OUT <= 0;  //95 / 108 = 0
    16'b01011111_01101101 : OUT <= 0;  //95 / 109 = 0
    16'b01011111_01101110 : OUT <= 0;  //95 / 110 = 0
    16'b01011111_01101111 : OUT <= 0;  //95 / 111 = 0
    16'b01011111_01110000 : OUT <= 0;  //95 / 112 = 0
    16'b01011111_01110001 : OUT <= 0;  //95 / 113 = 0
    16'b01011111_01110010 : OUT <= 0;  //95 / 114 = 0
    16'b01011111_01110011 : OUT <= 0;  //95 / 115 = 0
    16'b01011111_01110100 : OUT <= 0;  //95 / 116 = 0
    16'b01011111_01110101 : OUT <= 0;  //95 / 117 = 0
    16'b01011111_01110110 : OUT <= 0;  //95 / 118 = 0
    16'b01011111_01110111 : OUT <= 0;  //95 / 119 = 0
    16'b01011111_01111000 : OUT <= 0;  //95 / 120 = 0
    16'b01011111_01111001 : OUT <= 0;  //95 / 121 = 0
    16'b01011111_01111010 : OUT <= 0;  //95 / 122 = 0
    16'b01011111_01111011 : OUT <= 0;  //95 / 123 = 0
    16'b01011111_01111100 : OUT <= 0;  //95 / 124 = 0
    16'b01011111_01111101 : OUT <= 0;  //95 / 125 = 0
    16'b01011111_01111110 : OUT <= 0;  //95 / 126 = 0
    16'b01011111_01111111 : OUT <= 0;  //95 / 127 = 0
    16'b01011111_10000000 : OUT <= 0;  //95 / 128 = 0
    16'b01011111_10000001 : OUT <= 0;  //95 / 129 = 0
    16'b01011111_10000010 : OUT <= 0;  //95 / 130 = 0
    16'b01011111_10000011 : OUT <= 0;  //95 / 131 = 0
    16'b01011111_10000100 : OUT <= 0;  //95 / 132 = 0
    16'b01011111_10000101 : OUT <= 0;  //95 / 133 = 0
    16'b01011111_10000110 : OUT <= 0;  //95 / 134 = 0
    16'b01011111_10000111 : OUT <= 0;  //95 / 135 = 0
    16'b01011111_10001000 : OUT <= 0;  //95 / 136 = 0
    16'b01011111_10001001 : OUT <= 0;  //95 / 137 = 0
    16'b01011111_10001010 : OUT <= 0;  //95 / 138 = 0
    16'b01011111_10001011 : OUT <= 0;  //95 / 139 = 0
    16'b01011111_10001100 : OUT <= 0;  //95 / 140 = 0
    16'b01011111_10001101 : OUT <= 0;  //95 / 141 = 0
    16'b01011111_10001110 : OUT <= 0;  //95 / 142 = 0
    16'b01011111_10001111 : OUT <= 0;  //95 / 143 = 0
    16'b01011111_10010000 : OUT <= 0;  //95 / 144 = 0
    16'b01011111_10010001 : OUT <= 0;  //95 / 145 = 0
    16'b01011111_10010010 : OUT <= 0;  //95 / 146 = 0
    16'b01011111_10010011 : OUT <= 0;  //95 / 147 = 0
    16'b01011111_10010100 : OUT <= 0;  //95 / 148 = 0
    16'b01011111_10010101 : OUT <= 0;  //95 / 149 = 0
    16'b01011111_10010110 : OUT <= 0;  //95 / 150 = 0
    16'b01011111_10010111 : OUT <= 0;  //95 / 151 = 0
    16'b01011111_10011000 : OUT <= 0;  //95 / 152 = 0
    16'b01011111_10011001 : OUT <= 0;  //95 / 153 = 0
    16'b01011111_10011010 : OUT <= 0;  //95 / 154 = 0
    16'b01011111_10011011 : OUT <= 0;  //95 / 155 = 0
    16'b01011111_10011100 : OUT <= 0;  //95 / 156 = 0
    16'b01011111_10011101 : OUT <= 0;  //95 / 157 = 0
    16'b01011111_10011110 : OUT <= 0;  //95 / 158 = 0
    16'b01011111_10011111 : OUT <= 0;  //95 / 159 = 0
    16'b01011111_10100000 : OUT <= 0;  //95 / 160 = 0
    16'b01011111_10100001 : OUT <= 0;  //95 / 161 = 0
    16'b01011111_10100010 : OUT <= 0;  //95 / 162 = 0
    16'b01011111_10100011 : OUT <= 0;  //95 / 163 = 0
    16'b01011111_10100100 : OUT <= 0;  //95 / 164 = 0
    16'b01011111_10100101 : OUT <= 0;  //95 / 165 = 0
    16'b01011111_10100110 : OUT <= 0;  //95 / 166 = 0
    16'b01011111_10100111 : OUT <= 0;  //95 / 167 = 0
    16'b01011111_10101000 : OUT <= 0;  //95 / 168 = 0
    16'b01011111_10101001 : OUT <= 0;  //95 / 169 = 0
    16'b01011111_10101010 : OUT <= 0;  //95 / 170 = 0
    16'b01011111_10101011 : OUT <= 0;  //95 / 171 = 0
    16'b01011111_10101100 : OUT <= 0;  //95 / 172 = 0
    16'b01011111_10101101 : OUT <= 0;  //95 / 173 = 0
    16'b01011111_10101110 : OUT <= 0;  //95 / 174 = 0
    16'b01011111_10101111 : OUT <= 0;  //95 / 175 = 0
    16'b01011111_10110000 : OUT <= 0;  //95 / 176 = 0
    16'b01011111_10110001 : OUT <= 0;  //95 / 177 = 0
    16'b01011111_10110010 : OUT <= 0;  //95 / 178 = 0
    16'b01011111_10110011 : OUT <= 0;  //95 / 179 = 0
    16'b01011111_10110100 : OUT <= 0;  //95 / 180 = 0
    16'b01011111_10110101 : OUT <= 0;  //95 / 181 = 0
    16'b01011111_10110110 : OUT <= 0;  //95 / 182 = 0
    16'b01011111_10110111 : OUT <= 0;  //95 / 183 = 0
    16'b01011111_10111000 : OUT <= 0;  //95 / 184 = 0
    16'b01011111_10111001 : OUT <= 0;  //95 / 185 = 0
    16'b01011111_10111010 : OUT <= 0;  //95 / 186 = 0
    16'b01011111_10111011 : OUT <= 0;  //95 / 187 = 0
    16'b01011111_10111100 : OUT <= 0;  //95 / 188 = 0
    16'b01011111_10111101 : OUT <= 0;  //95 / 189 = 0
    16'b01011111_10111110 : OUT <= 0;  //95 / 190 = 0
    16'b01011111_10111111 : OUT <= 0;  //95 / 191 = 0
    16'b01011111_11000000 : OUT <= 0;  //95 / 192 = 0
    16'b01011111_11000001 : OUT <= 0;  //95 / 193 = 0
    16'b01011111_11000010 : OUT <= 0;  //95 / 194 = 0
    16'b01011111_11000011 : OUT <= 0;  //95 / 195 = 0
    16'b01011111_11000100 : OUT <= 0;  //95 / 196 = 0
    16'b01011111_11000101 : OUT <= 0;  //95 / 197 = 0
    16'b01011111_11000110 : OUT <= 0;  //95 / 198 = 0
    16'b01011111_11000111 : OUT <= 0;  //95 / 199 = 0
    16'b01011111_11001000 : OUT <= 0;  //95 / 200 = 0
    16'b01011111_11001001 : OUT <= 0;  //95 / 201 = 0
    16'b01011111_11001010 : OUT <= 0;  //95 / 202 = 0
    16'b01011111_11001011 : OUT <= 0;  //95 / 203 = 0
    16'b01011111_11001100 : OUT <= 0;  //95 / 204 = 0
    16'b01011111_11001101 : OUT <= 0;  //95 / 205 = 0
    16'b01011111_11001110 : OUT <= 0;  //95 / 206 = 0
    16'b01011111_11001111 : OUT <= 0;  //95 / 207 = 0
    16'b01011111_11010000 : OUT <= 0;  //95 / 208 = 0
    16'b01011111_11010001 : OUT <= 0;  //95 / 209 = 0
    16'b01011111_11010010 : OUT <= 0;  //95 / 210 = 0
    16'b01011111_11010011 : OUT <= 0;  //95 / 211 = 0
    16'b01011111_11010100 : OUT <= 0;  //95 / 212 = 0
    16'b01011111_11010101 : OUT <= 0;  //95 / 213 = 0
    16'b01011111_11010110 : OUT <= 0;  //95 / 214 = 0
    16'b01011111_11010111 : OUT <= 0;  //95 / 215 = 0
    16'b01011111_11011000 : OUT <= 0;  //95 / 216 = 0
    16'b01011111_11011001 : OUT <= 0;  //95 / 217 = 0
    16'b01011111_11011010 : OUT <= 0;  //95 / 218 = 0
    16'b01011111_11011011 : OUT <= 0;  //95 / 219 = 0
    16'b01011111_11011100 : OUT <= 0;  //95 / 220 = 0
    16'b01011111_11011101 : OUT <= 0;  //95 / 221 = 0
    16'b01011111_11011110 : OUT <= 0;  //95 / 222 = 0
    16'b01011111_11011111 : OUT <= 0;  //95 / 223 = 0
    16'b01011111_11100000 : OUT <= 0;  //95 / 224 = 0
    16'b01011111_11100001 : OUT <= 0;  //95 / 225 = 0
    16'b01011111_11100010 : OUT <= 0;  //95 / 226 = 0
    16'b01011111_11100011 : OUT <= 0;  //95 / 227 = 0
    16'b01011111_11100100 : OUT <= 0;  //95 / 228 = 0
    16'b01011111_11100101 : OUT <= 0;  //95 / 229 = 0
    16'b01011111_11100110 : OUT <= 0;  //95 / 230 = 0
    16'b01011111_11100111 : OUT <= 0;  //95 / 231 = 0
    16'b01011111_11101000 : OUT <= 0;  //95 / 232 = 0
    16'b01011111_11101001 : OUT <= 0;  //95 / 233 = 0
    16'b01011111_11101010 : OUT <= 0;  //95 / 234 = 0
    16'b01011111_11101011 : OUT <= 0;  //95 / 235 = 0
    16'b01011111_11101100 : OUT <= 0;  //95 / 236 = 0
    16'b01011111_11101101 : OUT <= 0;  //95 / 237 = 0
    16'b01011111_11101110 : OUT <= 0;  //95 / 238 = 0
    16'b01011111_11101111 : OUT <= 0;  //95 / 239 = 0
    16'b01011111_11110000 : OUT <= 0;  //95 / 240 = 0
    16'b01011111_11110001 : OUT <= 0;  //95 / 241 = 0
    16'b01011111_11110010 : OUT <= 0;  //95 / 242 = 0
    16'b01011111_11110011 : OUT <= 0;  //95 / 243 = 0
    16'b01011111_11110100 : OUT <= 0;  //95 / 244 = 0
    16'b01011111_11110101 : OUT <= 0;  //95 / 245 = 0
    16'b01011111_11110110 : OUT <= 0;  //95 / 246 = 0
    16'b01011111_11110111 : OUT <= 0;  //95 / 247 = 0
    16'b01011111_11111000 : OUT <= 0;  //95 / 248 = 0
    16'b01011111_11111001 : OUT <= 0;  //95 / 249 = 0
    16'b01011111_11111010 : OUT <= 0;  //95 / 250 = 0
    16'b01011111_11111011 : OUT <= 0;  //95 / 251 = 0
    16'b01011111_11111100 : OUT <= 0;  //95 / 252 = 0
    16'b01011111_11111101 : OUT <= 0;  //95 / 253 = 0
    16'b01011111_11111110 : OUT <= 0;  //95 / 254 = 0
    16'b01011111_11111111 : OUT <= 0;  //95 / 255 = 0
    16'b01100000_00000000 : OUT <= 0;  //96 / 0 = 0
    16'b01100000_00000001 : OUT <= 96;  //96 / 1 = 96
    16'b01100000_00000010 : OUT <= 48;  //96 / 2 = 48
    16'b01100000_00000011 : OUT <= 32;  //96 / 3 = 32
    16'b01100000_00000100 : OUT <= 24;  //96 / 4 = 24
    16'b01100000_00000101 : OUT <= 19;  //96 / 5 = 19
    16'b01100000_00000110 : OUT <= 16;  //96 / 6 = 16
    16'b01100000_00000111 : OUT <= 13;  //96 / 7 = 13
    16'b01100000_00001000 : OUT <= 12;  //96 / 8 = 12
    16'b01100000_00001001 : OUT <= 10;  //96 / 9 = 10
    16'b01100000_00001010 : OUT <= 9;  //96 / 10 = 9
    16'b01100000_00001011 : OUT <= 8;  //96 / 11 = 8
    16'b01100000_00001100 : OUT <= 8;  //96 / 12 = 8
    16'b01100000_00001101 : OUT <= 7;  //96 / 13 = 7
    16'b01100000_00001110 : OUT <= 6;  //96 / 14 = 6
    16'b01100000_00001111 : OUT <= 6;  //96 / 15 = 6
    16'b01100000_00010000 : OUT <= 6;  //96 / 16 = 6
    16'b01100000_00010001 : OUT <= 5;  //96 / 17 = 5
    16'b01100000_00010010 : OUT <= 5;  //96 / 18 = 5
    16'b01100000_00010011 : OUT <= 5;  //96 / 19 = 5
    16'b01100000_00010100 : OUT <= 4;  //96 / 20 = 4
    16'b01100000_00010101 : OUT <= 4;  //96 / 21 = 4
    16'b01100000_00010110 : OUT <= 4;  //96 / 22 = 4
    16'b01100000_00010111 : OUT <= 4;  //96 / 23 = 4
    16'b01100000_00011000 : OUT <= 4;  //96 / 24 = 4
    16'b01100000_00011001 : OUT <= 3;  //96 / 25 = 3
    16'b01100000_00011010 : OUT <= 3;  //96 / 26 = 3
    16'b01100000_00011011 : OUT <= 3;  //96 / 27 = 3
    16'b01100000_00011100 : OUT <= 3;  //96 / 28 = 3
    16'b01100000_00011101 : OUT <= 3;  //96 / 29 = 3
    16'b01100000_00011110 : OUT <= 3;  //96 / 30 = 3
    16'b01100000_00011111 : OUT <= 3;  //96 / 31 = 3
    16'b01100000_00100000 : OUT <= 3;  //96 / 32 = 3
    16'b01100000_00100001 : OUT <= 2;  //96 / 33 = 2
    16'b01100000_00100010 : OUT <= 2;  //96 / 34 = 2
    16'b01100000_00100011 : OUT <= 2;  //96 / 35 = 2
    16'b01100000_00100100 : OUT <= 2;  //96 / 36 = 2
    16'b01100000_00100101 : OUT <= 2;  //96 / 37 = 2
    16'b01100000_00100110 : OUT <= 2;  //96 / 38 = 2
    16'b01100000_00100111 : OUT <= 2;  //96 / 39 = 2
    16'b01100000_00101000 : OUT <= 2;  //96 / 40 = 2
    16'b01100000_00101001 : OUT <= 2;  //96 / 41 = 2
    16'b01100000_00101010 : OUT <= 2;  //96 / 42 = 2
    16'b01100000_00101011 : OUT <= 2;  //96 / 43 = 2
    16'b01100000_00101100 : OUT <= 2;  //96 / 44 = 2
    16'b01100000_00101101 : OUT <= 2;  //96 / 45 = 2
    16'b01100000_00101110 : OUT <= 2;  //96 / 46 = 2
    16'b01100000_00101111 : OUT <= 2;  //96 / 47 = 2
    16'b01100000_00110000 : OUT <= 2;  //96 / 48 = 2
    16'b01100000_00110001 : OUT <= 1;  //96 / 49 = 1
    16'b01100000_00110010 : OUT <= 1;  //96 / 50 = 1
    16'b01100000_00110011 : OUT <= 1;  //96 / 51 = 1
    16'b01100000_00110100 : OUT <= 1;  //96 / 52 = 1
    16'b01100000_00110101 : OUT <= 1;  //96 / 53 = 1
    16'b01100000_00110110 : OUT <= 1;  //96 / 54 = 1
    16'b01100000_00110111 : OUT <= 1;  //96 / 55 = 1
    16'b01100000_00111000 : OUT <= 1;  //96 / 56 = 1
    16'b01100000_00111001 : OUT <= 1;  //96 / 57 = 1
    16'b01100000_00111010 : OUT <= 1;  //96 / 58 = 1
    16'b01100000_00111011 : OUT <= 1;  //96 / 59 = 1
    16'b01100000_00111100 : OUT <= 1;  //96 / 60 = 1
    16'b01100000_00111101 : OUT <= 1;  //96 / 61 = 1
    16'b01100000_00111110 : OUT <= 1;  //96 / 62 = 1
    16'b01100000_00111111 : OUT <= 1;  //96 / 63 = 1
    16'b01100000_01000000 : OUT <= 1;  //96 / 64 = 1
    16'b01100000_01000001 : OUT <= 1;  //96 / 65 = 1
    16'b01100000_01000010 : OUT <= 1;  //96 / 66 = 1
    16'b01100000_01000011 : OUT <= 1;  //96 / 67 = 1
    16'b01100000_01000100 : OUT <= 1;  //96 / 68 = 1
    16'b01100000_01000101 : OUT <= 1;  //96 / 69 = 1
    16'b01100000_01000110 : OUT <= 1;  //96 / 70 = 1
    16'b01100000_01000111 : OUT <= 1;  //96 / 71 = 1
    16'b01100000_01001000 : OUT <= 1;  //96 / 72 = 1
    16'b01100000_01001001 : OUT <= 1;  //96 / 73 = 1
    16'b01100000_01001010 : OUT <= 1;  //96 / 74 = 1
    16'b01100000_01001011 : OUT <= 1;  //96 / 75 = 1
    16'b01100000_01001100 : OUT <= 1;  //96 / 76 = 1
    16'b01100000_01001101 : OUT <= 1;  //96 / 77 = 1
    16'b01100000_01001110 : OUT <= 1;  //96 / 78 = 1
    16'b01100000_01001111 : OUT <= 1;  //96 / 79 = 1
    16'b01100000_01010000 : OUT <= 1;  //96 / 80 = 1
    16'b01100000_01010001 : OUT <= 1;  //96 / 81 = 1
    16'b01100000_01010010 : OUT <= 1;  //96 / 82 = 1
    16'b01100000_01010011 : OUT <= 1;  //96 / 83 = 1
    16'b01100000_01010100 : OUT <= 1;  //96 / 84 = 1
    16'b01100000_01010101 : OUT <= 1;  //96 / 85 = 1
    16'b01100000_01010110 : OUT <= 1;  //96 / 86 = 1
    16'b01100000_01010111 : OUT <= 1;  //96 / 87 = 1
    16'b01100000_01011000 : OUT <= 1;  //96 / 88 = 1
    16'b01100000_01011001 : OUT <= 1;  //96 / 89 = 1
    16'b01100000_01011010 : OUT <= 1;  //96 / 90 = 1
    16'b01100000_01011011 : OUT <= 1;  //96 / 91 = 1
    16'b01100000_01011100 : OUT <= 1;  //96 / 92 = 1
    16'b01100000_01011101 : OUT <= 1;  //96 / 93 = 1
    16'b01100000_01011110 : OUT <= 1;  //96 / 94 = 1
    16'b01100000_01011111 : OUT <= 1;  //96 / 95 = 1
    16'b01100000_01100000 : OUT <= 1;  //96 / 96 = 1
    16'b01100000_01100001 : OUT <= 0;  //96 / 97 = 0
    16'b01100000_01100010 : OUT <= 0;  //96 / 98 = 0
    16'b01100000_01100011 : OUT <= 0;  //96 / 99 = 0
    16'b01100000_01100100 : OUT <= 0;  //96 / 100 = 0
    16'b01100000_01100101 : OUT <= 0;  //96 / 101 = 0
    16'b01100000_01100110 : OUT <= 0;  //96 / 102 = 0
    16'b01100000_01100111 : OUT <= 0;  //96 / 103 = 0
    16'b01100000_01101000 : OUT <= 0;  //96 / 104 = 0
    16'b01100000_01101001 : OUT <= 0;  //96 / 105 = 0
    16'b01100000_01101010 : OUT <= 0;  //96 / 106 = 0
    16'b01100000_01101011 : OUT <= 0;  //96 / 107 = 0
    16'b01100000_01101100 : OUT <= 0;  //96 / 108 = 0
    16'b01100000_01101101 : OUT <= 0;  //96 / 109 = 0
    16'b01100000_01101110 : OUT <= 0;  //96 / 110 = 0
    16'b01100000_01101111 : OUT <= 0;  //96 / 111 = 0
    16'b01100000_01110000 : OUT <= 0;  //96 / 112 = 0
    16'b01100000_01110001 : OUT <= 0;  //96 / 113 = 0
    16'b01100000_01110010 : OUT <= 0;  //96 / 114 = 0
    16'b01100000_01110011 : OUT <= 0;  //96 / 115 = 0
    16'b01100000_01110100 : OUT <= 0;  //96 / 116 = 0
    16'b01100000_01110101 : OUT <= 0;  //96 / 117 = 0
    16'b01100000_01110110 : OUT <= 0;  //96 / 118 = 0
    16'b01100000_01110111 : OUT <= 0;  //96 / 119 = 0
    16'b01100000_01111000 : OUT <= 0;  //96 / 120 = 0
    16'b01100000_01111001 : OUT <= 0;  //96 / 121 = 0
    16'b01100000_01111010 : OUT <= 0;  //96 / 122 = 0
    16'b01100000_01111011 : OUT <= 0;  //96 / 123 = 0
    16'b01100000_01111100 : OUT <= 0;  //96 / 124 = 0
    16'b01100000_01111101 : OUT <= 0;  //96 / 125 = 0
    16'b01100000_01111110 : OUT <= 0;  //96 / 126 = 0
    16'b01100000_01111111 : OUT <= 0;  //96 / 127 = 0
    16'b01100000_10000000 : OUT <= 0;  //96 / 128 = 0
    16'b01100000_10000001 : OUT <= 0;  //96 / 129 = 0
    16'b01100000_10000010 : OUT <= 0;  //96 / 130 = 0
    16'b01100000_10000011 : OUT <= 0;  //96 / 131 = 0
    16'b01100000_10000100 : OUT <= 0;  //96 / 132 = 0
    16'b01100000_10000101 : OUT <= 0;  //96 / 133 = 0
    16'b01100000_10000110 : OUT <= 0;  //96 / 134 = 0
    16'b01100000_10000111 : OUT <= 0;  //96 / 135 = 0
    16'b01100000_10001000 : OUT <= 0;  //96 / 136 = 0
    16'b01100000_10001001 : OUT <= 0;  //96 / 137 = 0
    16'b01100000_10001010 : OUT <= 0;  //96 / 138 = 0
    16'b01100000_10001011 : OUT <= 0;  //96 / 139 = 0
    16'b01100000_10001100 : OUT <= 0;  //96 / 140 = 0
    16'b01100000_10001101 : OUT <= 0;  //96 / 141 = 0
    16'b01100000_10001110 : OUT <= 0;  //96 / 142 = 0
    16'b01100000_10001111 : OUT <= 0;  //96 / 143 = 0
    16'b01100000_10010000 : OUT <= 0;  //96 / 144 = 0
    16'b01100000_10010001 : OUT <= 0;  //96 / 145 = 0
    16'b01100000_10010010 : OUT <= 0;  //96 / 146 = 0
    16'b01100000_10010011 : OUT <= 0;  //96 / 147 = 0
    16'b01100000_10010100 : OUT <= 0;  //96 / 148 = 0
    16'b01100000_10010101 : OUT <= 0;  //96 / 149 = 0
    16'b01100000_10010110 : OUT <= 0;  //96 / 150 = 0
    16'b01100000_10010111 : OUT <= 0;  //96 / 151 = 0
    16'b01100000_10011000 : OUT <= 0;  //96 / 152 = 0
    16'b01100000_10011001 : OUT <= 0;  //96 / 153 = 0
    16'b01100000_10011010 : OUT <= 0;  //96 / 154 = 0
    16'b01100000_10011011 : OUT <= 0;  //96 / 155 = 0
    16'b01100000_10011100 : OUT <= 0;  //96 / 156 = 0
    16'b01100000_10011101 : OUT <= 0;  //96 / 157 = 0
    16'b01100000_10011110 : OUT <= 0;  //96 / 158 = 0
    16'b01100000_10011111 : OUT <= 0;  //96 / 159 = 0
    16'b01100000_10100000 : OUT <= 0;  //96 / 160 = 0
    16'b01100000_10100001 : OUT <= 0;  //96 / 161 = 0
    16'b01100000_10100010 : OUT <= 0;  //96 / 162 = 0
    16'b01100000_10100011 : OUT <= 0;  //96 / 163 = 0
    16'b01100000_10100100 : OUT <= 0;  //96 / 164 = 0
    16'b01100000_10100101 : OUT <= 0;  //96 / 165 = 0
    16'b01100000_10100110 : OUT <= 0;  //96 / 166 = 0
    16'b01100000_10100111 : OUT <= 0;  //96 / 167 = 0
    16'b01100000_10101000 : OUT <= 0;  //96 / 168 = 0
    16'b01100000_10101001 : OUT <= 0;  //96 / 169 = 0
    16'b01100000_10101010 : OUT <= 0;  //96 / 170 = 0
    16'b01100000_10101011 : OUT <= 0;  //96 / 171 = 0
    16'b01100000_10101100 : OUT <= 0;  //96 / 172 = 0
    16'b01100000_10101101 : OUT <= 0;  //96 / 173 = 0
    16'b01100000_10101110 : OUT <= 0;  //96 / 174 = 0
    16'b01100000_10101111 : OUT <= 0;  //96 / 175 = 0
    16'b01100000_10110000 : OUT <= 0;  //96 / 176 = 0
    16'b01100000_10110001 : OUT <= 0;  //96 / 177 = 0
    16'b01100000_10110010 : OUT <= 0;  //96 / 178 = 0
    16'b01100000_10110011 : OUT <= 0;  //96 / 179 = 0
    16'b01100000_10110100 : OUT <= 0;  //96 / 180 = 0
    16'b01100000_10110101 : OUT <= 0;  //96 / 181 = 0
    16'b01100000_10110110 : OUT <= 0;  //96 / 182 = 0
    16'b01100000_10110111 : OUT <= 0;  //96 / 183 = 0
    16'b01100000_10111000 : OUT <= 0;  //96 / 184 = 0
    16'b01100000_10111001 : OUT <= 0;  //96 / 185 = 0
    16'b01100000_10111010 : OUT <= 0;  //96 / 186 = 0
    16'b01100000_10111011 : OUT <= 0;  //96 / 187 = 0
    16'b01100000_10111100 : OUT <= 0;  //96 / 188 = 0
    16'b01100000_10111101 : OUT <= 0;  //96 / 189 = 0
    16'b01100000_10111110 : OUT <= 0;  //96 / 190 = 0
    16'b01100000_10111111 : OUT <= 0;  //96 / 191 = 0
    16'b01100000_11000000 : OUT <= 0;  //96 / 192 = 0
    16'b01100000_11000001 : OUT <= 0;  //96 / 193 = 0
    16'b01100000_11000010 : OUT <= 0;  //96 / 194 = 0
    16'b01100000_11000011 : OUT <= 0;  //96 / 195 = 0
    16'b01100000_11000100 : OUT <= 0;  //96 / 196 = 0
    16'b01100000_11000101 : OUT <= 0;  //96 / 197 = 0
    16'b01100000_11000110 : OUT <= 0;  //96 / 198 = 0
    16'b01100000_11000111 : OUT <= 0;  //96 / 199 = 0
    16'b01100000_11001000 : OUT <= 0;  //96 / 200 = 0
    16'b01100000_11001001 : OUT <= 0;  //96 / 201 = 0
    16'b01100000_11001010 : OUT <= 0;  //96 / 202 = 0
    16'b01100000_11001011 : OUT <= 0;  //96 / 203 = 0
    16'b01100000_11001100 : OUT <= 0;  //96 / 204 = 0
    16'b01100000_11001101 : OUT <= 0;  //96 / 205 = 0
    16'b01100000_11001110 : OUT <= 0;  //96 / 206 = 0
    16'b01100000_11001111 : OUT <= 0;  //96 / 207 = 0
    16'b01100000_11010000 : OUT <= 0;  //96 / 208 = 0
    16'b01100000_11010001 : OUT <= 0;  //96 / 209 = 0
    16'b01100000_11010010 : OUT <= 0;  //96 / 210 = 0
    16'b01100000_11010011 : OUT <= 0;  //96 / 211 = 0
    16'b01100000_11010100 : OUT <= 0;  //96 / 212 = 0
    16'b01100000_11010101 : OUT <= 0;  //96 / 213 = 0
    16'b01100000_11010110 : OUT <= 0;  //96 / 214 = 0
    16'b01100000_11010111 : OUT <= 0;  //96 / 215 = 0
    16'b01100000_11011000 : OUT <= 0;  //96 / 216 = 0
    16'b01100000_11011001 : OUT <= 0;  //96 / 217 = 0
    16'b01100000_11011010 : OUT <= 0;  //96 / 218 = 0
    16'b01100000_11011011 : OUT <= 0;  //96 / 219 = 0
    16'b01100000_11011100 : OUT <= 0;  //96 / 220 = 0
    16'b01100000_11011101 : OUT <= 0;  //96 / 221 = 0
    16'b01100000_11011110 : OUT <= 0;  //96 / 222 = 0
    16'b01100000_11011111 : OUT <= 0;  //96 / 223 = 0
    16'b01100000_11100000 : OUT <= 0;  //96 / 224 = 0
    16'b01100000_11100001 : OUT <= 0;  //96 / 225 = 0
    16'b01100000_11100010 : OUT <= 0;  //96 / 226 = 0
    16'b01100000_11100011 : OUT <= 0;  //96 / 227 = 0
    16'b01100000_11100100 : OUT <= 0;  //96 / 228 = 0
    16'b01100000_11100101 : OUT <= 0;  //96 / 229 = 0
    16'b01100000_11100110 : OUT <= 0;  //96 / 230 = 0
    16'b01100000_11100111 : OUT <= 0;  //96 / 231 = 0
    16'b01100000_11101000 : OUT <= 0;  //96 / 232 = 0
    16'b01100000_11101001 : OUT <= 0;  //96 / 233 = 0
    16'b01100000_11101010 : OUT <= 0;  //96 / 234 = 0
    16'b01100000_11101011 : OUT <= 0;  //96 / 235 = 0
    16'b01100000_11101100 : OUT <= 0;  //96 / 236 = 0
    16'b01100000_11101101 : OUT <= 0;  //96 / 237 = 0
    16'b01100000_11101110 : OUT <= 0;  //96 / 238 = 0
    16'b01100000_11101111 : OUT <= 0;  //96 / 239 = 0
    16'b01100000_11110000 : OUT <= 0;  //96 / 240 = 0
    16'b01100000_11110001 : OUT <= 0;  //96 / 241 = 0
    16'b01100000_11110010 : OUT <= 0;  //96 / 242 = 0
    16'b01100000_11110011 : OUT <= 0;  //96 / 243 = 0
    16'b01100000_11110100 : OUT <= 0;  //96 / 244 = 0
    16'b01100000_11110101 : OUT <= 0;  //96 / 245 = 0
    16'b01100000_11110110 : OUT <= 0;  //96 / 246 = 0
    16'b01100000_11110111 : OUT <= 0;  //96 / 247 = 0
    16'b01100000_11111000 : OUT <= 0;  //96 / 248 = 0
    16'b01100000_11111001 : OUT <= 0;  //96 / 249 = 0
    16'b01100000_11111010 : OUT <= 0;  //96 / 250 = 0
    16'b01100000_11111011 : OUT <= 0;  //96 / 251 = 0
    16'b01100000_11111100 : OUT <= 0;  //96 / 252 = 0
    16'b01100000_11111101 : OUT <= 0;  //96 / 253 = 0
    16'b01100000_11111110 : OUT <= 0;  //96 / 254 = 0
    16'b01100000_11111111 : OUT <= 0;  //96 / 255 = 0
    16'b01100001_00000000 : OUT <= 0;  //97 / 0 = 0
    16'b01100001_00000001 : OUT <= 97;  //97 / 1 = 97
    16'b01100001_00000010 : OUT <= 48;  //97 / 2 = 48
    16'b01100001_00000011 : OUT <= 32;  //97 / 3 = 32
    16'b01100001_00000100 : OUT <= 24;  //97 / 4 = 24
    16'b01100001_00000101 : OUT <= 19;  //97 / 5 = 19
    16'b01100001_00000110 : OUT <= 16;  //97 / 6 = 16
    16'b01100001_00000111 : OUT <= 13;  //97 / 7 = 13
    16'b01100001_00001000 : OUT <= 12;  //97 / 8 = 12
    16'b01100001_00001001 : OUT <= 10;  //97 / 9 = 10
    16'b01100001_00001010 : OUT <= 9;  //97 / 10 = 9
    16'b01100001_00001011 : OUT <= 8;  //97 / 11 = 8
    16'b01100001_00001100 : OUT <= 8;  //97 / 12 = 8
    16'b01100001_00001101 : OUT <= 7;  //97 / 13 = 7
    16'b01100001_00001110 : OUT <= 6;  //97 / 14 = 6
    16'b01100001_00001111 : OUT <= 6;  //97 / 15 = 6
    16'b01100001_00010000 : OUT <= 6;  //97 / 16 = 6
    16'b01100001_00010001 : OUT <= 5;  //97 / 17 = 5
    16'b01100001_00010010 : OUT <= 5;  //97 / 18 = 5
    16'b01100001_00010011 : OUT <= 5;  //97 / 19 = 5
    16'b01100001_00010100 : OUT <= 4;  //97 / 20 = 4
    16'b01100001_00010101 : OUT <= 4;  //97 / 21 = 4
    16'b01100001_00010110 : OUT <= 4;  //97 / 22 = 4
    16'b01100001_00010111 : OUT <= 4;  //97 / 23 = 4
    16'b01100001_00011000 : OUT <= 4;  //97 / 24 = 4
    16'b01100001_00011001 : OUT <= 3;  //97 / 25 = 3
    16'b01100001_00011010 : OUT <= 3;  //97 / 26 = 3
    16'b01100001_00011011 : OUT <= 3;  //97 / 27 = 3
    16'b01100001_00011100 : OUT <= 3;  //97 / 28 = 3
    16'b01100001_00011101 : OUT <= 3;  //97 / 29 = 3
    16'b01100001_00011110 : OUT <= 3;  //97 / 30 = 3
    16'b01100001_00011111 : OUT <= 3;  //97 / 31 = 3
    16'b01100001_00100000 : OUT <= 3;  //97 / 32 = 3
    16'b01100001_00100001 : OUT <= 2;  //97 / 33 = 2
    16'b01100001_00100010 : OUT <= 2;  //97 / 34 = 2
    16'b01100001_00100011 : OUT <= 2;  //97 / 35 = 2
    16'b01100001_00100100 : OUT <= 2;  //97 / 36 = 2
    16'b01100001_00100101 : OUT <= 2;  //97 / 37 = 2
    16'b01100001_00100110 : OUT <= 2;  //97 / 38 = 2
    16'b01100001_00100111 : OUT <= 2;  //97 / 39 = 2
    16'b01100001_00101000 : OUT <= 2;  //97 / 40 = 2
    16'b01100001_00101001 : OUT <= 2;  //97 / 41 = 2
    16'b01100001_00101010 : OUT <= 2;  //97 / 42 = 2
    16'b01100001_00101011 : OUT <= 2;  //97 / 43 = 2
    16'b01100001_00101100 : OUT <= 2;  //97 / 44 = 2
    16'b01100001_00101101 : OUT <= 2;  //97 / 45 = 2
    16'b01100001_00101110 : OUT <= 2;  //97 / 46 = 2
    16'b01100001_00101111 : OUT <= 2;  //97 / 47 = 2
    16'b01100001_00110000 : OUT <= 2;  //97 / 48 = 2
    16'b01100001_00110001 : OUT <= 1;  //97 / 49 = 1
    16'b01100001_00110010 : OUT <= 1;  //97 / 50 = 1
    16'b01100001_00110011 : OUT <= 1;  //97 / 51 = 1
    16'b01100001_00110100 : OUT <= 1;  //97 / 52 = 1
    16'b01100001_00110101 : OUT <= 1;  //97 / 53 = 1
    16'b01100001_00110110 : OUT <= 1;  //97 / 54 = 1
    16'b01100001_00110111 : OUT <= 1;  //97 / 55 = 1
    16'b01100001_00111000 : OUT <= 1;  //97 / 56 = 1
    16'b01100001_00111001 : OUT <= 1;  //97 / 57 = 1
    16'b01100001_00111010 : OUT <= 1;  //97 / 58 = 1
    16'b01100001_00111011 : OUT <= 1;  //97 / 59 = 1
    16'b01100001_00111100 : OUT <= 1;  //97 / 60 = 1
    16'b01100001_00111101 : OUT <= 1;  //97 / 61 = 1
    16'b01100001_00111110 : OUT <= 1;  //97 / 62 = 1
    16'b01100001_00111111 : OUT <= 1;  //97 / 63 = 1
    16'b01100001_01000000 : OUT <= 1;  //97 / 64 = 1
    16'b01100001_01000001 : OUT <= 1;  //97 / 65 = 1
    16'b01100001_01000010 : OUT <= 1;  //97 / 66 = 1
    16'b01100001_01000011 : OUT <= 1;  //97 / 67 = 1
    16'b01100001_01000100 : OUT <= 1;  //97 / 68 = 1
    16'b01100001_01000101 : OUT <= 1;  //97 / 69 = 1
    16'b01100001_01000110 : OUT <= 1;  //97 / 70 = 1
    16'b01100001_01000111 : OUT <= 1;  //97 / 71 = 1
    16'b01100001_01001000 : OUT <= 1;  //97 / 72 = 1
    16'b01100001_01001001 : OUT <= 1;  //97 / 73 = 1
    16'b01100001_01001010 : OUT <= 1;  //97 / 74 = 1
    16'b01100001_01001011 : OUT <= 1;  //97 / 75 = 1
    16'b01100001_01001100 : OUT <= 1;  //97 / 76 = 1
    16'b01100001_01001101 : OUT <= 1;  //97 / 77 = 1
    16'b01100001_01001110 : OUT <= 1;  //97 / 78 = 1
    16'b01100001_01001111 : OUT <= 1;  //97 / 79 = 1
    16'b01100001_01010000 : OUT <= 1;  //97 / 80 = 1
    16'b01100001_01010001 : OUT <= 1;  //97 / 81 = 1
    16'b01100001_01010010 : OUT <= 1;  //97 / 82 = 1
    16'b01100001_01010011 : OUT <= 1;  //97 / 83 = 1
    16'b01100001_01010100 : OUT <= 1;  //97 / 84 = 1
    16'b01100001_01010101 : OUT <= 1;  //97 / 85 = 1
    16'b01100001_01010110 : OUT <= 1;  //97 / 86 = 1
    16'b01100001_01010111 : OUT <= 1;  //97 / 87 = 1
    16'b01100001_01011000 : OUT <= 1;  //97 / 88 = 1
    16'b01100001_01011001 : OUT <= 1;  //97 / 89 = 1
    16'b01100001_01011010 : OUT <= 1;  //97 / 90 = 1
    16'b01100001_01011011 : OUT <= 1;  //97 / 91 = 1
    16'b01100001_01011100 : OUT <= 1;  //97 / 92 = 1
    16'b01100001_01011101 : OUT <= 1;  //97 / 93 = 1
    16'b01100001_01011110 : OUT <= 1;  //97 / 94 = 1
    16'b01100001_01011111 : OUT <= 1;  //97 / 95 = 1
    16'b01100001_01100000 : OUT <= 1;  //97 / 96 = 1
    16'b01100001_01100001 : OUT <= 1;  //97 / 97 = 1
    16'b01100001_01100010 : OUT <= 0;  //97 / 98 = 0
    16'b01100001_01100011 : OUT <= 0;  //97 / 99 = 0
    16'b01100001_01100100 : OUT <= 0;  //97 / 100 = 0
    16'b01100001_01100101 : OUT <= 0;  //97 / 101 = 0
    16'b01100001_01100110 : OUT <= 0;  //97 / 102 = 0
    16'b01100001_01100111 : OUT <= 0;  //97 / 103 = 0
    16'b01100001_01101000 : OUT <= 0;  //97 / 104 = 0
    16'b01100001_01101001 : OUT <= 0;  //97 / 105 = 0
    16'b01100001_01101010 : OUT <= 0;  //97 / 106 = 0
    16'b01100001_01101011 : OUT <= 0;  //97 / 107 = 0
    16'b01100001_01101100 : OUT <= 0;  //97 / 108 = 0
    16'b01100001_01101101 : OUT <= 0;  //97 / 109 = 0
    16'b01100001_01101110 : OUT <= 0;  //97 / 110 = 0
    16'b01100001_01101111 : OUT <= 0;  //97 / 111 = 0
    16'b01100001_01110000 : OUT <= 0;  //97 / 112 = 0
    16'b01100001_01110001 : OUT <= 0;  //97 / 113 = 0
    16'b01100001_01110010 : OUT <= 0;  //97 / 114 = 0
    16'b01100001_01110011 : OUT <= 0;  //97 / 115 = 0
    16'b01100001_01110100 : OUT <= 0;  //97 / 116 = 0
    16'b01100001_01110101 : OUT <= 0;  //97 / 117 = 0
    16'b01100001_01110110 : OUT <= 0;  //97 / 118 = 0
    16'b01100001_01110111 : OUT <= 0;  //97 / 119 = 0
    16'b01100001_01111000 : OUT <= 0;  //97 / 120 = 0
    16'b01100001_01111001 : OUT <= 0;  //97 / 121 = 0
    16'b01100001_01111010 : OUT <= 0;  //97 / 122 = 0
    16'b01100001_01111011 : OUT <= 0;  //97 / 123 = 0
    16'b01100001_01111100 : OUT <= 0;  //97 / 124 = 0
    16'b01100001_01111101 : OUT <= 0;  //97 / 125 = 0
    16'b01100001_01111110 : OUT <= 0;  //97 / 126 = 0
    16'b01100001_01111111 : OUT <= 0;  //97 / 127 = 0
    16'b01100001_10000000 : OUT <= 0;  //97 / 128 = 0
    16'b01100001_10000001 : OUT <= 0;  //97 / 129 = 0
    16'b01100001_10000010 : OUT <= 0;  //97 / 130 = 0
    16'b01100001_10000011 : OUT <= 0;  //97 / 131 = 0
    16'b01100001_10000100 : OUT <= 0;  //97 / 132 = 0
    16'b01100001_10000101 : OUT <= 0;  //97 / 133 = 0
    16'b01100001_10000110 : OUT <= 0;  //97 / 134 = 0
    16'b01100001_10000111 : OUT <= 0;  //97 / 135 = 0
    16'b01100001_10001000 : OUT <= 0;  //97 / 136 = 0
    16'b01100001_10001001 : OUT <= 0;  //97 / 137 = 0
    16'b01100001_10001010 : OUT <= 0;  //97 / 138 = 0
    16'b01100001_10001011 : OUT <= 0;  //97 / 139 = 0
    16'b01100001_10001100 : OUT <= 0;  //97 / 140 = 0
    16'b01100001_10001101 : OUT <= 0;  //97 / 141 = 0
    16'b01100001_10001110 : OUT <= 0;  //97 / 142 = 0
    16'b01100001_10001111 : OUT <= 0;  //97 / 143 = 0
    16'b01100001_10010000 : OUT <= 0;  //97 / 144 = 0
    16'b01100001_10010001 : OUT <= 0;  //97 / 145 = 0
    16'b01100001_10010010 : OUT <= 0;  //97 / 146 = 0
    16'b01100001_10010011 : OUT <= 0;  //97 / 147 = 0
    16'b01100001_10010100 : OUT <= 0;  //97 / 148 = 0
    16'b01100001_10010101 : OUT <= 0;  //97 / 149 = 0
    16'b01100001_10010110 : OUT <= 0;  //97 / 150 = 0
    16'b01100001_10010111 : OUT <= 0;  //97 / 151 = 0
    16'b01100001_10011000 : OUT <= 0;  //97 / 152 = 0
    16'b01100001_10011001 : OUT <= 0;  //97 / 153 = 0
    16'b01100001_10011010 : OUT <= 0;  //97 / 154 = 0
    16'b01100001_10011011 : OUT <= 0;  //97 / 155 = 0
    16'b01100001_10011100 : OUT <= 0;  //97 / 156 = 0
    16'b01100001_10011101 : OUT <= 0;  //97 / 157 = 0
    16'b01100001_10011110 : OUT <= 0;  //97 / 158 = 0
    16'b01100001_10011111 : OUT <= 0;  //97 / 159 = 0
    16'b01100001_10100000 : OUT <= 0;  //97 / 160 = 0
    16'b01100001_10100001 : OUT <= 0;  //97 / 161 = 0
    16'b01100001_10100010 : OUT <= 0;  //97 / 162 = 0
    16'b01100001_10100011 : OUT <= 0;  //97 / 163 = 0
    16'b01100001_10100100 : OUT <= 0;  //97 / 164 = 0
    16'b01100001_10100101 : OUT <= 0;  //97 / 165 = 0
    16'b01100001_10100110 : OUT <= 0;  //97 / 166 = 0
    16'b01100001_10100111 : OUT <= 0;  //97 / 167 = 0
    16'b01100001_10101000 : OUT <= 0;  //97 / 168 = 0
    16'b01100001_10101001 : OUT <= 0;  //97 / 169 = 0
    16'b01100001_10101010 : OUT <= 0;  //97 / 170 = 0
    16'b01100001_10101011 : OUT <= 0;  //97 / 171 = 0
    16'b01100001_10101100 : OUT <= 0;  //97 / 172 = 0
    16'b01100001_10101101 : OUT <= 0;  //97 / 173 = 0
    16'b01100001_10101110 : OUT <= 0;  //97 / 174 = 0
    16'b01100001_10101111 : OUT <= 0;  //97 / 175 = 0
    16'b01100001_10110000 : OUT <= 0;  //97 / 176 = 0
    16'b01100001_10110001 : OUT <= 0;  //97 / 177 = 0
    16'b01100001_10110010 : OUT <= 0;  //97 / 178 = 0
    16'b01100001_10110011 : OUT <= 0;  //97 / 179 = 0
    16'b01100001_10110100 : OUT <= 0;  //97 / 180 = 0
    16'b01100001_10110101 : OUT <= 0;  //97 / 181 = 0
    16'b01100001_10110110 : OUT <= 0;  //97 / 182 = 0
    16'b01100001_10110111 : OUT <= 0;  //97 / 183 = 0
    16'b01100001_10111000 : OUT <= 0;  //97 / 184 = 0
    16'b01100001_10111001 : OUT <= 0;  //97 / 185 = 0
    16'b01100001_10111010 : OUT <= 0;  //97 / 186 = 0
    16'b01100001_10111011 : OUT <= 0;  //97 / 187 = 0
    16'b01100001_10111100 : OUT <= 0;  //97 / 188 = 0
    16'b01100001_10111101 : OUT <= 0;  //97 / 189 = 0
    16'b01100001_10111110 : OUT <= 0;  //97 / 190 = 0
    16'b01100001_10111111 : OUT <= 0;  //97 / 191 = 0
    16'b01100001_11000000 : OUT <= 0;  //97 / 192 = 0
    16'b01100001_11000001 : OUT <= 0;  //97 / 193 = 0
    16'b01100001_11000010 : OUT <= 0;  //97 / 194 = 0
    16'b01100001_11000011 : OUT <= 0;  //97 / 195 = 0
    16'b01100001_11000100 : OUT <= 0;  //97 / 196 = 0
    16'b01100001_11000101 : OUT <= 0;  //97 / 197 = 0
    16'b01100001_11000110 : OUT <= 0;  //97 / 198 = 0
    16'b01100001_11000111 : OUT <= 0;  //97 / 199 = 0
    16'b01100001_11001000 : OUT <= 0;  //97 / 200 = 0
    16'b01100001_11001001 : OUT <= 0;  //97 / 201 = 0
    16'b01100001_11001010 : OUT <= 0;  //97 / 202 = 0
    16'b01100001_11001011 : OUT <= 0;  //97 / 203 = 0
    16'b01100001_11001100 : OUT <= 0;  //97 / 204 = 0
    16'b01100001_11001101 : OUT <= 0;  //97 / 205 = 0
    16'b01100001_11001110 : OUT <= 0;  //97 / 206 = 0
    16'b01100001_11001111 : OUT <= 0;  //97 / 207 = 0
    16'b01100001_11010000 : OUT <= 0;  //97 / 208 = 0
    16'b01100001_11010001 : OUT <= 0;  //97 / 209 = 0
    16'b01100001_11010010 : OUT <= 0;  //97 / 210 = 0
    16'b01100001_11010011 : OUT <= 0;  //97 / 211 = 0
    16'b01100001_11010100 : OUT <= 0;  //97 / 212 = 0
    16'b01100001_11010101 : OUT <= 0;  //97 / 213 = 0
    16'b01100001_11010110 : OUT <= 0;  //97 / 214 = 0
    16'b01100001_11010111 : OUT <= 0;  //97 / 215 = 0
    16'b01100001_11011000 : OUT <= 0;  //97 / 216 = 0
    16'b01100001_11011001 : OUT <= 0;  //97 / 217 = 0
    16'b01100001_11011010 : OUT <= 0;  //97 / 218 = 0
    16'b01100001_11011011 : OUT <= 0;  //97 / 219 = 0
    16'b01100001_11011100 : OUT <= 0;  //97 / 220 = 0
    16'b01100001_11011101 : OUT <= 0;  //97 / 221 = 0
    16'b01100001_11011110 : OUT <= 0;  //97 / 222 = 0
    16'b01100001_11011111 : OUT <= 0;  //97 / 223 = 0
    16'b01100001_11100000 : OUT <= 0;  //97 / 224 = 0
    16'b01100001_11100001 : OUT <= 0;  //97 / 225 = 0
    16'b01100001_11100010 : OUT <= 0;  //97 / 226 = 0
    16'b01100001_11100011 : OUT <= 0;  //97 / 227 = 0
    16'b01100001_11100100 : OUT <= 0;  //97 / 228 = 0
    16'b01100001_11100101 : OUT <= 0;  //97 / 229 = 0
    16'b01100001_11100110 : OUT <= 0;  //97 / 230 = 0
    16'b01100001_11100111 : OUT <= 0;  //97 / 231 = 0
    16'b01100001_11101000 : OUT <= 0;  //97 / 232 = 0
    16'b01100001_11101001 : OUT <= 0;  //97 / 233 = 0
    16'b01100001_11101010 : OUT <= 0;  //97 / 234 = 0
    16'b01100001_11101011 : OUT <= 0;  //97 / 235 = 0
    16'b01100001_11101100 : OUT <= 0;  //97 / 236 = 0
    16'b01100001_11101101 : OUT <= 0;  //97 / 237 = 0
    16'b01100001_11101110 : OUT <= 0;  //97 / 238 = 0
    16'b01100001_11101111 : OUT <= 0;  //97 / 239 = 0
    16'b01100001_11110000 : OUT <= 0;  //97 / 240 = 0
    16'b01100001_11110001 : OUT <= 0;  //97 / 241 = 0
    16'b01100001_11110010 : OUT <= 0;  //97 / 242 = 0
    16'b01100001_11110011 : OUT <= 0;  //97 / 243 = 0
    16'b01100001_11110100 : OUT <= 0;  //97 / 244 = 0
    16'b01100001_11110101 : OUT <= 0;  //97 / 245 = 0
    16'b01100001_11110110 : OUT <= 0;  //97 / 246 = 0
    16'b01100001_11110111 : OUT <= 0;  //97 / 247 = 0
    16'b01100001_11111000 : OUT <= 0;  //97 / 248 = 0
    16'b01100001_11111001 : OUT <= 0;  //97 / 249 = 0
    16'b01100001_11111010 : OUT <= 0;  //97 / 250 = 0
    16'b01100001_11111011 : OUT <= 0;  //97 / 251 = 0
    16'b01100001_11111100 : OUT <= 0;  //97 / 252 = 0
    16'b01100001_11111101 : OUT <= 0;  //97 / 253 = 0
    16'b01100001_11111110 : OUT <= 0;  //97 / 254 = 0
    16'b01100001_11111111 : OUT <= 0;  //97 / 255 = 0
    16'b01100010_00000000 : OUT <= 0;  //98 / 0 = 0
    16'b01100010_00000001 : OUT <= 98;  //98 / 1 = 98
    16'b01100010_00000010 : OUT <= 49;  //98 / 2 = 49
    16'b01100010_00000011 : OUT <= 32;  //98 / 3 = 32
    16'b01100010_00000100 : OUT <= 24;  //98 / 4 = 24
    16'b01100010_00000101 : OUT <= 19;  //98 / 5 = 19
    16'b01100010_00000110 : OUT <= 16;  //98 / 6 = 16
    16'b01100010_00000111 : OUT <= 14;  //98 / 7 = 14
    16'b01100010_00001000 : OUT <= 12;  //98 / 8 = 12
    16'b01100010_00001001 : OUT <= 10;  //98 / 9 = 10
    16'b01100010_00001010 : OUT <= 9;  //98 / 10 = 9
    16'b01100010_00001011 : OUT <= 8;  //98 / 11 = 8
    16'b01100010_00001100 : OUT <= 8;  //98 / 12 = 8
    16'b01100010_00001101 : OUT <= 7;  //98 / 13 = 7
    16'b01100010_00001110 : OUT <= 7;  //98 / 14 = 7
    16'b01100010_00001111 : OUT <= 6;  //98 / 15 = 6
    16'b01100010_00010000 : OUT <= 6;  //98 / 16 = 6
    16'b01100010_00010001 : OUT <= 5;  //98 / 17 = 5
    16'b01100010_00010010 : OUT <= 5;  //98 / 18 = 5
    16'b01100010_00010011 : OUT <= 5;  //98 / 19 = 5
    16'b01100010_00010100 : OUT <= 4;  //98 / 20 = 4
    16'b01100010_00010101 : OUT <= 4;  //98 / 21 = 4
    16'b01100010_00010110 : OUT <= 4;  //98 / 22 = 4
    16'b01100010_00010111 : OUT <= 4;  //98 / 23 = 4
    16'b01100010_00011000 : OUT <= 4;  //98 / 24 = 4
    16'b01100010_00011001 : OUT <= 3;  //98 / 25 = 3
    16'b01100010_00011010 : OUT <= 3;  //98 / 26 = 3
    16'b01100010_00011011 : OUT <= 3;  //98 / 27 = 3
    16'b01100010_00011100 : OUT <= 3;  //98 / 28 = 3
    16'b01100010_00011101 : OUT <= 3;  //98 / 29 = 3
    16'b01100010_00011110 : OUT <= 3;  //98 / 30 = 3
    16'b01100010_00011111 : OUT <= 3;  //98 / 31 = 3
    16'b01100010_00100000 : OUT <= 3;  //98 / 32 = 3
    16'b01100010_00100001 : OUT <= 2;  //98 / 33 = 2
    16'b01100010_00100010 : OUT <= 2;  //98 / 34 = 2
    16'b01100010_00100011 : OUT <= 2;  //98 / 35 = 2
    16'b01100010_00100100 : OUT <= 2;  //98 / 36 = 2
    16'b01100010_00100101 : OUT <= 2;  //98 / 37 = 2
    16'b01100010_00100110 : OUT <= 2;  //98 / 38 = 2
    16'b01100010_00100111 : OUT <= 2;  //98 / 39 = 2
    16'b01100010_00101000 : OUT <= 2;  //98 / 40 = 2
    16'b01100010_00101001 : OUT <= 2;  //98 / 41 = 2
    16'b01100010_00101010 : OUT <= 2;  //98 / 42 = 2
    16'b01100010_00101011 : OUT <= 2;  //98 / 43 = 2
    16'b01100010_00101100 : OUT <= 2;  //98 / 44 = 2
    16'b01100010_00101101 : OUT <= 2;  //98 / 45 = 2
    16'b01100010_00101110 : OUT <= 2;  //98 / 46 = 2
    16'b01100010_00101111 : OUT <= 2;  //98 / 47 = 2
    16'b01100010_00110000 : OUT <= 2;  //98 / 48 = 2
    16'b01100010_00110001 : OUT <= 2;  //98 / 49 = 2
    16'b01100010_00110010 : OUT <= 1;  //98 / 50 = 1
    16'b01100010_00110011 : OUT <= 1;  //98 / 51 = 1
    16'b01100010_00110100 : OUT <= 1;  //98 / 52 = 1
    16'b01100010_00110101 : OUT <= 1;  //98 / 53 = 1
    16'b01100010_00110110 : OUT <= 1;  //98 / 54 = 1
    16'b01100010_00110111 : OUT <= 1;  //98 / 55 = 1
    16'b01100010_00111000 : OUT <= 1;  //98 / 56 = 1
    16'b01100010_00111001 : OUT <= 1;  //98 / 57 = 1
    16'b01100010_00111010 : OUT <= 1;  //98 / 58 = 1
    16'b01100010_00111011 : OUT <= 1;  //98 / 59 = 1
    16'b01100010_00111100 : OUT <= 1;  //98 / 60 = 1
    16'b01100010_00111101 : OUT <= 1;  //98 / 61 = 1
    16'b01100010_00111110 : OUT <= 1;  //98 / 62 = 1
    16'b01100010_00111111 : OUT <= 1;  //98 / 63 = 1
    16'b01100010_01000000 : OUT <= 1;  //98 / 64 = 1
    16'b01100010_01000001 : OUT <= 1;  //98 / 65 = 1
    16'b01100010_01000010 : OUT <= 1;  //98 / 66 = 1
    16'b01100010_01000011 : OUT <= 1;  //98 / 67 = 1
    16'b01100010_01000100 : OUT <= 1;  //98 / 68 = 1
    16'b01100010_01000101 : OUT <= 1;  //98 / 69 = 1
    16'b01100010_01000110 : OUT <= 1;  //98 / 70 = 1
    16'b01100010_01000111 : OUT <= 1;  //98 / 71 = 1
    16'b01100010_01001000 : OUT <= 1;  //98 / 72 = 1
    16'b01100010_01001001 : OUT <= 1;  //98 / 73 = 1
    16'b01100010_01001010 : OUT <= 1;  //98 / 74 = 1
    16'b01100010_01001011 : OUT <= 1;  //98 / 75 = 1
    16'b01100010_01001100 : OUT <= 1;  //98 / 76 = 1
    16'b01100010_01001101 : OUT <= 1;  //98 / 77 = 1
    16'b01100010_01001110 : OUT <= 1;  //98 / 78 = 1
    16'b01100010_01001111 : OUT <= 1;  //98 / 79 = 1
    16'b01100010_01010000 : OUT <= 1;  //98 / 80 = 1
    16'b01100010_01010001 : OUT <= 1;  //98 / 81 = 1
    16'b01100010_01010010 : OUT <= 1;  //98 / 82 = 1
    16'b01100010_01010011 : OUT <= 1;  //98 / 83 = 1
    16'b01100010_01010100 : OUT <= 1;  //98 / 84 = 1
    16'b01100010_01010101 : OUT <= 1;  //98 / 85 = 1
    16'b01100010_01010110 : OUT <= 1;  //98 / 86 = 1
    16'b01100010_01010111 : OUT <= 1;  //98 / 87 = 1
    16'b01100010_01011000 : OUT <= 1;  //98 / 88 = 1
    16'b01100010_01011001 : OUT <= 1;  //98 / 89 = 1
    16'b01100010_01011010 : OUT <= 1;  //98 / 90 = 1
    16'b01100010_01011011 : OUT <= 1;  //98 / 91 = 1
    16'b01100010_01011100 : OUT <= 1;  //98 / 92 = 1
    16'b01100010_01011101 : OUT <= 1;  //98 / 93 = 1
    16'b01100010_01011110 : OUT <= 1;  //98 / 94 = 1
    16'b01100010_01011111 : OUT <= 1;  //98 / 95 = 1
    16'b01100010_01100000 : OUT <= 1;  //98 / 96 = 1
    16'b01100010_01100001 : OUT <= 1;  //98 / 97 = 1
    16'b01100010_01100010 : OUT <= 1;  //98 / 98 = 1
    16'b01100010_01100011 : OUT <= 0;  //98 / 99 = 0
    16'b01100010_01100100 : OUT <= 0;  //98 / 100 = 0
    16'b01100010_01100101 : OUT <= 0;  //98 / 101 = 0
    16'b01100010_01100110 : OUT <= 0;  //98 / 102 = 0
    16'b01100010_01100111 : OUT <= 0;  //98 / 103 = 0
    16'b01100010_01101000 : OUT <= 0;  //98 / 104 = 0
    16'b01100010_01101001 : OUT <= 0;  //98 / 105 = 0
    16'b01100010_01101010 : OUT <= 0;  //98 / 106 = 0
    16'b01100010_01101011 : OUT <= 0;  //98 / 107 = 0
    16'b01100010_01101100 : OUT <= 0;  //98 / 108 = 0
    16'b01100010_01101101 : OUT <= 0;  //98 / 109 = 0
    16'b01100010_01101110 : OUT <= 0;  //98 / 110 = 0
    16'b01100010_01101111 : OUT <= 0;  //98 / 111 = 0
    16'b01100010_01110000 : OUT <= 0;  //98 / 112 = 0
    16'b01100010_01110001 : OUT <= 0;  //98 / 113 = 0
    16'b01100010_01110010 : OUT <= 0;  //98 / 114 = 0
    16'b01100010_01110011 : OUT <= 0;  //98 / 115 = 0
    16'b01100010_01110100 : OUT <= 0;  //98 / 116 = 0
    16'b01100010_01110101 : OUT <= 0;  //98 / 117 = 0
    16'b01100010_01110110 : OUT <= 0;  //98 / 118 = 0
    16'b01100010_01110111 : OUT <= 0;  //98 / 119 = 0
    16'b01100010_01111000 : OUT <= 0;  //98 / 120 = 0
    16'b01100010_01111001 : OUT <= 0;  //98 / 121 = 0
    16'b01100010_01111010 : OUT <= 0;  //98 / 122 = 0
    16'b01100010_01111011 : OUT <= 0;  //98 / 123 = 0
    16'b01100010_01111100 : OUT <= 0;  //98 / 124 = 0
    16'b01100010_01111101 : OUT <= 0;  //98 / 125 = 0
    16'b01100010_01111110 : OUT <= 0;  //98 / 126 = 0
    16'b01100010_01111111 : OUT <= 0;  //98 / 127 = 0
    16'b01100010_10000000 : OUT <= 0;  //98 / 128 = 0
    16'b01100010_10000001 : OUT <= 0;  //98 / 129 = 0
    16'b01100010_10000010 : OUT <= 0;  //98 / 130 = 0
    16'b01100010_10000011 : OUT <= 0;  //98 / 131 = 0
    16'b01100010_10000100 : OUT <= 0;  //98 / 132 = 0
    16'b01100010_10000101 : OUT <= 0;  //98 / 133 = 0
    16'b01100010_10000110 : OUT <= 0;  //98 / 134 = 0
    16'b01100010_10000111 : OUT <= 0;  //98 / 135 = 0
    16'b01100010_10001000 : OUT <= 0;  //98 / 136 = 0
    16'b01100010_10001001 : OUT <= 0;  //98 / 137 = 0
    16'b01100010_10001010 : OUT <= 0;  //98 / 138 = 0
    16'b01100010_10001011 : OUT <= 0;  //98 / 139 = 0
    16'b01100010_10001100 : OUT <= 0;  //98 / 140 = 0
    16'b01100010_10001101 : OUT <= 0;  //98 / 141 = 0
    16'b01100010_10001110 : OUT <= 0;  //98 / 142 = 0
    16'b01100010_10001111 : OUT <= 0;  //98 / 143 = 0
    16'b01100010_10010000 : OUT <= 0;  //98 / 144 = 0
    16'b01100010_10010001 : OUT <= 0;  //98 / 145 = 0
    16'b01100010_10010010 : OUT <= 0;  //98 / 146 = 0
    16'b01100010_10010011 : OUT <= 0;  //98 / 147 = 0
    16'b01100010_10010100 : OUT <= 0;  //98 / 148 = 0
    16'b01100010_10010101 : OUT <= 0;  //98 / 149 = 0
    16'b01100010_10010110 : OUT <= 0;  //98 / 150 = 0
    16'b01100010_10010111 : OUT <= 0;  //98 / 151 = 0
    16'b01100010_10011000 : OUT <= 0;  //98 / 152 = 0
    16'b01100010_10011001 : OUT <= 0;  //98 / 153 = 0
    16'b01100010_10011010 : OUT <= 0;  //98 / 154 = 0
    16'b01100010_10011011 : OUT <= 0;  //98 / 155 = 0
    16'b01100010_10011100 : OUT <= 0;  //98 / 156 = 0
    16'b01100010_10011101 : OUT <= 0;  //98 / 157 = 0
    16'b01100010_10011110 : OUT <= 0;  //98 / 158 = 0
    16'b01100010_10011111 : OUT <= 0;  //98 / 159 = 0
    16'b01100010_10100000 : OUT <= 0;  //98 / 160 = 0
    16'b01100010_10100001 : OUT <= 0;  //98 / 161 = 0
    16'b01100010_10100010 : OUT <= 0;  //98 / 162 = 0
    16'b01100010_10100011 : OUT <= 0;  //98 / 163 = 0
    16'b01100010_10100100 : OUT <= 0;  //98 / 164 = 0
    16'b01100010_10100101 : OUT <= 0;  //98 / 165 = 0
    16'b01100010_10100110 : OUT <= 0;  //98 / 166 = 0
    16'b01100010_10100111 : OUT <= 0;  //98 / 167 = 0
    16'b01100010_10101000 : OUT <= 0;  //98 / 168 = 0
    16'b01100010_10101001 : OUT <= 0;  //98 / 169 = 0
    16'b01100010_10101010 : OUT <= 0;  //98 / 170 = 0
    16'b01100010_10101011 : OUT <= 0;  //98 / 171 = 0
    16'b01100010_10101100 : OUT <= 0;  //98 / 172 = 0
    16'b01100010_10101101 : OUT <= 0;  //98 / 173 = 0
    16'b01100010_10101110 : OUT <= 0;  //98 / 174 = 0
    16'b01100010_10101111 : OUT <= 0;  //98 / 175 = 0
    16'b01100010_10110000 : OUT <= 0;  //98 / 176 = 0
    16'b01100010_10110001 : OUT <= 0;  //98 / 177 = 0
    16'b01100010_10110010 : OUT <= 0;  //98 / 178 = 0
    16'b01100010_10110011 : OUT <= 0;  //98 / 179 = 0
    16'b01100010_10110100 : OUT <= 0;  //98 / 180 = 0
    16'b01100010_10110101 : OUT <= 0;  //98 / 181 = 0
    16'b01100010_10110110 : OUT <= 0;  //98 / 182 = 0
    16'b01100010_10110111 : OUT <= 0;  //98 / 183 = 0
    16'b01100010_10111000 : OUT <= 0;  //98 / 184 = 0
    16'b01100010_10111001 : OUT <= 0;  //98 / 185 = 0
    16'b01100010_10111010 : OUT <= 0;  //98 / 186 = 0
    16'b01100010_10111011 : OUT <= 0;  //98 / 187 = 0
    16'b01100010_10111100 : OUT <= 0;  //98 / 188 = 0
    16'b01100010_10111101 : OUT <= 0;  //98 / 189 = 0
    16'b01100010_10111110 : OUT <= 0;  //98 / 190 = 0
    16'b01100010_10111111 : OUT <= 0;  //98 / 191 = 0
    16'b01100010_11000000 : OUT <= 0;  //98 / 192 = 0
    16'b01100010_11000001 : OUT <= 0;  //98 / 193 = 0
    16'b01100010_11000010 : OUT <= 0;  //98 / 194 = 0
    16'b01100010_11000011 : OUT <= 0;  //98 / 195 = 0
    16'b01100010_11000100 : OUT <= 0;  //98 / 196 = 0
    16'b01100010_11000101 : OUT <= 0;  //98 / 197 = 0
    16'b01100010_11000110 : OUT <= 0;  //98 / 198 = 0
    16'b01100010_11000111 : OUT <= 0;  //98 / 199 = 0
    16'b01100010_11001000 : OUT <= 0;  //98 / 200 = 0
    16'b01100010_11001001 : OUT <= 0;  //98 / 201 = 0
    16'b01100010_11001010 : OUT <= 0;  //98 / 202 = 0
    16'b01100010_11001011 : OUT <= 0;  //98 / 203 = 0
    16'b01100010_11001100 : OUT <= 0;  //98 / 204 = 0
    16'b01100010_11001101 : OUT <= 0;  //98 / 205 = 0
    16'b01100010_11001110 : OUT <= 0;  //98 / 206 = 0
    16'b01100010_11001111 : OUT <= 0;  //98 / 207 = 0
    16'b01100010_11010000 : OUT <= 0;  //98 / 208 = 0
    16'b01100010_11010001 : OUT <= 0;  //98 / 209 = 0
    16'b01100010_11010010 : OUT <= 0;  //98 / 210 = 0
    16'b01100010_11010011 : OUT <= 0;  //98 / 211 = 0
    16'b01100010_11010100 : OUT <= 0;  //98 / 212 = 0
    16'b01100010_11010101 : OUT <= 0;  //98 / 213 = 0
    16'b01100010_11010110 : OUT <= 0;  //98 / 214 = 0
    16'b01100010_11010111 : OUT <= 0;  //98 / 215 = 0
    16'b01100010_11011000 : OUT <= 0;  //98 / 216 = 0
    16'b01100010_11011001 : OUT <= 0;  //98 / 217 = 0
    16'b01100010_11011010 : OUT <= 0;  //98 / 218 = 0
    16'b01100010_11011011 : OUT <= 0;  //98 / 219 = 0
    16'b01100010_11011100 : OUT <= 0;  //98 / 220 = 0
    16'b01100010_11011101 : OUT <= 0;  //98 / 221 = 0
    16'b01100010_11011110 : OUT <= 0;  //98 / 222 = 0
    16'b01100010_11011111 : OUT <= 0;  //98 / 223 = 0
    16'b01100010_11100000 : OUT <= 0;  //98 / 224 = 0
    16'b01100010_11100001 : OUT <= 0;  //98 / 225 = 0
    16'b01100010_11100010 : OUT <= 0;  //98 / 226 = 0
    16'b01100010_11100011 : OUT <= 0;  //98 / 227 = 0
    16'b01100010_11100100 : OUT <= 0;  //98 / 228 = 0
    16'b01100010_11100101 : OUT <= 0;  //98 / 229 = 0
    16'b01100010_11100110 : OUT <= 0;  //98 / 230 = 0
    16'b01100010_11100111 : OUT <= 0;  //98 / 231 = 0
    16'b01100010_11101000 : OUT <= 0;  //98 / 232 = 0
    16'b01100010_11101001 : OUT <= 0;  //98 / 233 = 0
    16'b01100010_11101010 : OUT <= 0;  //98 / 234 = 0
    16'b01100010_11101011 : OUT <= 0;  //98 / 235 = 0
    16'b01100010_11101100 : OUT <= 0;  //98 / 236 = 0
    16'b01100010_11101101 : OUT <= 0;  //98 / 237 = 0
    16'b01100010_11101110 : OUT <= 0;  //98 / 238 = 0
    16'b01100010_11101111 : OUT <= 0;  //98 / 239 = 0
    16'b01100010_11110000 : OUT <= 0;  //98 / 240 = 0
    16'b01100010_11110001 : OUT <= 0;  //98 / 241 = 0
    16'b01100010_11110010 : OUT <= 0;  //98 / 242 = 0
    16'b01100010_11110011 : OUT <= 0;  //98 / 243 = 0
    16'b01100010_11110100 : OUT <= 0;  //98 / 244 = 0
    16'b01100010_11110101 : OUT <= 0;  //98 / 245 = 0
    16'b01100010_11110110 : OUT <= 0;  //98 / 246 = 0
    16'b01100010_11110111 : OUT <= 0;  //98 / 247 = 0
    16'b01100010_11111000 : OUT <= 0;  //98 / 248 = 0
    16'b01100010_11111001 : OUT <= 0;  //98 / 249 = 0
    16'b01100010_11111010 : OUT <= 0;  //98 / 250 = 0
    16'b01100010_11111011 : OUT <= 0;  //98 / 251 = 0
    16'b01100010_11111100 : OUT <= 0;  //98 / 252 = 0
    16'b01100010_11111101 : OUT <= 0;  //98 / 253 = 0
    16'b01100010_11111110 : OUT <= 0;  //98 / 254 = 0
    16'b01100010_11111111 : OUT <= 0;  //98 / 255 = 0
    16'b01100011_00000000 : OUT <= 0;  //99 / 0 = 0
    16'b01100011_00000001 : OUT <= 99;  //99 / 1 = 99
    16'b01100011_00000010 : OUT <= 49;  //99 / 2 = 49
    16'b01100011_00000011 : OUT <= 33;  //99 / 3 = 33
    16'b01100011_00000100 : OUT <= 24;  //99 / 4 = 24
    16'b01100011_00000101 : OUT <= 19;  //99 / 5 = 19
    16'b01100011_00000110 : OUT <= 16;  //99 / 6 = 16
    16'b01100011_00000111 : OUT <= 14;  //99 / 7 = 14
    16'b01100011_00001000 : OUT <= 12;  //99 / 8 = 12
    16'b01100011_00001001 : OUT <= 11;  //99 / 9 = 11
    16'b01100011_00001010 : OUT <= 9;  //99 / 10 = 9
    16'b01100011_00001011 : OUT <= 9;  //99 / 11 = 9
    16'b01100011_00001100 : OUT <= 8;  //99 / 12 = 8
    16'b01100011_00001101 : OUT <= 7;  //99 / 13 = 7
    16'b01100011_00001110 : OUT <= 7;  //99 / 14 = 7
    16'b01100011_00001111 : OUT <= 6;  //99 / 15 = 6
    16'b01100011_00010000 : OUT <= 6;  //99 / 16 = 6
    16'b01100011_00010001 : OUT <= 5;  //99 / 17 = 5
    16'b01100011_00010010 : OUT <= 5;  //99 / 18 = 5
    16'b01100011_00010011 : OUT <= 5;  //99 / 19 = 5
    16'b01100011_00010100 : OUT <= 4;  //99 / 20 = 4
    16'b01100011_00010101 : OUT <= 4;  //99 / 21 = 4
    16'b01100011_00010110 : OUT <= 4;  //99 / 22 = 4
    16'b01100011_00010111 : OUT <= 4;  //99 / 23 = 4
    16'b01100011_00011000 : OUT <= 4;  //99 / 24 = 4
    16'b01100011_00011001 : OUT <= 3;  //99 / 25 = 3
    16'b01100011_00011010 : OUT <= 3;  //99 / 26 = 3
    16'b01100011_00011011 : OUT <= 3;  //99 / 27 = 3
    16'b01100011_00011100 : OUT <= 3;  //99 / 28 = 3
    16'b01100011_00011101 : OUT <= 3;  //99 / 29 = 3
    16'b01100011_00011110 : OUT <= 3;  //99 / 30 = 3
    16'b01100011_00011111 : OUT <= 3;  //99 / 31 = 3
    16'b01100011_00100000 : OUT <= 3;  //99 / 32 = 3
    16'b01100011_00100001 : OUT <= 3;  //99 / 33 = 3
    16'b01100011_00100010 : OUT <= 2;  //99 / 34 = 2
    16'b01100011_00100011 : OUT <= 2;  //99 / 35 = 2
    16'b01100011_00100100 : OUT <= 2;  //99 / 36 = 2
    16'b01100011_00100101 : OUT <= 2;  //99 / 37 = 2
    16'b01100011_00100110 : OUT <= 2;  //99 / 38 = 2
    16'b01100011_00100111 : OUT <= 2;  //99 / 39 = 2
    16'b01100011_00101000 : OUT <= 2;  //99 / 40 = 2
    16'b01100011_00101001 : OUT <= 2;  //99 / 41 = 2
    16'b01100011_00101010 : OUT <= 2;  //99 / 42 = 2
    16'b01100011_00101011 : OUT <= 2;  //99 / 43 = 2
    16'b01100011_00101100 : OUT <= 2;  //99 / 44 = 2
    16'b01100011_00101101 : OUT <= 2;  //99 / 45 = 2
    16'b01100011_00101110 : OUT <= 2;  //99 / 46 = 2
    16'b01100011_00101111 : OUT <= 2;  //99 / 47 = 2
    16'b01100011_00110000 : OUT <= 2;  //99 / 48 = 2
    16'b01100011_00110001 : OUT <= 2;  //99 / 49 = 2
    16'b01100011_00110010 : OUT <= 1;  //99 / 50 = 1
    16'b01100011_00110011 : OUT <= 1;  //99 / 51 = 1
    16'b01100011_00110100 : OUT <= 1;  //99 / 52 = 1
    16'b01100011_00110101 : OUT <= 1;  //99 / 53 = 1
    16'b01100011_00110110 : OUT <= 1;  //99 / 54 = 1
    16'b01100011_00110111 : OUT <= 1;  //99 / 55 = 1
    16'b01100011_00111000 : OUT <= 1;  //99 / 56 = 1
    16'b01100011_00111001 : OUT <= 1;  //99 / 57 = 1
    16'b01100011_00111010 : OUT <= 1;  //99 / 58 = 1
    16'b01100011_00111011 : OUT <= 1;  //99 / 59 = 1
    16'b01100011_00111100 : OUT <= 1;  //99 / 60 = 1
    16'b01100011_00111101 : OUT <= 1;  //99 / 61 = 1
    16'b01100011_00111110 : OUT <= 1;  //99 / 62 = 1
    16'b01100011_00111111 : OUT <= 1;  //99 / 63 = 1
    16'b01100011_01000000 : OUT <= 1;  //99 / 64 = 1
    16'b01100011_01000001 : OUT <= 1;  //99 / 65 = 1
    16'b01100011_01000010 : OUT <= 1;  //99 / 66 = 1
    16'b01100011_01000011 : OUT <= 1;  //99 / 67 = 1
    16'b01100011_01000100 : OUT <= 1;  //99 / 68 = 1
    16'b01100011_01000101 : OUT <= 1;  //99 / 69 = 1
    16'b01100011_01000110 : OUT <= 1;  //99 / 70 = 1
    16'b01100011_01000111 : OUT <= 1;  //99 / 71 = 1
    16'b01100011_01001000 : OUT <= 1;  //99 / 72 = 1
    16'b01100011_01001001 : OUT <= 1;  //99 / 73 = 1
    16'b01100011_01001010 : OUT <= 1;  //99 / 74 = 1
    16'b01100011_01001011 : OUT <= 1;  //99 / 75 = 1
    16'b01100011_01001100 : OUT <= 1;  //99 / 76 = 1
    16'b01100011_01001101 : OUT <= 1;  //99 / 77 = 1
    16'b01100011_01001110 : OUT <= 1;  //99 / 78 = 1
    16'b01100011_01001111 : OUT <= 1;  //99 / 79 = 1
    16'b01100011_01010000 : OUT <= 1;  //99 / 80 = 1
    16'b01100011_01010001 : OUT <= 1;  //99 / 81 = 1
    16'b01100011_01010010 : OUT <= 1;  //99 / 82 = 1
    16'b01100011_01010011 : OUT <= 1;  //99 / 83 = 1
    16'b01100011_01010100 : OUT <= 1;  //99 / 84 = 1
    16'b01100011_01010101 : OUT <= 1;  //99 / 85 = 1
    16'b01100011_01010110 : OUT <= 1;  //99 / 86 = 1
    16'b01100011_01010111 : OUT <= 1;  //99 / 87 = 1
    16'b01100011_01011000 : OUT <= 1;  //99 / 88 = 1
    16'b01100011_01011001 : OUT <= 1;  //99 / 89 = 1
    16'b01100011_01011010 : OUT <= 1;  //99 / 90 = 1
    16'b01100011_01011011 : OUT <= 1;  //99 / 91 = 1
    16'b01100011_01011100 : OUT <= 1;  //99 / 92 = 1
    16'b01100011_01011101 : OUT <= 1;  //99 / 93 = 1
    16'b01100011_01011110 : OUT <= 1;  //99 / 94 = 1
    16'b01100011_01011111 : OUT <= 1;  //99 / 95 = 1
    16'b01100011_01100000 : OUT <= 1;  //99 / 96 = 1
    16'b01100011_01100001 : OUT <= 1;  //99 / 97 = 1
    16'b01100011_01100010 : OUT <= 1;  //99 / 98 = 1
    16'b01100011_01100011 : OUT <= 1;  //99 / 99 = 1
    16'b01100011_01100100 : OUT <= 0;  //99 / 100 = 0
    16'b01100011_01100101 : OUT <= 0;  //99 / 101 = 0
    16'b01100011_01100110 : OUT <= 0;  //99 / 102 = 0
    16'b01100011_01100111 : OUT <= 0;  //99 / 103 = 0
    16'b01100011_01101000 : OUT <= 0;  //99 / 104 = 0
    16'b01100011_01101001 : OUT <= 0;  //99 / 105 = 0
    16'b01100011_01101010 : OUT <= 0;  //99 / 106 = 0
    16'b01100011_01101011 : OUT <= 0;  //99 / 107 = 0
    16'b01100011_01101100 : OUT <= 0;  //99 / 108 = 0
    16'b01100011_01101101 : OUT <= 0;  //99 / 109 = 0
    16'b01100011_01101110 : OUT <= 0;  //99 / 110 = 0
    16'b01100011_01101111 : OUT <= 0;  //99 / 111 = 0
    16'b01100011_01110000 : OUT <= 0;  //99 / 112 = 0
    16'b01100011_01110001 : OUT <= 0;  //99 / 113 = 0
    16'b01100011_01110010 : OUT <= 0;  //99 / 114 = 0
    16'b01100011_01110011 : OUT <= 0;  //99 / 115 = 0
    16'b01100011_01110100 : OUT <= 0;  //99 / 116 = 0
    16'b01100011_01110101 : OUT <= 0;  //99 / 117 = 0
    16'b01100011_01110110 : OUT <= 0;  //99 / 118 = 0
    16'b01100011_01110111 : OUT <= 0;  //99 / 119 = 0
    16'b01100011_01111000 : OUT <= 0;  //99 / 120 = 0
    16'b01100011_01111001 : OUT <= 0;  //99 / 121 = 0
    16'b01100011_01111010 : OUT <= 0;  //99 / 122 = 0
    16'b01100011_01111011 : OUT <= 0;  //99 / 123 = 0
    16'b01100011_01111100 : OUT <= 0;  //99 / 124 = 0
    16'b01100011_01111101 : OUT <= 0;  //99 / 125 = 0
    16'b01100011_01111110 : OUT <= 0;  //99 / 126 = 0
    16'b01100011_01111111 : OUT <= 0;  //99 / 127 = 0
    16'b01100011_10000000 : OUT <= 0;  //99 / 128 = 0
    16'b01100011_10000001 : OUT <= 0;  //99 / 129 = 0
    16'b01100011_10000010 : OUT <= 0;  //99 / 130 = 0
    16'b01100011_10000011 : OUT <= 0;  //99 / 131 = 0
    16'b01100011_10000100 : OUT <= 0;  //99 / 132 = 0
    16'b01100011_10000101 : OUT <= 0;  //99 / 133 = 0
    16'b01100011_10000110 : OUT <= 0;  //99 / 134 = 0
    16'b01100011_10000111 : OUT <= 0;  //99 / 135 = 0
    16'b01100011_10001000 : OUT <= 0;  //99 / 136 = 0
    16'b01100011_10001001 : OUT <= 0;  //99 / 137 = 0
    16'b01100011_10001010 : OUT <= 0;  //99 / 138 = 0
    16'b01100011_10001011 : OUT <= 0;  //99 / 139 = 0
    16'b01100011_10001100 : OUT <= 0;  //99 / 140 = 0
    16'b01100011_10001101 : OUT <= 0;  //99 / 141 = 0
    16'b01100011_10001110 : OUT <= 0;  //99 / 142 = 0
    16'b01100011_10001111 : OUT <= 0;  //99 / 143 = 0
    16'b01100011_10010000 : OUT <= 0;  //99 / 144 = 0
    16'b01100011_10010001 : OUT <= 0;  //99 / 145 = 0
    16'b01100011_10010010 : OUT <= 0;  //99 / 146 = 0
    16'b01100011_10010011 : OUT <= 0;  //99 / 147 = 0
    16'b01100011_10010100 : OUT <= 0;  //99 / 148 = 0
    16'b01100011_10010101 : OUT <= 0;  //99 / 149 = 0
    16'b01100011_10010110 : OUT <= 0;  //99 / 150 = 0
    16'b01100011_10010111 : OUT <= 0;  //99 / 151 = 0
    16'b01100011_10011000 : OUT <= 0;  //99 / 152 = 0
    16'b01100011_10011001 : OUT <= 0;  //99 / 153 = 0
    16'b01100011_10011010 : OUT <= 0;  //99 / 154 = 0
    16'b01100011_10011011 : OUT <= 0;  //99 / 155 = 0
    16'b01100011_10011100 : OUT <= 0;  //99 / 156 = 0
    16'b01100011_10011101 : OUT <= 0;  //99 / 157 = 0
    16'b01100011_10011110 : OUT <= 0;  //99 / 158 = 0
    16'b01100011_10011111 : OUT <= 0;  //99 / 159 = 0
    16'b01100011_10100000 : OUT <= 0;  //99 / 160 = 0
    16'b01100011_10100001 : OUT <= 0;  //99 / 161 = 0
    16'b01100011_10100010 : OUT <= 0;  //99 / 162 = 0
    16'b01100011_10100011 : OUT <= 0;  //99 / 163 = 0
    16'b01100011_10100100 : OUT <= 0;  //99 / 164 = 0
    16'b01100011_10100101 : OUT <= 0;  //99 / 165 = 0
    16'b01100011_10100110 : OUT <= 0;  //99 / 166 = 0
    16'b01100011_10100111 : OUT <= 0;  //99 / 167 = 0
    16'b01100011_10101000 : OUT <= 0;  //99 / 168 = 0
    16'b01100011_10101001 : OUT <= 0;  //99 / 169 = 0
    16'b01100011_10101010 : OUT <= 0;  //99 / 170 = 0
    16'b01100011_10101011 : OUT <= 0;  //99 / 171 = 0
    16'b01100011_10101100 : OUT <= 0;  //99 / 172 = 0
    16'b01100011_10101101 : OUT <= 0;  //99 / 173 = 0
    16'b01100011_10101110 : OUT <= 0;  //99 / 174 = 0
    16'b01100011_10101111 : OUT <= 0;  //99 / 175 = 0
    16'b01100011_10110000 : OUT <= 0;  //99 / 176 = 0
    16'b01100011_10110001 : OUT <= 0;  //99 / 177 = 0
    16'b01100011_10110010 : OUT <= 0;  //99 / 178 = 0
    16'b01100011_10110011 : OUT <= 0;  //99 / 179 = 0
    16'b01100011_10110100 : OUT <= 0;  //99 / 180 = 0
    16'b01100011_10110101 : OUT <= 0;  //99 / 181 = 0
    16'b01100011_10110110 : OUT <= 0;  //99 / 182 = 0
    16'b01100011_10110111 : OUT <= 0;  //99 / 183 = 0
    16'b01100011_10111000 : OUT <= 0;  //99 / 184 = 0
    16'b01100011_10111001 : OUT <= 0;  //99 / 185 = 0
    16'b01100011_10111010 : OUT <= 0;  //99 / 186 = 0
    16'b01100011_10111011 : OUT <= 0;  //99 / 187 = 0
    16'b01100011_10111100 : OUT <= 0;  //99 / 188 = 0
    16'b01100011_10111101 : OUT <= 0;  //99 / 189 = 0
    16'b01100011_10111110 : OUT <= 0;  //99 / 190 = 0
    16'b01100011_10111111 : OUT <= 0;  //99 / 191 = 0
    16'b01100011_11000000 : OUT <= 0;  //99 / 192 = 0
    16'b01100011_11000001 : OUT <= 0;  //99 / 193 = 0
    16'b01100011_11000010 : OUT <= 0;  //99 / 194 = 0
    16'b01100011_11000011 : OUT <= 0;  //99 / 195 = 0
    16'b01100011_11000100 : OUT <= 0;  //99 / 196 = 0
    16'b01100011_11000101 : OUT <= 0;  //99 / 197 = 0
    16'b01100011_11000110 : OUT <= 0;  //99 / 198 = 0
    16'b01100011_11000111 : OUT <= 0;  //99 / 199 = 0
    16'b01100011_11001000 : OUT <= 0;  //99 / 200 = 0
    16'b01100011_11001001 : OUT <= 0;  //99 / 201 = 0
    16'b01100011_11001010 : OUT <= 0;  //99 / 202 = 0
    16'b01100011_11001011 : OUT <= 0;  //99 / 203 = 0
    16'b01100011_11001100 : OUT <= 0;  //99 / 204 = 0
    16'b01100011_11001101 : OUT <= 0;  //99 / 205 = 0
    16'b01100011_11001110 : OUT <= 0;  //99 / 206 = 0
    16'b01100011_11001111 : OUT <= 0;  //99 / 207 = 0
    16'b01100011_11010000 : OUT <= 0;  //99 / 208 = 0
    16'b01100011_11010001 : OUT <= 0;  //99 / 209 = 0
    16'b01100011_11010010 : OUT <= 0;  //99 / 210 = 0
    16'b01100011_11010011 : OUT <= 0;  //99 / 211 = 0
    16'b01100011_11010100 : OUT <= 0;  //99 / 212 = 0
    16'b01100011_11010101 : OUT <= 0;  //99 / 213 = 0
    16'b01100011_11010110 : OUT <= 0;  //99 / 214 = 0
    16'b01100011_11010111 : OUT <= 0;  //99 / 215 = 0
    16'b01100011_11011000 : OUT <= 0;  //99 / 216 = 0
    16'b01100011_11011001 : OUT <= 0;  //99 / 217 = 0
    16'b01100011_11011010 : OUT <= 0;  //99 / 218 = 0
    16'b01100011_11011011 : OUT <= 0;  //99 / 219 = 0
    16'b01100011_11011100 : OUT <= 0;  //99 / 220 = 0
    16'b01100011_11011101 : OUT <= 0;  //99 / 221 = 0
    16'b01100011_11011110 : OUT <= 0;  //99 / 222 = 0
    16'b01100011_11011111 : OUT <= 0;  //99 / 223 = 0
    16'b01100011_11100000 : OUT <= 0;  //99 / 224 = 0
    16'b01100011_11100001 : OUT <= 0;  //99 / 225 = 0
    16'b01100011_11100010 : OUT <= 0;  //99 / 226 = 0
    16'b01100011_11100011 : OUT <= 0;  //99 / 227 = 0
    16'b01100011_11100100 : OUT <= 0;  //99 / 228 = 0
    16'b01100011_11100101 : OUT <= 0;  //99 / 229 = 0
    16'b01100011_11100110 : OUT <= 0;  //99 / 230 = 0
    16'b01100011_11100111 : OUT <= 0;  //99 / 231 = 0
    16'b01100011_11101000 : OUT <= 0;  //99 / 232 = 0
    16'b01100011_11101001 : OUT <= 0;  //99 / 233 = 0
    16'b01100011_11101010 : OUT <= 0;  //99 / 234 = 0
    16'b01100011_11101011 : OUT <= 0;  //99 / 235 = 0
    16'b01100011_11101100 : OUT <= 0;  //99 / 236 = 0
    16'b01100011_11101101 : OUT <= 0;  //99 / 237 = 0
    16'b01100011_11101110 : OUT <= 0;  //99 / 238 = 0
    16'b01100011_11101111 : OUT <= 0;  //99 / 239 = 0
    16'b01100011_11110000 : OUT <= 0;  //99 / 240 = 0
    16'b01100011_11110001 : OUT <= 0;  //99 / 241 = 0
    16'b01100011_11110010 : OUT <= 0;  //99 / 242 = 0
    16'b01100011_11110011 : OUT <= 0;  //99 / 243 = 0
    16'b01100011_11110100 : OUT <= 0;  //99 / 244 = 0
    16'b01100011_11110101 : OUT <= 0;  //99 / 245 = 0
    16'b01100011_11110110 : OUT <= 0;  //99 / 246 = 0
    16'b01100011_11110111 : OUT <= 0;  //99 / 247 = 0
    16'b01100011_11111000 : OUT <= 0;  //99 / 248 = 0
    16'b01100011_11111001 : OUT <= 0;  //99 / 249 = 0
    16'b01100011_11111010 : OUT <= 0;  //99 / 250 = 0
    16'b01100011_11111011 : OUT <= 0;  //99 / 251 = 0
    16'b01100011_11111100 : OUT <= 0;  //99 / 252 = 0
    16'b01100011_11111101 : OUT <= 0;  //99 / 253 = 0
    16'b01100011_11111110 : OUT <= 0;  //99 / 254 = 0
    16'b01100011_11111111 : OUT <= 0;  //99 / 255 = 0
    16'b01100100_00000000 : OUT <= 0;  //100 / 0 = 0
    16'b01100100_00000001 : OUT <= 100;  //100 / 1 = 100
    16'b01100100_00000010 : OUT <= 50;  //100 / 2 = 50
    16'b01100100_00000011 : OUT <= 33;  //100 / 3 = 33
    16'b01100100_00000100 : OUT <= 25;  //100 / 4 = 25
    16'b01100100_00000101 : OUT <= 20;  //100 / 5 = 20
    16'b01100100_00000110 : OUT <= 16;  //100 / 6 = 16
    16'b01100100_00000111 : OUT <= 14;  //100 / 7 = 14
    16'b01100100_00001000 : OUT <= 12;  //100 / 8 = 12
    16'b01100100_00001001 : OUT <= 11;  //100 / 9 = 11
    16'b01100100_00001010 : OUT <= 10;  //100 / 10 = 10
    16'b01100100_00001011 : OUT <= 9;  //100 / 11 = 9
    16'b01100100_00001100 : OUT <= 8;  //100 / 12 = 8
    16'b01100100_00001101 : OUT <= 7;  //100 / 13 = 7
    16'b01100100_00001110 : OUT <= 7;  //100 / 14 = 7
    16'b01100100_00001111 : OUT <= 6;  //100 / 15 = 6
    16'b01100100_00010000 : OUT <= 6;  //100 / 16 = 6
    16'b01100100_00010001 : OUT <= 5;  //100 / 17 = 5
    16'b01100100_00010010 : OUT <= 5;  //100 / 18 = 5
    16'b01100100_00010011 : OUT <= 5;  //100 / 19 = 5
    16'b01100100_00010100 : OUT <= 5;  //100 / 20 = 5
    16'b01100100_00010101 : OUT <= 4;  //100 / 21 = 4
    16'b01100100_00010110 : OUT <= 4;  //100 / 22 = 4
    16'b01100100_00010111 : OUT <= 4;  //100 / 23 = 4
    16'b01100100_00011000 : OUT <= 4;  //100 / 24 = 4
    16'b01100100_00011001 : OUT <= 4;  //100 / 25 = 4
    16'b01100100_00011010 : OUT <= 3;  //100 / 26 = 3
    16'b01100100_00011011 : OUT <= 3;  //100 / 27 = 3
    16'b01100100_00011100 : OUT <= 3;  //100 / 28 = 3
    16'b01100100_00011101 : OUT <= 3;  //100 / 29 = 3
    16'b01100100_00011110 : OUT <= 3;  //100 / 30 = 3
    16'b01100100_00011111 : OUT <= 3;  //100 / 31 = 3
    16'b01100100_00100000 : OUT <= 3;  //100 / 32 = 3
    16'b01100100_00100001 : OUT <= 3;  //100 / 33 = 3
    16'b01100100_00100010 : OUT <= 2;  //100 / 34 = 2
    16'b01100100_00100011 : OUT <= 2;  //100 / 35 = 2
    16'b01100100_00100100 : OUT <= 2;  //100 / 36 = 2
    16'b01100100_00100101 : OUT <= 2;  //100 / 37 = 2
    16'b01100100_00100110 : OUT <= 2;  //100 / 38 = 2
    16'b01100100_00100111 : OUT <= 2;  //100 / 39 = 2
    16'b01100100_00101000 : OUT <= 2;  //100 / 40 = 2
    16'b01100100_00101001 : OUT <= 2;  //100 / 41 = 2
    16'b01100100_00101010 : OUT <= 2;  //100 / 42 = 2
    16'b01100100_00101011 : OUT <= 2;  //100 / 43 = 2
    16'b01100100_00101100 : OUT <= 2;  //100 / 44 = 2
    16'b01100100_00101101 : OUT <= 2;  //100 / 45 = 2
    16'b01100100_00101110 : OUT <= 2;  //100 / 46 = 2
    16'b01100100_00101111 : OUT <= 2;  //100 / 47 = 2
    16'b01100100_00110000 : OUT <= 2;  //100 / 48 = 2
    16'b01100100_00110001 : OUT <= 2;  //100 / 49 = 2
    16'b01100100_00110010 : OUT <= 2;  //100 / 50 = 2
    16'b01100100_00110011 : OUT <= 1;  //100 / 51 = 1
    16'b01100100_00110100 : OUT <= 1;  //100 / 52 = 1
    16'b01100100_00110101 : OUT <= 1;  //100 / 53 = 1
    16'b01100100_00110110 : OUT <= 1;  //100 / 54 = 1
    16'b01100100_00110111 : OUT <= 1;  //100 / 55 = 1
    16'b01100100_00111000 : OUT <= 1;  //100 / 56 = 1
    16'b01100100_00111001 : OUT <= 1;  //100 / 57 = 1
    16'b01100100_00111010 : OUT <= 1;  //100 / 58 = 1
    16'b01100100_00111011 : OUT <= 1;  //100 / 59 = 1
    16'b01100100_00111100 : OUT <= 1;  //100 / 60 = 1
    16'b01100100_00111101 : OUT <= 1;  //100 / 61 = 1
    16'b01100100_00111110 : OUT <= 1;  //100 / 62 = 1
    16'b01100100_00111111 : OUT <= 1;  //100 / 63 = 1
    16'b01100100_01000000 : OUT <= 1;  //100 / 64 = 1
    16'b01100100_01000001 : OUT <= 1;  //100 / 65 = 1
    16'b01100100_01000010 : OUT <= 1;  //100 / 66 = 1
    16'b01100100_01000011 : OUT <= 1;  //100 / 67 = 1
    16'b01100100_01000100 : OUT <= 1;  //100 / 68 = 1
    16'b01100100_01000101 : OUT <= 1;  //100 / 69 = 1
    16'b01100100_01000110 : OUT <= 1;  //100 / 70 = 1
    16'b01100100_01000111 : OUT <= 1;  //100 / 71 = 1
    16'b01100100_01001000 : OUT <= 1;  //100 / 72 = 1
    16'b01100100_01001001 : OUT <= 1;  //100 / 73 = 1
    16'b01100100_01001010 : OUT <= 1;  //100 / 74 = 1
    16'b01100100_01001011 : OUT <= 1;  //100 / 75 = 1
    16'b01100100_01001100 : OUT <= 1;  //100 / 76 = 1
    16'b01100100_01001101 : OUT <= 1;  //100 / 77 = 1
    16'b01100100_01001110 : OUT <= 1;  //100 / 78 = 1
    16'b01100100_01001111 : OUT <= 1;  //100 / 79 = 1
    16'b01100100_01010000 : OUT <= 1;  //100 / 80 = 1
    16'b01100100_01010001 : OUT <= 1;  //100 / 81 = 1
    16'b01100100_01010010 : OUT <= 1;  //100 / 82 = 1
    16'b01100100_01010011 : OUT <= 1;  //100 / 83 = 1
    16'b01100100_01010100 : OUT <= 1;  //100 / 84 = 1
    16'b01100100_01010101 : OUT <= 1;  //100 / 85 = 1
    16'b01100100_01010110 : OUT <= 1;  //100 / 86 = 1
    16'b01100100_01010111 : OUT <= 1;  //100 / 87 = 1
    16'b01100100_01011000 : OUT <= 1;  //100 / 88 = 1
    16'b01100100_01011001 : OUT <= 1;  //100 / 89 = 1
    16'b01100100_01011010 : OUT <= 1;  //100 / 90 = 1
    16'b01100100_01011011 : OUT <= 1;  //100 / 91 = 1
    16'b01100100_01011100 : OUT <= 1;  //100 / 92 = 1
    16'b01100100_01011101 : OUT <= 1;  //100 / 93 = 1
    16'b01100100_01011110 : OUT <= 1;  //100 / 94 = 1
    16'b01100100_01011111 : OUT <= 1;  //100 / 95 = 1
    16'b01100100_01100000 : OUT <= 1;  //100 / 96 = 1
    16'b01100100_01100001 : OUT <= 1;  //100 / 97 = 1
    16'b01100100_01100010 : OUT <= 1;  //100 / 98 = 1
    16'b01100100_01100011 : OUT <= 1;  //100 / 99 = 1
    16'b01100100_01100100 : OUT <= 1;  //100 / 100 = 1
    16'b01100100_01100101 : OUT <= 0;  //100 / 101 = 0
    16'b01100100_01100110 : OUT <= 0;  //100 / 102 = 0
    16'b01100100_01100111 : OUT <= 0;  //100 / 103 = 0
    16'b01100100_01101000 : OUT <= 0;  //100 / 104 = 0
    16'b01100100_01101001 : OUT <= 0;  //100 / 105 = 0
    16'b01100100_01101010 : OUT <= 0;  //100 / 106 = 0
    16'b01100100_01101011 : OUT <= 0;  //100 / 107 = 0
    16'b01100100_01101100 : OUT <= 0;  //100 / 108 = 0
    16'b01100100_01101101 : OUT <= 0;  //100 / 109 = 0
    16'b01100100_01101110 : OUT <= 0;  //100 / 110 = 0
    16'b01100100_01101111 : OUT <= 0;  //100 / 111 = 0
    16'b01100100_01110000 : OUT <= 0;  //100 / 112 = 0
    16'b01100100_01110001 : OUT <= 0;  //100 / 113 = 0
    16'b01100100_01110010 : OUT <= 0;  //100 / 114 = 0
    16'b01100100_01110011 : OUT <= 0;  //100 / 115 = 0
    16'b01100100_01110100 : OUT <= 0;  //100 / 116 = 0
    16'b01100100_01110101 : OUT <= 0;  //100 / 117 = 0
    16'b01100100_01110110 : OUT <= 0;  //100 / 118 = 0
    16'b01100100_01110111 : OUT <= 0;  //100 / 119 = 0
    16'b01100100_01111000 : OUT <= 0;  //100 / 120 = 0
    16'b01100100_01111001 : OUT <= 0;  //100 / 121 = 0
    16'b01100100_01111010 : OUT <= 0;  //100 / 122 = 0
    16'b01100100_01111011 : OUT <= 0;  //100 / 123 = 0
    16'b01100100_01111100 : OUT <= 0;  //100 / 124 = 0
    16'b01100100_01111101 : OUT <= 0;  //100 / 125 = 0
    16'b01100100_01111110 : OUT <= 0;  //100 / 126 = 0
    16'b01100100_01111111 : OUT <= 0;  //100 / 127 = 0
    16'b01100100_10000000 : OUT <= 0;  //100 / 128 = 0
    16'b01100100_10000001 : OUT <= 0;  //100 / 129 = 0
    16'b01100100_10000010 : OUT <= 0;  //100 / 130 = 0
    16'b01100100_10000011 : OUT <= 0;  //100 / 131 = 0
    16'b01100100_10000100 : OUT <= 0;  //100 / 132 = 0
    16'b01100100_10000101 : OUT <= 0;  //100 / 133 = 0
    16'b01100100_10000110 : OUT <= 0;  //100 / 134 = 0
    16'b01100100_10000111 : OUT <= 0;  //100 / 135 = 0
    16'b01100100_10001000 : OUT <= 0;  //100 / 136 = 0
    16'b01100100_10001001 : OUT <= 0;  //100 / 137 = 0
    16'b01100100_10001010 : OUT <= 0;  //100 / 138 = 0
    16'b01100100_10001011 : OUT <= 0;  //100 / 139 = 0
    16'b01100100_10001100 : OUT <= 0;  //100 / 140 = 0
    16'b01100100_10001101 : OUT <= 0;  //100 / 141 = 0
    16'b01100100_10001110 : OUT <= 0;  //100 / 142 = 0
    16'b01100100_10001111 : OUT <= 0;  //100 / 143 = 0
    16'b01100100_10010000 : OUT <= 0;  //100 / 144 = 0
    16'b01100100_10010001 : OUT <= 0;  //100 / 145 = 0
    16'b01100100_10010010 : OUT <= 0;  //100 / 146 = 0
    16'b01100100_10010011 : OUT <= 0;  //100 / 147 = 0
    16'b01100100_10010100 : OUT <= 0;  //100 / 148 = 0
    16'b01100100_10010101 : OUT <= 0;  //100 / 149 = 0
    16'b01100100_10010110 : OUT <= 0;  //100 / 150 = 0
    16'b01100100_10010111 : OUT <= 0;  //100 / 151 = 0
    16'b01100100_10011000 : OUT <= 0;  //100 / 152 = 0
    16'b01100100_10011001 : OUT <= 0;  //100 / 153 = 0
    16'b01100100_10011010 : OUT <= 0;  //100 / 154 = 0
    16'b01100100_10011011 : OUT <= 0;  //100 / 155 = 0
    16'b01100100_10011100 : OUT <= 0;  //100 / 156 = 0
    16'b01100100_10011101 : OUT <= 0;  //100 / 157 = 0
    16'b01100100_10011110 : OUT <= 0;  //100 / 158 = 0
    16'b01100100_10011111 : OUT <= 0;  //100 / 159 = 0
    16'b01100100_10100000 : OUT <= 0;  //100 / 160 = 0
    16'b01100100_10100001 : OUT <= 0;  //100 / 161 = 0
    16'b01100100_10100010 : OUT <= 0;  //100 / 162 = 0
    16'b01100100_10100011 : OUT <= 0;  //100 / 163 = 0
    16'b01100100_10100100 : OUT <= 0;  //100 / 164 = 0
    16'b01100100_10100101 : OUT <= 0;  //100 / 165 = 0
    16'b01100100_10100110 : OUT <= 0;  //100 / 166 = 0
    16'b01100100_10100111 : OUT <= 0;  //100 / 167 = 0
    16'b01100100_10101000 : OUT <= 0;  //100 / 168 = 0
    16'b01100100_10101001 : OUT <= 0;  //100 / 169 = 0
    16'b01100100_10101010 : OUT <= 0;  //100 / 170 = 0
    16'b01100100_10101011 : OUT <= 0;  //100 / 171 = 0
    16'b01100100_10101100 : OUT <= 0;  //100 / 172 = 0
    16'b01100100_10101101 : OUT <= 0;  //100 / 173 = 0
    16'b01100100_10101110 : OUT <= 0;  //100 / 174 = 0
    16'b01100100_10101111 : OUT <= 0;  //100 / 175 = 0
    16'b01100100_10110000 : OUT <= 0;  //100 / 176 = 0
    16'b01100100_10110001 : OUT <= 0;  //100 / 177 = 0
    16'b01100100_10110010 : OUT <= 0;  //100 / 178 = 0
    16'b01100100_10110011 : OUT <= 0;  //100 / 179 = 0
    16'b01100100_10110100 : OUT <= 0;  //100 / 180 = 0
    16'b01100100_10110101 : OUT <= 0;  //100 / 181 = 0
    16'b01100100_10110110 : OUT <= 0;  //100 / 182 = 0
    16'b01100100_10110111 : OUT <= 0;  //100 / 183 = 0
    16'b01100100_10111000 : OUT <= 0;  //100 / 184 = 0
    16'b01100100_10111001 : OUT <= 0;  //100 / 185 = 0
    16'b01100100_10111010 : OUT <= 0;  //100 / 186 = 0
    16'b01100100_10111011 : OUT <= 0;  //100 / 187 = 0
    16'b01100100_10111100 : OUT <= 0;  //100 / 188 = 0
    16'b01100100_10111101 : OUT <= 0;  //100 / 189 = 0
    16'b01100100_10111110 : OUT <= 0;  //100 / 190 = 0
    16'b01100100_10111111 : OUT <= 0;  //100 / 191 = 0
    16'b01100100_11000000 : OUT <= 0;  //100 / 192 = 0
    16'b01100100_11000001 : OUT <= 0;  //100 / 193 = 0
    16'b01100100_11000010 : OUT <= 0;  //100 / 194 = 0
    16'b01100100_11000011 : OUT <= 0;  //100 / 195 = 0
    16'b01100100_11000100 : OUT <= 0;  //100 / 196 = 0
    16'b01100100_11000101 : OUT <= 0;  //100 / 197 = 0
    16'b01100100_11000110 : OUT <= 0;  //100 / 198 = 0
    16'b01100100_11000111 : OUT <= 0;  //100 / 199 = 0
    16'b01100100_11001000 : OUT <= 0;  //100 / 200 = 0
    16'b01100100_11001001 : OUT <= 0;  //100 / 201 = 0
    16'b01100100_11001010 : OUT <= 0;  //100 / 202 = 0
    16'b01100100_11001011 : OUT <= 0;  //100 / 203 = 0
    16'b01100100_11001100 : OUT <= 0;  //100 / 204 = 0
    16'b01100100_11001101 : OUT <= 0;  //100 / 205 = 0
    16'b01100100_11001110 : OUT <= 0;  //100 / 206 = 0
    16'b01100100_11001111 : OUT <= 0;  //100 / 207 = 0
    16'b01100100_11010000 : OUT <= 0;  //100 / 208 = 0
    16'b01100100_11010001 : OUT <= 0;  //100 / 209 = 0
    16'b01100100_11010010 : OUT <= 0;  //100 / 210 = 0
    16'b01100100_11010011 : OUT <= 0;  //100 / 211 = 0
    16'b01100100_11010100 : OUT <= 0;  //100 / 212 = 0
    16'b01100100_11010101 : OUT <= 0;  //100 / 213 = 0
    16'b01100100_11010110 : OUT <= 0;  //100 / 214 = 0
    16'b01100100_11010111 : OUT <= 0;  //100 / 215 = 0
    16'b01100100_11011000 : OUT <= 0;  //100 / 216 = 0
    16'b01100100_11011001 : OUT <= 0;  //100 / 217 = 0
    16'b01100100_11011010 : OUT <= 0;  //100 / 218 = 0
    16'b01100100_11011011 : OUT <= 0;  //100 / 219 = 0
    16'b01100100_11011100 : OUT <= 0;  //100 / 220 = 0
    16'b01100100_11011101 : OUT <= 0;  //100 / 221 = 0
    16'b01100100_11011110 : OUT <= 0;  //100 / 222 = 0
    16'b01100100_11011111 : OUT <= 0;  //100 / 223 = 0
    16'b01100100_11100000 : OUT <= 0;  //100 / 224 = 0
    16'b01100100_11100001 : OUT <= 0;  //100 / 225 = 0
    16'b01100100_11100010 : OUT <= 0;  //100 / 226 = 0
    16'b01100100_11100011 : OUT <= 0;  //100 / 227 = 0
    16'b01100100_11100100 : OUT <= 0;  //100 / 228 = 0
    16'b01100100_11100101 : OUT <= 0;  //100 / 229 = 0
    16'b01100100_11100110 : OUT <= 0;  //100 / 230 = 0
    16'b01100100_11100111 : OUT <= 0;  //100 / 231 = 0
    16'b01100100_11101000 : OUT <= 0;  //100 / 232 = 0
    16'b01100100_11101001 : OUT <= 0;  //100 / 233 = 0
    16'b01100100_11101010 : OUT <= 0;  //100 / 234 = 0
    16'b01100100_11101011 : OUT <= 0;  //100 / 235 = 0
    16'b01100100_11101100 : OUT <= 0;  //100 / 236 = 0
    16'b01100100_11101101 : OUT <= 0;  //100 / 237 = 0
    16'b01100100_11101110 : OUT <= 0;  //100 / 238 = 0
    16'b01100100_11101111 : OUT <= 0;  //100 / 239 = 0
    16'b01100100_11110000 : OUT <= 0;  //100 / 240 = 0
    16'b01100100_11110001 : OUT <= 0;  //100 / 241 = 0
    16'b01100100_11110010 : OUT <= 0;  //100 / 242 = 0
    16'b01100100_11110011 : OUT <= 0;  //100 / 243 = 0
    16'b01100100_11110100 : OUT <= 0;  //100 / 244 = 0
    16'b01100100_11110101 : OUT <= 0;  //100 / 245 = 0
    16'b01100100_11110110 : OUT <= 0;  //100 / 246 = 0
    16'b01100100_11110111 : OUT <= 0;  //100 / 247 = 0
    16'b01100100_11111000 : OUT <= 0;  //100 / 248 = 0
    16'b01100100_11111001 : OUT <= 0;  //100 / 249 = 0
    16'b01100100_11111010 : OUT <= 0;  //100 / 250 = 0
    16'b01100100_11111011 : OUT <= 0;  //100 / 251 = 0
    16'b01100100_11111100 : OUT <= 0;  //100 / 252 = 0
    16'b01100100_11111101 : OUT <= 0;  //100 / 253 = 0
    16'b01100100_11111110 : OUT <= 0;  //100 / 254 = 0
    16'b01100100_11111111 : OUT <= 0;  //100 / 255 = 0
    16'b01100101_00000000 : OUT <= 0;  //101 / 0 = 0
    16'b01100101_00000001 : OUT <= 101;  //101 / 1 = 101
    16'b01100101_00000010 : OUT <= 50;  //101 / 2 = 50
    16'b01100101_00000011 : OUT <= 33;  //101 / 3 = 33
    16'b01100101_00000100 : OUT <= 25;  //101 / 4 = 25
    16'b01100101_00000101 : OUT <= 20;  //101 / 5 = 20
    16'b01100101_00000110 : OUT <= 16;  //101 / 6 = 16
    16'b01100101_00000111 : OUT <= 14;  //101 / 7 = 14
    16'b01100101_00001000 : OUT <= 12;  //101 / 8 = 12
    16'b01100101_00001001 : OUT <= 11;  //101 / 9 = 11
    16'b01100101_00001010 : OUT <= 10;  //101 / 10 = 10
    16'b01100101_00001011 : OUT <= 9;  //101 / 11 = 9
    16'b01100101_00001100 : OUT <= 8;  //101 / 12 = 8
    16'b01100101_00001101 : OUT <= 7;  //101 / 13 = 7
    16'b01100101_00001110 : OUT <= 7;  //101 / 14 = 7
    16'b01100101_00001111 : OUT <= 6;  //101 / 15 = 6
    16'b01100101_00010000 : OUT <= 6;  //101 / 16 = 6
    16'b01100101_00010001 : OUT <= 5;  //101 / 17 = 5
    16'b01100101_00010010 : OUT <= 5;  //101 / 18 = 5
    16'b01100101_00010011 : OUT <= 5;  //101 / 19 = 5
    16'b01100101_00010100 : OUT <= 5;  //101 / 20 = 5
    16'b01100101_00010101 : OUT <= 4;  //101 / 21 = 4
    16'b01100101_00010110 : OUT <= 4;  //101 / 22 = 4
    16'b01100101_00010111 : OUT <= 4;  //101 / 23 = 4
    16'b01100101_00011000 : OUT <= 4;  //101 / 24 = 4
    16'b01100101_00011001 : OUT <= 4;  //101 / 25 = 4
    16'b01100101_00011010 : OUT <= 3;  //101 / 26 = 3
    16'b01100101_00011011 : OUT <= 3;  //101 / 27 = 3
    16'b01100101_00011100 : OUT <= 3;  //101 / 28 = 3
    16'b01100101_00011101 : OUT <= 3;  //101 / 29 = 3
    16'b01100101_00011110 : OUT <= 3;  //101 / 30 = 3
    16'b01100101_00011111 : OUT <= 3;  //101 / 31 = 3
    16'b01100101_00100000 : OUT <= 3;  //101 / 32 = 3
    16'b01100101_00100001 : OUT <= 3;  //101 / 33 = 3
    16'b01100101_00100010 : OUT <= 2;  //101 / 34 = 2
    16'b01100101_00100011 : OUT <= 2;  //101 / 35 = 2
    16'b01100101_00100100 : OUT <= 2;  //101 / 36 = 2
    16'b01100101_00100101 : OUT <= 2;  //101 / 37 = 2
    16'b01100101_00100110 : OUT <= 2;  //101 / 38 = 2
    16'b01100101_00100111 : OUT <= 2;  //101 / 39 = 2
    16'b01100101_00101000 : OUT <= 2;  //101 / 40 = 2
    16'b01100101_00101001 : OUT <= 2;  //101 / 41 = 2
    16'b01100101_00101010 : OUT <= 2;  //101 / 42 = 2
    16'b01100101_00101011 : OUT <= 2;  //101 / 43 = 2
    16'b01100101_00101100 : OUT <= 2;  //101 / 44 = 2
    16'b01100101_00101101 : OUT <= 2;  //101 / 45 = 2
    16'b01100101_00101110 : OUT <= 2;  //101 / 46 = 2
    16'b01100101_00101111 : OUT <= 2;  //101 / 47 = 2
    16'b01100101_00110000 : OUT <= 2;  //101 / 48 = 2
    16'b01100101_00110001 : OUT <= 2;  //101 / 49 = 2
    16'b01100101_00110010 : OUT <= 2;  //101 / 50 = 2
    16'b01100101_00110011 : OUT <= 1;  //101 / 51 = 1
    16'b01100101_00110100 : OUT <= 1;  //101 / 52 = 1
    16'b01100101_00110101 : OUT <= 1;  //101 / 53 = 1
    16'b01100101_00110110 : OUT <= 1;  //101 / 54 = 1
    16'b01100101_00110111 : OUT <= 1;  //101 / 55 = 1
    16'b01100101_00111000 : OUT <= 1;  //101 / 56 = 1
    16'b01100101_00111001 : OUT <= 1;  //101 / 57 = 1
    16'b01100101_00111010 : OUT <= 1;  //101 / 58 = 1
    16'b01100101_00111011 : OUT <= 1;  //101 / 59 = 1
    16'b01100101_00111100 : OUT <= 1;  //101 / 60 = 1
    16'b01100101_00111101 : OUT <= 1;  //101 / 61 = 1
    16'b01100101_00111110 : OUT <= 1;  //101 / 62 = 1
    16'b01100101_00111111 : OUT <= 1;  //101 / 63 = 1
    16'b01100101_01000000 : OUT <= 1;  //101 / 64 = 1
    16'b01100101_01000001 : OUT <= 1;  //101 / 65 = 1
    16'b01100101_01000010 : OUT <= 1;  //101 / 66 = 1
    16'b01100101_01000011 : OUT <= 1;  //101 / 67 = 1
    16'b01100101_01000100 : OUT <= 1;  //101 / 68 = 1
    16'b01100101_01000101 : OUT <= 1;  //101 / 69 = 1
    16'b01100101_01000110 : OUT <= 1;  //101 / 70 = 1
    16'b01100101_01000111 : OUT <= 1;  //101 / 71 = 1
    16'b01100101_01001000 : OUT <= 1;  //101 / 72 = 1
    16'b01100101_01001001 : OUT <= 1;  //101 / 73 = 1
    16'b01100101_01001010 : OUT <= 1;  //101 / 74 = 1
    16'b01100101_01001011 : OUT <= 1;  //101 / 75 = 1
    16'b01100101_01001100 : OUT <= 1;  //101 / 76 = 1
    16'b01100101_01001101 : OUT <= 1;  //101 / 77 = 1
    16'b01100101_01001110 : OUT <= 1;  //101 / 78 = 1
    16'b01100101_01001111 : OUT <= 1;  //101 / 79 = 1
    16'b01100101_01010000 : OUT <= 1;  //101 / 80 = 1
    16'b01100101_01010001 : OUT <= 1;  //101 / 81 = 1
    16'b01100101_01010010 : OUT <= 1;  //101 / 82 = 1
    16'b01100101_01010011 : OUT <= 1;  //101 / 83 = 1
    16'b01100101_01010100 : OUT <= 1;  //101 / 84 = 1
    16'b01100101_01010101 : OUT <= 1;  //101 / 85 = 1
    16'b01100101_01010110 : OUT <= 1;  //101 / 86 = 1
    16'b01100101_01010111 : OUT <= 1;  //101 / 87 = 1
    16'b01100101_01011000 : OUT <= 1;  //101 / 88 = 1
    16'b01100101_01011001 : OUT <= 1;  //101 / 89 = 1
    16'b01100101_01011010 : OUT <= 1;  //101 / 90 = 1
    16'b01100101_01011011 : OUT <= 1;  //101 / 91 = 1
    16'b01100101_01011100 : OUT <= 1;  //101 / 92 = 1
    16'b01100101_01011101 : OUT <= 1;  //101 / 93 = 1
    16'b01100101_01011110 : OUT <= 1;  //101 / 94 = 1
    16'b01100101_01011111 : OUT <= 1;  //101 / 95 = 1
    16'b01100101_01100000 : OUT <= 1;  //101 / 96 = 1
    16'b01100101_01100001 : OUT <= 1;  //101 / 97 = 1
    16'b01100101_01100010 : OUT <= 1;  //101 / 98 = 1
    16'b01100101_01100011 : OUT <= 1;  //101 / 99 = 1
    16'b01100101_01100100 : OUT <= 1;  //101 / 100 = 1
    16'b01100101_01100101 : OUT <= 1;  //101 / 101 = 1
    16'b01100101_01100110 : OUT <= 0;  //101 / 102 = 0
    16'b01100101_01100111 : OUT <= 0;  //101 / 103 = 0
    16'b01100101_01101000 : OUT <= 0;  //101 / 104 = 0
    16'b01100101_01101001 : OUT <= 0;  //101 / 105 = 0
    16'b01100101_01101010 : OUT <= 0;  //101 / 106 = 0
    16'b01100101_01101011 : OUT <= 0;  //101 / 107 = 0
    16'b01100101_01101100 : OUT <= 0;  //101 / 108 = 0
    16'b01100101_01101101 : OUT <= 0;  //101 / 109 = 0
    16'b01100101_01101110 : OUT <= 0;  //101 / 110 = 0
    16'b01100101_01101111 : OUT <= 0;  //101 / 111 = 0
    16'b01100101_01110000 : OUT <= 0;  //101 / 112 = 0
    16'b01100101_01110001 : OUT <= 0;  //101 / 113 = 0
    16'b01100101_01110010 : OUT <= 0;  //101 / 114 = 0
    16'b01100101_01110011 : OUT <= 0;  //101 / 115 = 0
    16'b01100101_01110100 : OUT <= 0;  //101 / 116 = 0
    16'b01100101_01110101 : OUT <= 0;  //101 / 117 = 0
    16'b01100101_01110110 : OUT <= 0;  //101 / 118 = 0
    16'b01100101_01110111 : OUT <= 0;  //101 / 119 = 0
    16'b01100101_01111000 : OUT <= 0;  //101 / 120 = 0
    16'b01100101_01111001 : OUT <= 0;  //101 / 121 = 0
    16'b01100101_01111010 : OUT <= 0;  //101 / 122 = 0
    16'b01100101_01111011 : OUT <= 0;  //101 / 123 = 0
    16'b01100101_01111100 : OUT <= 0;  //101 / 124 = 0
    16'b01100101_01111101 : OUT <= 0;  //101 / 125 = 0
    16'b01100101_01111110 : OUT <= 0;  //101 / 126 = 0
    16'b01100101_01111111 : OUT <= 0;  //101 / 127 = 0
    16'b01100101_10000000 : OUT <= 0;  //101 / 128 = 0
    16'b01100101_10000001 : OUT <= 0;  //101 / 129 = 0
    16'b01100101_10000010 : OUT <= 0;  //101 / 130 = 0
    16'b01100101_10000011 : OUT <= 0;  //101 / 131 = 0
    16'b01100101_10000100 : OUT <= 0;  //101 / 132 = 0
    16'b01100101_10000101 : OUT <= 0;  //101 / 133 = 0
    16'b01100101_10000110 : OUT <= 0;  //101 / 134 = 0
    16'b01100101_10000111 : OUT <= 0;  //101 / 135 = 0
    16'b01100101_10001000 : OUT <= 0;  //101 / 136 = 0
    16'b01100101_10001001 : OUT <= 0;  //101 / 137 = 0
    16'b01100101_10001010 : OUT <= 0;  //101 / 138 = 0
    16'b01100101_10001011 : OUT <= 0;  //101 / 139 = 0
    16'b01100101_10001100 : OUT <= 0;  //101 / 140 = 0
    16'b01100101_10001101 : OUT <= 0;  //101 / 141 = 0
    16'b01100101_10001110 : OUT <= 0;  //101 / 142 = 0
    16'b01100101_10001111 : OUT <= 0;  //101 / 143 = 0
    16'b01100101_10010000 : OUT <= 0;  //101 / 144 = 0
    16'b01100101_10010001 : OUT <= 0;  //101 / 145 = 0
    16'b01100101_10010010 : OUT <= 0;  //101 / 146 = 0
    16'b01100101_10010011 : OUT <= 0;  //101 / 147 = 0
    16'b01100101_10010100 : OUT <= 0;  //101 / 148 = 0
    16'b01100101_10010101 : OUT <= 0;  //101 / 149 = 0
    16'b01100101_10010110 : OUT <= 0;  //101 / 150 = 0
    16'b01100101_10010111 : OUT <= 0;  //101 / 151 = 0
    16'b01100101_10011000 : OUT <= 0;  //101 / 152 = 0
    16'b01100101_10011001 : OUT <= 0;  //101 / 153 = 0
    16'b01100101_10011010 : OUT <= 0;  //101 / 154 = 0
    16'b01100101_10011011 : OUT <= 0;  //101 / 155 = 0
    16'b01100101_10011100 : OUT <= 0;  //101 / 156 = 0
    16'b01100101_10011101 : OUT <= 0;  //101 / 157 = 0
    16'b01100101_10011110 : OUT <= 0;  //101 / 158 = 0
    16'b01100101_10011111 : OUT <= 0;  //101 / 159 = 0
    16'b01100101_10100000 : OUT <= 0;  //101 / 160 = 0
    16'b01100101_10100001 : OUT <= 0;  //101 / 161 = 0
    16'b01100101_10100010 : OUT <= 0;  //101 / 162 = 0
    16'b01100101_10100011 : OUT <= 0;  //101 / 163 = 0
    16'b01100101_10100100 : OUT <= 0;  //101 / 164 = 0
    16'b01100101_10100101 : OUT <= 0;  //101 / 165 = 0
    16'b01100101_10100110 : OUT <= 0;  //101 / 166 = 0
    16'b01100101_10100111 : OUT <= 0;  //101 / 167 = 0
    16'b01100101_10101000 : OUT <= 0;  //101 / 168 = 0
    16'b01100101_10101001 : OUT <= 0;  //101 / 169 = 0
    16'b01100101_10101010 : OUT <= 0;  //101 / 170 = 0
    16'b01100101_10101011 : OUT <= 0;  //101 / 171 = 0
    16'b01100101_10101100 : OUT <= 0;  //101 / 172 = 0
    16'b01100101_10101101 : OUT <= 0;  //101 / 173 = 0
    16'b01100101_10101110 : OUT <= 0;  //101 / 174 = 0
    16'b01100101_10101111 : OUT <= 0;  //101 / 175 = 0
    16'b01100101_10110000 : OUT <= 0;  //101 / 176 = 0
    16'b01100101_10110001 : OUT <= 0;  //101 / 177 = 0
    16'b01100101_10110010 : OUT <= 0;  //101 / 178 = 0
    16'b01100101_10110011 : OUT <= 0;  //101 / 179 = 0
    16'b01100101_10110100 : OUT <= 0;  //101 / 180 = 0
    16'b01100101_10110101 : OUT <= 0;  //101 / 181 = 0
    16'b01100101_10110110 : OUT <= 0;  //101 / 182 = 0
    16'b01100101_10110111 : OUT <= 0;  //101 / 183 = 0
    16'b01100101_10111000 : OUT <= 0;  //101 / 184 = 0
    16'b01100101_10111001 : OUT <= 0;  //101 / 185 = 0
    16'b01100101_10111010 : OUT <= 0;  //101 / 186 = 0
    16'b01100101_10111011 : OUT <= 0;  //101 / 187 = 0
    16'b01100101_10111100 : OUT <= 0;  //101 / 188 = 0
    16'b01100101_10111101 : OUT <= 0;  //101 / 189 = 0
    16'b01100101_10111110 : OUT <= 0;  //101 / 190 = 0
    16'b01100101_10111111 : OUT <= 0;  //101 / 191 = 0
    16'b01100101_11000000 : OUT <= 0;  //101 / 192 = 0
    16'b01100101_11000001 : OUT <= 0;  //101 / 193 = 0
    16'b01100101_11000010 : OUT <= 0;  //101 / 194 = 0
    16'b01100101_11000011 : OUT <= 0;  //101 / 195 = 0
    16'b01100101_11000100 : OUT <= 0;  //101 / 196 = 0
    16'b01100101_11000101 : OUT <= 0;  //101 / 197 = 0
    16'b01100101_11000110 : OUT <= 0;  //101 / 198 = 0
    16'b01100101_11000111 : OUT <= 0;  //101 / 199 = 0
    16'b01100101_11001000 : OUT <= 0;  //101 / 200 = 0
    16'b01100101_11001001 : OUT <= 0;  //101 / 201 = 0
    16'b01100101_11001010 : OUT <= 0;  //101 / 202 = 0
    16'b01100101_11001011 : OUT <= 0;  //101 / 203 = 0
    16'b01100101_11001100 : OUT <= 0;  //101 / 204 = 0
    16'b01100101_11001101 : OUT <= 0;  //101 / 205 = 0
    16'b01100101_11001110 : OUT <= 0;  //101 / 206 = 0
    16'b01100101_11001111 : OUT <= 0;  //101 / 207 = 0
    16'b01100101_11010000 : OUT <= 0;  //101 / 208 = 0
    16'b01100101_11010001 : OUT <= 0;  //101 / 209 = 0
    16'b01100101_11010010 : OUT <= 0;  //101 / 210 = 0
    16'b01100101_11010011 : OUT <= 0;  //101 / 211 = 0
    16'b01100101_11010100 : OUT <= 0;  //101 / 212 = 0
    16'b01100101_11010101 : OUT <= 0;  //101 / 213 = 0
    16'b01100101_11010110 : OUT <= 0;  //101 / 214 = 0
    16'b01100101_11010111 : OUT <= 0;  //101 / 215 = 0
    16'b01100101_11011000 : OUT <= 0;  //101 / 216 = 0
    16'b01100101_11011001 : OUT <= 0;  //101 / 217 = 0
    16'b01100101_11011010 : OUT <= 0;  //101 / 218 = 0
    16'b01100101_11011011 : OUT <= 0;  //101 / 219 = 0
    16'b01100101_11011100 : OUT <= 0;  //101 / 220 = 0
    16'b01100101_11011101 : OUT <= 0;  //101 / 221 = 0
    16'b01100101_11011110 : OUT <= 0;  //101 / 222 = 0
    16'b01100101_11011111 : OUT <= 0;  //101 / 223 = 0
    16'b01100101_11100000 : OUT <= 0;  //101 / 224 = 0
    16'b01100101_11100001 : OUT <= 0;  //101 / 225 = 0
    16'b01100101_11100010 : OUT <= 0;  //101 / 226 = 0
    16'b01100101_11100011 : OUT <= 0;  //101 / 227 = 0
    16'b01100101_11100100 : OUT <= 0;  //101 / 228 = 0
    16'b01100101_11100101 : OUT <= 0;  //101 / 229 = 0
    16'b01100101_11100110 : OUT <= 0;  //101 / 230 = 0
    16'b01100101_11100111 : OUT <= 0;  //101 / 231 = 0
    16'b01100101_11101000 : OUT <= 0;  //101 / 232 = 0
    16'b01100101_11101001 : OUT <= 0;  //101 / 233 = 0
    16'b01100101_11101010 : OUT <= 0;  //101 / 234 = 0
    16'b01100101_11101011 : OUT <= 0;  //101 / 235 = 0
    16'b01100101_11101100 : OUT <= 0;  //101 / 236 = 0
    16'b01100101_11101101 : OUT <= 0;  //101 / 237 = 0
    16'b01100101_11101110 : OUT <= 0;  //101 / 238 = 0
    16'b01100101_11101111 : OUT <= 0;  //101 / 239 = 0
    16'b01100101_11110000 : OUT <= 0;  //101 / 240 = 0
    16'b01100101_11110001 : OUT <= 0;  //101 / 241 = 0
    16'b01100101_11110010 : OUT <= 0;  //101 / 242 = 0
    16'b01100101_11110011 : OUT <= 0;  //101 / 243 = 0
    16'b01100101_11110100 : OUT <= 0;  //101 / 244 = 0
    16'b01100101_11110101 : OUT <= 0;  //101 / 245 = 0
    16'b01100101_11110110 : OUT <= 0;  //101 / 246 = 0
    16'b01100101_11110111 : OUT <= 0;  //101 / 247 = 0
    16'b01100101_11111000 : OUT <= 0;  //101 / 248 = 0
    16'b01100101_11111001 : OUT <= 0;  //101 / 249 = 0
    16'b01100101_11111010 : OUT <= 0;  //101 / 250 = 0
    16'b01100101_11111011 : OUT <= 0;  //101 / 251 = 0
    16'b01100101_11111100 : OUT <= 0;  //101 / 252 = 0
    16'b01100101_11111101 : OUT <= 0;  //101 / 253 = 0
    16'b01100101_11111110 : OUT <= 0;  //101 / 254 = 0
    16'b01100101_11111111 : OUT <= 0;  //101 / 255 = 0
    16'b01100110_00000000 : OUT <= 0;  //102 / 0 = 0
    16'b01100110_00000001 : OUT <= 102;  //102 / 1 = 102
    16'b01100110_00000010 : OUT <= 51;  //102 / 2 = 51
    16'b01100110_00000011 : OUT <= 34;  //102 / 3 = 34
    16'b01100110_00000100 : OUT <= 25;  //102 / 4 = 25
    16'b01100110_00000101 : OUT <= 20;  //102 / 5 = 20
    16'b01100110_00000110 : OUT <= 17;  //102 / 6 = 17
    16'b01100110_00000111 : OUT <= 14;  //102 / 7 = 14
    16'b01100110_00001000 : OUT <= 12;  //102 / 8 = 12
    16'b01100110_00001001 : OUT <= 11;  //102 / 9 = 11
    16'b01100110_00001010 : OUT <= 10;  //102 / 10 = 10
    16'b01100110_00001011 : OUT <= 9;  //102 / 11 = 9
    16'b01100110_00001100 : OUT <= 8;  //102 / 12 = 8
    16'b01100110_00001101 : OUT <= 7;  //102 / 13 = 7
    16'b01100110_00001110 : OUT <= 7;  //102 / 14 = 7
    16'b01100110_00001111 : OUT <= 6;  //102 / 15 = 6
    16'b01100110_00010000 : OUT <= 6;  //102 / 16 = 6
    16'b01100110_00010001 : OUT <= 6;  //102 / 17 = 6
    16'b01100110_00010010 : OUT <= 5;  //102 / 18 = 5
    16'b01100110_00010011 : OUT <= 5;  //102 / 19 = 5
    16'b01100110_00010100 : OUT <= 5;  //102 / 20 = 5
    16'b01100110_00010101 : OUT <= 4;  //102 / 21 = 4
    16'b01100110_00010110 : OUT <= 4;  //102 / 22 = 4
    16'b01100110_00010111 : OUT <= 4;  //102 / 23 = 4
    16'b01100110_00011000 : OUT <= 4;  //102 / 24 = 4
    16'b01100110_00011001 : OUT <= 4;  //102 / 25 = 4
    16'b01100110_00011010 : OUT <= 3;  //102 / 26 = 3
    16'b01100110_00011011 : OUT <= 3;  //102 / 27 = 3
    16'b01100110_00011100 : OUT <= 3;  //102 / 28 = 3
    16'b01100110_00011101 : OUT <= 3;  //102 / 29 = 3
    16'b01100110_00011110 : OUT <= 3;  //102 / 30 = 3
    16'b01100110_00011111 : OUT <= 3;  //102 / 31 = 3
    16'b01100110_00100000 : OUT <= 3;  //102 / 32 = 3
    16'b01100110_00100001 : OUT <= 3;  //102 / 33 = 3
    16'b01100110_00100010 : OUT <= 3;  //102 / 34 = 3
    16'b01100110_00100011 : OUT <= 2;  //102 / 35 = 2
    16'b01100110_00100100 : OUT <= 2;  //102 / 36 = 2
    16'b01100110_00100101 : OUT <= 2;  //102 / 37 = 2
    16'b01100110_00100110 : OUT <= 2;  //102 / 38 = 2
    16'b01100110_00100111 : OUT <= 2;  //102 / 39 = 2
    16'b01100110_00101000 : OUT <= 2;  //102 / 40 = 2
    16'b01100110_00101001 : OUT <= 2;  //102 / 41 = 2
    16'b01100110_00101010 : OUT <= 2;  //102 / 42 = 2
    16'b01100110_00101011 : OUT <= 2;  //102 / 43 = 2
    16'b01100110_00101100 : OUT <= 2;  //102 / 44 = 2
    16'b01100110_00101101 : OUT <= 2;  //102 / 45 = 2
    16'b01100110_00101110 : OUT <= 2;  //102 / 46 = 2
    16'b01100110_00101111 : OUT <= 2;  //102 / 47 = 2
    16'b01100110_00110000 : OUT <= 2;  //102 / 48 = 2
    16'b01100110_00110001 : OUT <= 2;  //102 / 49 = 2
    16'b01100110_00110010 : OUT <= 2;  //102 / 50 = 2
    16'b01100110_00110011 : OUT <= 2;  //102 / 51 = 2
    16'b01100110_00110100 : OUT <= 1;  //102 / 52 = 1
    16'b01100110_00110101 : OUT <= 1;  //102 / 53 = 1
    16'b01100110_00110110 : OUT <= 1;  //102 / 54 = 1
    16'b01100110_00110111 : OUT <= 1;  //102 / 55 = 1
    16'b01100110_00111000 : OUT <= 1;  //102 / 56 = 1
    16'b01100110_00111001 : OUT <= 1;  //102 / 57 = 1
    16'b01100110_00111010 : OUT <= 1;  //102 / 58 = 1
    16'b01100110_00111011 : OUT <= 1;  //102 / 59 = 1
    16'b01100110_00111100 : OUT <= 1;  //102 / 60 = 1
    16'b01100110_00111101 : OUT <= 1;  //102 / 61 = 1
    16'b01100110_00111110 : OUT <= 1;  //102 / 62 = 1
    16'b01100110_00111111 : OUT <= 1;  //102 / 63 = 1
    16'b01100110_01000000 : OUT <= 1;  //102 / 64 = 1
    16'b01100110_01000001 : OUT <= 1;  //102 / 65 = 1
    16'b01100110_01000010 : OUT <= 1;  //102 / 66 = 1
    16'b01100110_01000011 : OUT <= 1;  //102 / 67 = 1
    16'b01100110_01000100 : OUT <= 1;  //102 / 68 = 1
    16'b01100110_01000101 : OUT <= 1;  //102 / 69 = 1
    16'b01100110_01000110 : OUT <= 1;  //102 / 70 = 1
    16'b01100110_01000111 : OUT <= 1;  //102 / 71 = 1
    16'b01100110_01001000 : OUT <= 1;  //102 / 72 = 1
    16'b01100110_01001001 : OUT <= 1;  //102 / 73 = 1
    16'b01100110_01001010 : OUT <= 1;  //102 / 74 = 1
    16'b01100110_01001011 : OUT <= 1;  //102 / 75 = 1
    16'b01100110_01001100 : OUT <= 1;  //102 / 76 = 1
    16'b01100110_01001101 : OUT <= 1;  //102 / 77 = 1
    16'b01100110_01001110 : OUT <= 1;  //102 / 78 = 1
    16'b01100110_01001111 : OUT <= 1;  //102 / 79 = 1
    16'b01100110_01010000 : OUT <= 1;  //102 / 80 = 1
    16'b01100110_01010001 : OUT <= 1;  //102 / 81 = 1
    16'b01100110_01010010 : OUT <= 1;  //102 / 82 = 1
    16'b01100110_01010011 : OUT <= 1;  //102 / 83 = 1
    16'b01100110_01010100 : OUT <= 1;  //102 / 84 = 1
    16'b01100110_01010101 : OUT <= 1;  //102 / 85 = 1
    16'b01100110_01010110 : OUT <= 1;  //102 / 86 = 1
    16'b01100110_01010111 : OUT <= 1;  //102 / 87 = 1
    16'b01100110_01011000 : OUT <= 1;  //102 / 88 = 1
    16'b01100110_01011001 : OUT <= 1;  //102 / 89 = 1
    16'b01100110_01011010 : OUT <= 1;  //102 / 90 = 1
    16'b01100110_01011011 : OUT <= 1;  //102 / 91 = 1
    16'b01100110_01011100 : OUT <= 1;  //102 / 92 = 1
    16'b01100110_01011101 : OUT <= 1;  //102 / 93 = 1
    16'b01100110_01011110 : OUT <= 1;  //102 / 94 = 1
    16'b01100110_01011111 : OUT <= 1;  //102 / 95 = 1
    16'b01100110_01100000 : OUT <= 1;  //102 / 96 = 1
    16'b01100110_01100001 : OUT <= 1;  //102 / 97 = 1
    16'b01100110_01100010 : OUT <= 1;  //102 / 98 = 1
    16'b01100110_01100011 : OUT <= 1;  //102 / 99 = 1
    16'b01100110_01100100 : OUT <= 1;  //102 / 100 = 1
    16'b01100110_01100101 : OUT <= 1;  //102 / 101 = 1
    16'b01100110_01100110 : OUT <= 1;  //102 / 102 = 1
    16'b01100110_01100111 : OUT <= 0;  //102 / 103 = 0
    16'b01100110_01101000 : OUT <= 0;  //102 / 104 = 0
    16'b01100110_01101001 : OUT <= 0;  //102 / 105 = 0
    16'b01100110_01101010 : OUT <= 0;  //102 / 106 = 0
    16'b01100110_01101011 : OUT <= 0;  //102 / 107 = 0
    16'b01100110_01101100 : OUT <= 0;  //102 / 108 = 0
    16'b01100110_01101101 : OUT <= 0;  //102 / 109 = 0
    16'b01100110_01101110 : OUT <= 0;  //102 / 110 = 0
    16'b01100110_01101111 : OUT <= 0;  //102 / 111 = 0
    16'b01100110_01110000 : OUT <= 0;  //102 / 112 = 0
    16'b01100110_01110001 : OUT <= 0;  //102 / 113 = 0
    16'b01100110_01110010 : OUT <= 0;  //102 / 114 = 0
    16'b01100110_01110011 : OUT <= 0;  //102 / 115 = 0
    16'b01100110_01110100 : OUT <= 0;  //102 / 116 = 0
    16'b01100110_01110101 : OUT <= 0;  //102 / 117 = 0
    16'b01100110_01110110 : OUT <= 0;  //102 / 118 = 0
    16'b01100110_01110111 : OUT <= 0;  //102 / 119 = 0
    16'b01100110_01111000 : OUT <= 0;  //102 / 120 = 0
    16'b01100110_01111001 : OUT <= 0;  //102 / 121 = 0
    16'b01100110_01111010 : OUT <= 0;  //102 / 122 = 0
    16'b01100110_01111011 : OUT <= 0;  //102 / 123 = 0
    16'b01100110_01111100 : OUT <= 0;  //102 / 124 = 0
    16'b01100110_01111101 : OUT <= 0;  //102 / 125 = 0
    16'b01100110_01111110 : OUT <= 0;  //102 / 126 = 0
    16'b01100110_01111111 : OUT <= 0;  //102 / 127 = 0
    16'b01100110_10000000 : OUT <= 0;  //102 / 128 = 0
    16'b01100110_10000001 : OUT <= 0;  //102 / 129 = 0
    16'b01100110_10000010 : OUT <= 0;  //102 / 130 = 0
    16'b01100110_10000011 : OUT <= 0;  //102 / 131 = 0
    16'b01100110_10000100 : OUT <= 0;  //102 / 132 = 0
    16'b01100110_10000101 : OUT <= 0;  //102 / 133 = 0
    16'b01100110_10000110 : OUT <= 0;  //102 / 134 = 0
    16'b01100110_10000111 : OUT <= 0;  //102 / 135 = 0
    16'b01100110_10001000 : OUT <= 0;  //102 / 136 = 0
    16'b01100110_10001001 : OUT <= 0;  //102 / 137 = 0
    16'b01100110_10001010 : OUT <= 0;  //102 / 138 = 0
    16'b01100110_10001011 : OUT <= 0;  //102 / 139 = 0
    16'b01100110_10001100 : OUT <= 0;  //102 / 140 = 0
    16'b01100110_10001101 : OUT <= 0;  //102 / 141 = 0
    16'b01100110_10001110 : OUT <= 0;  //102 / 142 = 0
    16'b01100110_10001111 : OUT <= 0;  //102 / 143 = 0
    16'b01100110_10010000 : OUT <= 0;  //102 / 144 = 0
    16'b01100110_10010001 : OUT <= 0;  //102 / 145 = 0
    16'b01100110_10010010 : OUT <= 0;  //102 / 146 = 0
    16'b01100110_10010011 : OUT <= 0;  //102 / 147 = 0
    16'b01100110_10010100 : OUT <= 0;  //102 / 148 = 0
    16'b01100110_10010101 : OUT <= 0;  //102 / 149 = 0
    16'b01100110_10010110 : OUT <= 0;  //102 / 150 = 0
    16'b01100110_10010111 : OUT <= 0;  //102 / 151 = 0
    16'b01100110_10011000 : OUT <= 0;  //102 / 152 = 0
    16'b01100110_10011001 : OUT <= 0;  //102 / 153 = 0
    16'b01100110_10011010 : OUT <= 0;  //102 / 154 = 0
    16'b01100110_10011011 : OUT <= 0;  //102 / 155 = 0
    16'b01100110_10011100 : OUT <= 0;  //102 / 156 = 0
    16'b01100110_10011101 : OUT <= 0;  //102 / 157 = 0
    16'b01100110_10011110 : OUT <= 0;  //102 / 158 = 0
    16'b01100110_10011111 : OUT <= 0;  //102 / 159 = 0
    16'b01100110_10100000 : OUT <= 0;  //102 / 160 = 0
    16'b01100110_10100001 : OUT <= 0;  //102 / 161 = 0
    16'b01100110_10100010 : OUT <= 0;  //102 / 162 = 0
    16'b01100110_10100011 : OUT <= 0;  //102 / 163 = 0
    16'b01100110_10100100 : OUT <= 0;  //102 / 164 = 0
    16'b01100110_10100101 : OUT <= 0;  //102 / 165 = 0
    16'b01100110_10100110 : OUT <= 0;  //102 / 166 = 0
    16'b01100110_10100111 : OUT <= 0;  //102 / 167 = 0
    16'b01100110_10101000 : OUT <= 0;  //102 / 168 = 0
    16'b01100110_10101001 : OUT <= 0;  //102 / 169 = 0
    16'b01100110_10101010 : OUT <= 0;  //102 / 170 = 0
    16'b01100110_10101011 : OUT <= 0;  //102 / 171 = 0
    16'b01100110_10101100 : OUT <= 0;  //102 / 172 = 0
    16'b01100110_10101101 : OUT <= 0;  //102 / 173 = 0
    16'b01100110_10101110 : OUT <= 0;  //102 / 174 = 0
    16'b01100110_10101111 : OUT <= 0;  //102 / 175 = 0
    16'b01100110_10110000 : OUT <= 0;  //102 / 176 = 0
    16'b01100110_10110001 : OUT <= 0;  //102 / 177 = 0
    16'b01100110_10110010 : OUT <= 0;  //102 / 178 = 0
    16'b01100110_10110011 : OUT <= 0;  //102 / 179 = 0
    16'b01100110_10110100 : OUT <= 0;  //102 / 180 = 0
    16'b01100110_10110101 : OUT <= 0;  //102 / 181 = 0
    16'b01100110_10110110 : OUT <= 0;  //102 / 182 = 0
    16'b01100110_10110111 : OUT <= 0;  //102 / 183 = 0
    16'b01100110_10111000 : OUT <= 0;  //102 / 184 = 0
    16'b01100110_10111001 : OUT <= 0;  //102 / 185 = 0
    16'b01100110_10111010 : OUT <= 0;  //102 / 186 = 0
    16'b01100110_10111011 : OUT <= 0;  //102 / 187 = 0
    16'b01100110_10111100 : OUT <= 0;  //102 / 188 = 0
    16'b01100110_10111101 : OUT <= 0;  //102 / 189 = 0
    16'b01100110_10111110 : OUT <= 0;  //102 / 190 = 0
    16'b01100110_10111111 : OUT <= 0;  //102 / 191 = 0
    16'b01100110_11000000 : OUT <= 0;  //102 / 192 = 0
    16'b01100110_11000001 : OUT <= 0;  //102 / 193 = 0
    16'b01100110_11000010 : OUT <= 0;  //102 / 194 = 0
    16'b01100110_11000011 : OUT <= 0;  //102 / 195 = 0
    16'b01100110_11000100 : OUT <= 0;  //102 / 196 = 0
    16'b01100110_11000101 : OUT <= 0;  //102 / 197 = 0
    16'b01100110_11000110 : OUT <= 0;  //102 / 198 = 0
    16'b01100110_11000111 : OUT <= 0;  //102 / 199 = 0
    16'b01100110_11001000 : OUT <= 0;  //102 / 200 = 0
    16'b01100110_11001001 : OUT <= 0;  //102 / 201 = 0
    16'b01100110_11001010 : OUT <= 0;  //102 / 202 = 0
    16'b01100110_11001011 : OUT <= 0;  //102 / 203 = 0
    16'b01100110_11001100 : OUT <= 0;  //102 / 204 = 0
    16'b01100110_11001101 : OUT <= 0;  //102 / 205 = 0
    16'b01100110_11001110 : OUT <= 0;  //102 / 206 = 0
    16'b01100110_11001111 : OUT <= 0;  //102 / 207 = 0
    16'b01100110_11010000 : OUT <= 0;  //102 / 208 = 0
    16'b01100110_11010001 : OUT <= 0;  //102 / 209 = 0
    16'b01100110_11010010 : OUT <= 0;  //102 / 210 = 0
    16'b01100110_11010011 : OUT <= 0;  //102 / 211 = 0
    16'b01100110_11010100 : OUT <= 0;  //102 / 212 = 0
    16'b01100110_11010101 : OUT <= 0;  //102 / 213 = 0
    16'b01100110_11010110 : OUT <= 0;  //102 / 214 = 0
    16'b01100110_11010111 : OUT <= 0;  //102 / 215 = 0
    16'b01100110_11011000 : OUT <= 0;  //102 / 216 = 0
    16'b01100110_11011001 : OUT <= 0;  //102 / 217 = 0
    16'b01100110_11011010 : OUT <= 0;  //102 / 218 = 0
    16'b01100110_11011011 : OUT <= 0;  //102 / 219 = 0
    16'b01100110_11011100 : OUT <= 0;  //102 / 220 = 0
    16'b01100110_11011101 : OUT <= 0;  //102 / 221 = 0
    16'b01100110_11011110 : OUT <= 0;  //102 / 222 = 0
    16'b01100110_11011111 : OUT <= 0;  //102 / 223 = 0
    16'b01100110_11100000 : OUT <= 0;  //102 / 224 = 0
    16'b01100110_11100001 : OUT <= 0;  //102 / 225 = 0
    16'b01100110_11100010 : OUT <= 0;  //102 / 226 = 0
    16'b01100110_11100011 : OUT <= 0;  //102 / 227 = 0
    16'b01100110_11100100 : OUT <= 0;  //102 / 228 = 0
    16'b01100110_11100101 : OUT <= 0;  //102 / 229 = 0
    16'b01100110_11100110 : OUT <= 0;  //102 / 230 = 0
    16'b01100110_11100111 : OUT <= 0;  //102 / 231 = 0
    16'b01100110_11101000 : OUT <= 0;  //102 / 232 = 0
    16'b01100110_11101001 : OUT <= 0;  //102 / 233 = 0
    16'b01100110_11101010 : OUT <= 0;  //102 / 234 = 0
    16'b01100110_11101011 : OUT <= 0;  //102 / 235 = 0
    16'b01100110_11101100 : OUT <= 0;  //102 / 236 = 0
    16'b01100110_11101101 : OUT <= 0;  //102 / 237 = 0
    16'b01100110_11101110 : OUT <= 0;  //102 / 238 = 0
    16'b01100110_11101111 : OUT <= 0;  //102 / 239 = 0
    16'b01100110_11110000 : OUT <= 0;  //102 / 240 = 0
    16'b01100110_11110001 : OUT <= 0;  //102 / 241 = 0
    16'b01100110_11110010 : OUT <= 0;  //102 / 242 = 0
    16'b01100110_11110011 : OUT <= 0;  //102 / 243 = 0
    16'b01100110_11110100 : OUT <= 0;  //102 / 244 = 0
    16'b01100110_11110101 : OUT <= 0;  //102 / 245 = 0
    16'b01100110_11110110 : OUT <= 0;  //102 / 246 = 0
    16'b01100110_11110111 : OUT <= 0;  //102 / 247 = 0
    16'b01100110_11111000 : OUT <= 0;  //102 / 248 = 0
    16'b01100110_11111001 : OUT <= 0;  //102 / 249 = 0
    16'b01100110_11111010 : OUT <= 0;  //102 / 250 = 0
    16'b01100110_11111011 : OUT <= 0;  //102 / 251 = 0
    16'b01100110_11111100 : OUT <= 0;  //102 / 252 = 0
    16'b01100110_11111101 : OUT <= 0;  //102 / 253 = 0
    16'b01100110_11111110 : OUT <= 0;  //102 / 254 = 0
    16'b01100110_11111111 : OUT <= 0;  //102 / 255 = 0
    16'b01100111_00000000 : OUT <= 0;  //103 / 0 = 0
    16'b01100111_00000001 : OUT <= 103;  //103 / 1 = 103
    16'b01100111_00000010 : OUT <= 51;  //103 / 2 = 51
    16'b01100111_00000011 : OUT <= 34;  //103 / 3 = 34
    16'b01100111_00000100 : OUT <= 25;  //103 / 4 = 25
    16'b01100111_00000101 : OUT <= 20;  //103 / 5 = 20
    16'b01100111_00000110 : OUT <= 17;  //103 / 6 = 17
    16'b01100111_00000111 : OUT <= 14;  //103 / 7 = 14
    16'b01100111_00001000 : OUT <= 12;  //103 / 8 = 12
    16'b01100111_00001001 : OUT <= 11;  //103 / 9 = 11
    16'b01100111_00001010 : OUT <= 10;  //103 / 10 = 10
    16'b01100111_00001011 : OUT <= 9;  //103 / 11 = 9
    16'b01100111_00001100 : OUT <= 8;  //103 / 12 = 8
    16'b01100111_00001101 : OUT <= 7;  //103 / 13 = 7
    16'b01100111_00001110 : OUT <= 7;  //103 / 14 = 7
    16'b01100111_00001111 : OUT <= 6;  //103 / 15 = 6
    16'b01100111_00010000 : OUT <= 6;  //103 / 16 = 6
    16'b01100111_00010001 : OUT <= 6;  //103 / 17 = 6
    16'b01100111_00010010 : OUT <= 5;  //103 / 18 = 5
    16'b01100111_00010011 : OUT <= 5;  //103 / 19 = 5
    16'b01100111_00010100 : OUT <= 5;  //103 / 20 = 5
    16'b01100111_00010101 : OUT <= 4;  //103 / 21 = 4
    16'b01100111_00010110 : OUT <= 4;  //103 / 22 = 4
    16'b01100111_00010111 : OUT <= 4;  //103 / 23 = 4
    16'b01100111_00011000 : OUT <= 4;  //103 / 24 = 4
    16'b01100111_00011001 : OUT <= 4;  //103 / 25 = 4
    16'b01100111_00011010 : OUT <= 3;  //103 / 26 = 3
    16'b01100111_00011011 : OUT <= 3;  //103 / 27 = 3
    16'b01100111_00011100 : OUT <= 3;  //103 / 28 = 3
    16'b01100111_00011101 : OUT <= 3;  //103 / 29 = 3
    16'b01100111_00011110 : OUT <= 3;  //103 / 30 = 3
    16'b01100111_00011111 : OUT <= 3;  //103 / 31 = 3
    16'b01100111_00100000 : OUT <= 3;  //103 / 32 = 3
    16'b01100111_00100001 : OUT <= 3;  //103 / 33 = 3
    16'b01100111_00100010 : OUT <= 3;  //103 / 34 = 3
    16'b01100111_00100011 : OUT <= 2;  //103 / 35 = 2
    16'b01100111_00100100 : OUT <= 2;  //103 / 36 = 2
    16'b01100111_00100101 : OUT <= 2;  //103 / 37 = 2
    16'b01100111_00100110 : OUT <= 2;  //103 / 38 = 2
    16'b01100111_00100111 : OUT <= 2;  //103 / 39 = 2
    16'b01100111_00101000 : OUT <= 2;  //103 / 40 = 2
    16'b01100111_00101001 : OUT <= 2;  //103 / 41 = 2
    16'b01100111_00101010 : OUT <= 2;  //103 / 42 = 2
    16'b01100111_00101011 : OUT <= 2;  //103 / 43 = 2
    16'b01100111_00101100 : OUT <= 2;  //103 / 44 = 2
    16'b01100111_00101101 : OUT <= 2;  //103 / 45 = 2
    16'b01100111_00101110 : OUT <= 2;  //103 / 46 = 2
    16'b01100111_00101111 : OUT <= 2;  //103 / 47 = 2
    16'b01100111_00110000 : OUT <= 2;  //103 / 48 = 2
    16'b01100111_00110001 : OUT <= 2;  //103 / 49 = 2
    16'b01100111_00110010 : OUT <= 2;  //103 / 50 = 2
    16'b01100111_00110011 : OUT <= 2;  //103 / 51 = 2
    16'b01100111_00110100 : OUT <= 1;  //103 / 52 = 1
    16'b01100111_00110101 : OUT <= 1;  //103 / 53 = 1
    16'b01100111_00110110 : OUT <= 1;  //103 / 54 = 1
    16'b01100111_00110111 : OUT <= 1;  //103 / 55 = 1
    16'b01100111_00111000 : OUT <= 1;  //103 / 56 = 1
    16'b01100111_00111001 : OUT <= 1;  //103 / 57 = 1
    16'b01100111_00111010 : OUT <= 1;  //103 / 58 = 1
    16'b01100111_00111011 : OUT <= 1;  //103 / 59 = 1
    16'b01100111_00111100 : OUT <= 1;  //103 / 60 = 1
    16'b01100111_00111101 : OUT <= 1;  //103 / 61 = 1
    16'b01100111_00111110 : OUT <= 1;  //103 / 62 = 1
    16'b01100111_00111111 : OUT <= 1;  //103 / 63 = 1
    16'b01100111_01000000 : OUT <= 1;  //103 / 64 = 1
    16'b01100111_01000001 : OUT <= 1;  //103 / 65 = 1
    16'b01100111_01000010 : OUT <= 1;  //103 / 66 = 1
    16'b01100111_01000011 : OUT <= 1;  //103 / 67 = 1
    16'b01100111_01000100 : OUT <= 1;  //103 / 68 = 1
    16'b01100111_01000101 : OUT <= 1;  //103 / 69 = 1
    16'b01100111_01000110 : OUT <= 1;  //103 / 70 = 1
    16'b01100111_01000111 : OUT <= 1;  //103 / 71 = 1
    16'b01100111_01001000 : OUT <= 1;  //103 / 72 = 1
    16'b01100111_01001001 : OUT <= 1;  //103 / 73 = 1
    16'b01100111_01001010 : OUT <= 1;  //103 / 74 = 1
    16'b01100111_01001011 : OUT <= 1;  //103 / 75 = 1
    16'b01100111_01001100 : OUT <= 1;  //103 / 76 = 1
    16'b01100111_01001101 : OUT <= 1;  //103 / 77 = 1
    16'b01100111_01001110 : OUT <= 1;  //103 / 78 = 1
    16'b01100111_01001111 : OUT <= 1;  //103 / 79 = 1
    16'b01100111_01010000 : OUT <= 1;  //103 / 80 = 1
    16'b01100111_01010001 : OUT <= 1;  //103 / 81 = 1
    16'b01100111_01010010 : OUT <= 1;  //103 / 82 = 1
    16'b01100111_01010011 : OUT <= 1;  //103 / 83 = 1
    16'b01100111_01010100 : OUT <= 1;  //103 / 84 = 1
    16'b01100111_01010101 : OUT <= 1;  //103 / 85 = 1
    16'b01100111_01010110 : OUT <= 1;  //103 / 86 = 1
    16'b01100111_01010111 : OUT <= 1;  //103 / 87 = 1
    16'b01100111_01011000 : OUT <= 1;  //103 / 88 = 1
    16'b01100111_01011001 : OUT <= 1;  //103 / 89 = 1
    16'b01100111_01011010 : OUT <= 1;  //103 / 90 = 1
    16'b01100111_01011011 : OUT <= 1;  //103 / 91 = 1
    16'b01100111_01011100 : OUT <= 1;  //103 / 92 = 1
    16'b01100111_01011101 : OUT <= 1;  //103 / 93 = 1
    16'b01100111_01011110 : OUT <= 1;  //103 / 94 = 1
    16'b01100111_01011111 : OUT <= 1;  //103 / 95 = 1
    16'b01100111_01100000 : OUT <= 1;  //103 / 96 = 1
    16'b01100111_01100001 : OUT <= 1;  //103 / 97 = 1
    16'b01100111_01100010 : OUT <= 1;  //103 / 98 = 1
    16'b01100111_01100011 : OUT <= 1;  //103 / 99 = 1
    16'b01100111_01100100 : OUT <= 1;  //103 / 100 = 1
    16'b01100111_01100101 : OUT <= 1;  //103 / 101 = 1
    16'b01100111_01100110 : OUT <= 1;  //103 / 102 = 1
    16'b01100111_01100111 : OUT <= 1;  //103 / 103 = 1
    16'b01100111_01101000 : OUT <= 0;  //103 / 104 = 0
    16'b01100111_01101001 : OUT <= 0;  //103 / 105 = 0
    16'b01100111_01101010 : OUT <= 0;  //103 / 106 = 0
    16'b01100111_01101011 : OUT <= 0;  //103 / 107 = 0
    16'b01100111_01101100 : OUT <= 0;  //103 / 108 = 0
    16'b01100111_01101101 : OUT <= 0;  //103 / 109 = 0
    16'b01100111_01101110 : OUT <= 0;  //103 / 110 = 0
    16'b01100111_01101111 : OUT <= 0;  //103 / 111 = 0
    16'b01100111_01110000 : OUT <= 0;  //103 / 112 = 0
    16'b01100111_01110001 : OUT <= 0;  //103 / 113 = 0
    16'b01100111_01110010 : OUT <= 0;  //103 / 114 = 0
    16'b01100111_01110011 : OUT <= 0;  //103 / 115 = 0
    16'b01100111_01110100 : OUT <= 0;  //103 / 116 = 0
    16'b01100111_01110101 : OUT <= 0;  //103 / 117 = 0
    16'b01100111_01110110 : OUT <= 0;  //103 / 118 = 0
    16'b01100111_01110111 : OUT <= 0;  //103 / 119 = 0
    16'b01100111_01111000 : OUT <= 0;  //103 / 120 = 0
    16'b01100111_01111001 : OUT <= 0;  //103 / 121 = 0
    16'b01100111_01111010 : OUT <= 0;  //103 / 122 = 0
    16'b01100111_01111011 : OUT <= 0;  //103 / 123 = 0
    16'b01100111_01111100 : OUT <= 0;  //103 / 124 = 0
    16'b01100111_01111101 : OUT <= 0;  //103 / 125 = 0
    16'b01100111_01111110 : OUT <= 0;  //103 / 126 = 0
    16'b01100111_01111111 : OUT <= 0;  //103 / 127 = 0
    16'b01100111_10000000 : OUT <= 0;  //103 / 128 = 0
    16'b01100111_10000001 : OUT <= 0;  //103 / 129 = 0
    16'b01100111_10000010 : OUT <= 0;  //103 / 130 = 0
    16'b01100111_10000011 : OUT <= 0;  //103 / 131 = 0
    16'b01100111_10000100 : OUT <= 0;  //103 / 132 = 0
    16'b01100111_10000101 : OUT <= 0;  //103 / 133 = 0
    16'b01100111_10000110 : OUT <= 0;  //103 / 134 = 0
    16'b01100111_10000111 : OUT <= 0;  //103 / 135 = 0
    16'b01100111_10001000 : OUT <= 0;  //103 / 136 = 0
    16'b01100111_10001001 : OUT <= 0;  //103 / 137 = 0
    16'b01100111_10001010 : OUT <= 0;  //103 / 138 = 0
    16'b01100111_10001011 : OUT <= 0;  //103 / 139 = 0
    16'b01100111_10001100 : OUT <= 0;  //103 / 140 = 0
    16'b01100111_10001101 : OUT <= 0;  //103 / 141 = 0
    16'b01100111_10001110 : OUT <= 0;  //103 / 142 = 0
    16'b01100111_10001111 : OUT <= 0;  //103 / 143 = 0
    16'b01100111_10010000 : OUT <= 0;  //103 / 144 = 0
    16'b01100111_10010001 : OUT <= 0;  //103 / 145 = 0
    16'b01100111_10010010 : OUT <= 0;  //103 / 146 = 0
    16'b01100111_10010011 : OUT <= 0;  //103 / 147 = 0
    16'b01100111_10010100 : OUT <= 0;  //103 / 148 = 0
    16'b01100111_10010101 : OUT <= 0;  //103 / 149 = 0
    16'b01100111_10010110 : OUT <= 0;  //103 / 150 = 0
    16'b01100111_10010111 : OUT <= 0;  //103 / 151 = 0
    16'b01100111_10011000 : OUT <= 0;  //103 / 152 = 0
    16'b01100111_10011001 : OUT <= 0;  //103 / 153 = 0
    16'b01100111_10011010 : OUT <= 0;  //103 / 154 = 0
    16'b01100111_10011011 : OUT <= 0;  //103 / 155 = 0
    16'b01100111_10011100 : OUT <= 0;  //103 / 156 = 0
    16'b01100111_10011101 : OUT <= 0;  //103 / 157 = 0
    16'b01100111_10011110 : OUT <= 0;  //103 / 158 = 0
    16'b01100111_10011111 : OUT <= 0;  //103 / 159 = 0
    16'b01100111_10100000 : OUT <= 0;  //103 / 160 = 0
    16'b01100111_10100001 : OUT <= 0;  //103 / 161 = 0
    16'b01100111_10100010 : OUT <= 0;  //103 / 162 = 0
    16'b01100111_10100011 : OUT <= 0;  //103 / 163 = 0
    16'b01100111_10100100 : OUT <= 0;  //103 / 164 = 0
    16'b01100111_10100101 : OUT <= 0;  //103 / 165 = 0
    16'b01100111_10100110 : OUT <= 0;  //103 / 166 = 0
    16'b01100111_10100111 : OUT <= 0;  //103 / 167 = 0
    16'b01100111_10101000 : OUT <= 0;  //103 / 168 = 0
    16'b01100111_10101001 : OUT <= 0;  //103 / 169 = 0
    16'b01100111_10101010 : OUT <= 0;  //103 / 170 = 0
    16'b01100111_10101011 : OUT <= 0;  //103 / 171 = 0
    16'b01100111_10101100 : OUT <= 0;  //103 / 172 = 0
    16'b01100111_10101101 : OUT <= 0;  //103 / 173 = 0
    16'b01100111_10101110 : OUT <= 0;  //103 / 174 = 0
    16'b01100111_10101111 : OUT <= 0;  //103 / 175 = 0
    16'b01100111_10110000 : OUT <= 0;  //103 / 176 = 0
    16'b01100111_10110001 : OUT <= 0;  //103 / 177 = 0
    16'b01100111_10110010 : OUT <= 0;  //103 / 178 = 0
    16'b01100111_10110011 : OUT <= 0;  //103 / 179 = 0
    16'b01100111_10110100 : OUT <= 0;  //103 / 180 = 0
    16'b01100111_10110101 : OUT <= 0;  //103 / 181 = 0
    16'b01100111_10110110 : OUT <= 0;  //103 / 182 = 0
    16'b01100111_10110111 : OUT <= 0;  //103 / 183 = 0
    16'b01100111_10111000 : OUT <= 0;  //103 / 184 = 0
    16'b01100111_10111001 : OUT <= 0;  //103 / 185 = 0
    16'b01100111_10111010 : OUT <= 0;  //103 / 186 = 0
    16'b01100111_10111011 : OUT <= 0;  //103 / 187 = 0
    16'b01100111_10111100 : OUT <= 0;  //103 / 188 = 0
    16'b01100111_10111101 : OUT <= 0;  //103 / 189 = 0
    16'b01100111_10111110 : OUT <= 0;  //103 / 190 = 0
    16'b01100111_10111111 : OUT <= 0;  //103 / 191 = 0
    16'b01100111_11000000 : OUT <= 0;  //103 / 192 = 0
    16'b01100111_11000001 : OUT <= 0;  //103 / 193 = 0
    16'b01100111_11000010 : OUT <= 0;  //103 / 194 = 0
    16'b01100111_11000011 : OUT <= 0;  //103 / 195 = 0
    16'b01100111_11000100 : OUT <= 0;  //103 / 196 = 0
    16'b01100111_11000101 : OUT <= 0;  //103 / 197 = 0
    16'b01100111_11000110 : OUT <= 0;  //103 / 198 = 0
    16'b01100111_11000111 : OUT <= 0;  //103 / 199 = 0
    16'b01100111_11001000 : OUT <= 0;  //103 / 200 = 0
    16'b01100111_11001001 : OUT <= 0;  //103 / 201 = 0
    16'b01100111_11001010 : OUT <= 0;  //103 / 202 = 0
    16'b01100111_11001011 : OUT <= 0;  //103 / 203 = 0
    16'b01100111_11001100 : OUT <= 0;  //103 / 204 = 0
    16'b01100111_11001101 : OUT <= 0;  //103 / 205 = 0
    16'b01100111_11001110 : OUT <= 0;  //103 / 206 = 0
    16'b01100111_11001111 : OUT <= 0;  //103 / 207 = 0
    16'b01100111_11010000 : OUT <= 0;  //103 / 208 = 0
    16'b01100111_11010001 : OUT <= 0;  //103 / 209 = 0
    16'b01100111_11010010 : OUT <= 0;  //103 / 210 = 0
    16'b01100111_11010011 : OUT <= 0;  //103 / 211 = 0
    16'b01100111_11010100 : OUT <= 0;  //103 / 212 = 0
    16'b01100111_11010101 : OUT <= 0;  //103 / 213 = 0
    16'b01100111_11010110 : OUT <= 0;  //103 / 214 = 0
    16'b01100111_11010111 : OUT <= 0;  //103 / 215 = 0
    16'b01100111_11011000 : OUT <= 0;  //103 / 216 = 0
    16'b01100111_11011001 : OUT <= 0;  //103 / 217 = 0
    16'b01100111_11011010 : OUT <= 0;  //103 / 218 = 0
    16'b01100111_11011011 : OUT <= 0;  //103 / 219 = 0
    16'b01100111_11011100 : OUT <= 0;  //103 / 220 = 0
    16'b01100111_11011101 : OUT <= 0;  //103 / 221 = 0
    16'b01100111_11011110 : OUT <= 0;  //103 / 222 = 0
    16'b01100111_11011111 : OUT <= 0;  //103 / 223 = 0
    16'b01100111_11100000 : OUT <= 0;  //103 / 224 = 0
    16'b01100111_11100001 : OUT <= 0;  //103 / 225 = 0
    16'b01100111_11100010 : OUT <= 0;  //103 / 226 = 0
    16'b01100111_11100011 : OUT <= 0;  //103 / 227 = 0
    16'b01100111_11100100 : OUT <= 0;  //103 / 228 = 0
    16'b01100111_11100101 : OUT <= 0;  //103 / 229 = 0
    16'b01100111_11100110 : OUT <= 0;  //103 / 230 = 0
    16'b01100111_11100111 : OUT <= 0;  //103 / 231 = 0
    16'b01100111_11101000 : OUT <= 0;  //103 / 232 = 0
    16'b01100111_11101001 : OUT <= 0;  //103 / 233 = 0
    16'b01100111_11101010 : OUT <= 0;  //103 / 234 = 0
    16'b01100111_11101011 : OUT <= 0;  //103 / 235 = 0
    16'b01100111_11101100 : OUT <= 0;  //103 / 236 = 0
    16'b01100111_11101101 : OUT <= 0;  //103 / 237 = 0
    16'b01100111_11101110 : OUT <= 0;  //103 / 238 = 0
    16'b01100111_11101111 : OUT <= 0;  //103 / 239 = 0
    16'b01100111_11110000 : OUT <= 0;  //103 / 240 = 0
    16'b01100111_11110001 : OUT <= 0;  //103 / 241 = 0
    16'b01100111_11110010 : OUT <= 0;  //103 / 242 = 0
    16'b01100111_11110011 : OUT <= 0;  //103 / 243 = 0
    16'b01100111_11110100 : OUT <= 0;  //103 / 244 = 0
    16'b01100111_11110101 : OUT <= 0;  //103 / 245 = 0
    16'b01100111_11110110 : OUT <= 0;  //103 / 246 = 0
    16'b01100111_11110111 : OUT <= 0;  //103 / 247 = 0
    16'b01100111_11111000 : OUT <= 0;  //103 / 248 = 0
    16'b01100111_11111001 : OUT <= 0;  //103 / 249 = 0
    16'b01100111_11111010 : OUT <= 0;  //103 / 250 = 0
    16'b01100111_11111011 : OUT <= 0;  //103 / 251 = 0
    16'b01100111_11111100 : OUT <= 0;  //103 / 252 = 0
    16'b01100111_11111101 : OUT <= 0;  //103 / 253 = 0
    16'b01100111_11111110 : OUT <= 0;  //103 / 254 = 0
    16'b01100111_11111111 : OUT <= 0;  //103 / 255 = 0
    16'b01101000_00000000 : OUT <= 0;  //104 / 0 = 0
    16'b01101000_00000001 : OUT <= 104;  //104 / 1 = 104
    16'b01101000_00000010 : OUT <= 52;  //104 / 2 = 52
    16'b01101000_00000011 : OUT <= 34;  //104 / 3 = 34
    16'b01101000_00000100 : OUT <= 26;  //104 / 4 = 26
    16'b01101000_00000101 : OUT <= 20;  //104 / 5 = 20
    16'b01101000_00000110 : OUT <= 17;  //104 / 6 = 17
    16'b01101000_00000111 : OUT <= 14;  //104 / 7 = 14
    16'b01101000_00001000 : OUT <= 13;  //104 / 8 = 13
    16'b01101000_00001001 : OUT <= 11;  //104 / 9 = 11
    16'b01101000_00001010 : OUT <= 10;  //104 / 10 = 10
    16'b01101000_00001011 : OUT <= 9;  //104 / 11 = 9
    16'b01101000_00001100 : OUT <= 8;  //104 / 12 = 8
    16'b01101000_00001101 : OUT <= 8;  //104 / 13 = 8
    16'b01101000_00001110 : OUT <= 7;  //104 / 14 = 7
    16'b01101000_00001111 : OUT <= 6;  //104 / 15 = 6
    16'b01101000_00010000 : OUT <= 6;  //104 / 16 = 6
    16'b01101000_00010001 : OUT <= 6;  //104 / 17 = 6
    16'b01101000_00010010 : OUT <= 5;  //104 / 18 = 5
    16'b01101000_00010011 : OUT <= 5;  //104 / 19 = 5
    16'b01101000_00010100 : OUT <= 5;  //104 / 20 = 5
    16'b01101000_00010101 : OUT <= 4;  //104 / 21 = 4
    16'b01101000_00010110 : OUT <= 4;  //104 / 22 = 4
    16'b01101000_00010111 : OUT <= 4;  //104 / 23 = 4
    16'b01101000_00011000 : OUT <= 4;  //104 / 24 = 4
    16'b01101000_00011001 : OUT <= 4;  //104 / 25 = 4
    16'b01101000_00011010 : OUT <= 4;  //104 / 26 = 4
    16'b01101000_00011011 : OUT <= 3;  //104 / 27 = 3
    16'b01101000_00011100 : OUT <= 3;  //104 / 28 = 3
    16'b01101000_00011101 : OUT <= 3;  //104 / 29 = 3
    16'b01101000_00011110 : OUT <= 3;  //104 / 30 = 3
    16'b01101000_00011111 : OUT <= 3;  //104 / 31 = 3
    16'b01101000_00100000 : OUT <= 3;  //104 / 32 = 3
    16'b01101000_00100001 : OUT <= 3;  //104 / 33 = 3
    16'b01101000_00100010 : OUT <= 3;  //104 / 34 = 3
    16'b01101000_00100011 : OUT <= 2;  //104 / 35 = 2
    16'b01101000_00100100 : OUT <= 2;  //104 / 36 = 2
    16'b01101000_00100101 : OUT <= 2;  //104 / 37 = 2
    16'b01101000_00100110 : OUT <= 2;  //104 / 38 = 2
    16'b01101000_00100111 : OUT <= 2;  //104 / 39 = 2
    16'b01101000_00101000 : OUT <= 2;  //104 / 40 = 2
    16'b01101000_00101001 : OUT <= 2;  //104 / 41 = 2
    16'b01101000_00101010 : OUT <= 2;  //104 / 42 = 2
    16'b01101000_00101011 : OUT <= 2;  //104 / 43 = 2
    16'b01101000_00101100 : OUT <= 2;  //104 / 44 = 2
    16'b01101000_00101101 : OUT <= 2;  //104 / 45 = 2
    16'b01101000_00101110 : OUT <= 2;  //104 / 46 = 2
    16'b01101000_00101111 : OUT <= 2;  //104 / 47 = 2
    16'b01101000_00110000 : OUT <= 2;  //104 / 48 = 2
    16'b01101000_00110001 : OUT <= 2;  //104 / 49 = 2
    16'b01101000_00110010 : OUT <= 2;  //104 / 50 = 2
    16'b01101000_00110011 : OUT <= 2;  //104 / 51 = 2
    16'b01101000_00110100 : OUT <= 2;  //104 / 52 = 2
    16'b01101000_00110101 : OUT <= 1;  //104 / 53 = 1
    16'b01101000_00110110 : OUT <= 1;  //104 / 54 = 1
    16'b01101000_00110111 : OUT <= 1;  //104 / 55 = 1
    16'b01101000_00111000 : OUT <= 1;  //104 / 56 = 1
    16'b01101000_00111001 : OUT <= 1;  //104 / 57 = 1
    16'b01101000_00111010 : OUT <= 1;  //104 / 58 = 1
    16'b01101000_00111011 : OUT <= 1;  //104 / 59 = 1
    16'b01101000_00111100 : OUT <= 1;  //104 / 60 = 1
    16'b01101000_00111101 : OUT <= 1;  //104 / 61 = 1
    16'b01101000_00111110 : OUT <= 1;  //104 / 62 = 1
    16'b01101000_00111111 : OUT <= 1;  //104 / 63 = 1
    16'b01101000_01000000 : OUT <= 1;  //104 / 64 = 1
    16'b01101000_01000001 : OUT <= 1;  //104 / 65 = 1
    16'b01101000_01000010 : OUT <= 1;  //104 / 66 = 1
    16'b01101000_01000011 : OUT <= 1;  //104 / 67 = 1
    16'b01101000_01000100 : OUT <= 1;  //104 / 68 = 1
    16'b01101000_01000101 : OUT <= 1;  //104 / 69 = 1
    16'b01101000_01000110 : OUT <= 1;  //104 / 70 = 1
    16'b01101000_01000111 : OUT <= 1;  //104 / 71 = 1
    16'b01101000_01001000 : OUT <= 1;  //104 / 72 = 1
    16'b01101000_01001001 : OUT <= 1;  //104 / 73 = 1
    16'b01101000_01001010 : OUT <= 1;  //104 / 74 = 1
    16'b01101000_01001011 : OUT <= 1;  //104 / 75 = 1
    16'b01101000_01001100 : OUT <= 1;  //104 / 76 = 1
    16'b01101000_01001101 : OUT <= 1;  //104 / 77 = 1
    16'b01101000_01001110 : OUT <= 1;  //104 / 78 = 1
    16'b01101000_01001111 : OUT <= 1;  //104 / 79 = 1
    16'b01101000_01010000 : OUT <= 1;  //104 / 80 = 1
    16'b01101000_01010001 : OUT <= 1;  //104 / 81 = 1
    16'b01101000_01010010 : OUT <= 1;  //104 / 82 = 1
    16'b01101000_01010011 : OUT <= 1;  //104 / 83 = 1
    16'b01101000_01010100 : OUT <= 1;  //104 / 84 = 1
    16'b01101000_01010101 : OUT <= 1;  //104 / 85 = 1
    16'b01101000_01010110 : OUT <= 1;  //104 / 86 = 1
    16'b01101000_01010111 : OUT <= 1;  //104 / 87 = 1
    16'b01101000_01011000 : OUT <= 1;  //104 / 88 = 1
    16'b01101000_01011001 : OUT <= 1;  //104 / 89 = 1
    16'b01101000_01011010 : OUT <= 1;  //104 / 90 = 1
    16'b01101000_01011011 : OUT <= 1;  //104 / 91 = 1
    16'b01101000_01011100 : OUT <= 1;  //104 / 92 = 1
    16'b01101000_01011101 : OUT <= 1;  //104 / 93 = 1
    16'b01101000_01011110 : OUT <= 1;  //104 / 94 = 1
    16'b01101000_01011111 : OUT <= 1;  //104 / 95 = 1
    16'b01101000_01100000 : OUT <= 1;  //104 / 96 = 1
    16'b01101000_01100001 : OUT <= 1;  //104 / 97 = 1
    16'b01101000_01100010 : OUT <= 1;  //104 / 98 = 1
    16'b01101000_01100011 : OUT <= 1;  //104 / 99 = 1
    16'b01101000_01100100 : OUT <= 1;  //104 / 100 = 1
    16'b01101000_01100101 : OUT <= 1;  //104 / 101 = 1
    16'b01101000_01100110 : OUT <= 1;  //104 / 102 = 1
    16'b01101000_01100111 : OUT <= 1;  //104 / 103 = 1
    16'b01101000_01101000 : OUT <= 1;  //104 / 104 = 1
    16'b01101000_01101001 : OUT <= 0;  //104 / 105 = 0
    16'b01101000_01101010 : OUT <= 0;  //104 / 106 = 0
    16'b01101000_01101011 : OUT <= 0;  //104 / 107 = 0
    16'b01101000_01101100 : OUT <= 0;  //104 / 108 = 0
    16'b01101000_01101101 : OUT <= 0;  //104 / 109 = 0
    16'b01101000_01101110 : OUT <= 0;  //104 / 110 = 0
    16'b01101000_01101111 : OUT <= 0;  //104 / 111 = 0
    16'b01101000_01110000 : OUT <= 0;  //104 / 112 = 0
    16'b01101000_01110001 : OUT <= 0;  //104 / 113 = 0
    16'b01101000_01110010 : OUT <= 0;  //104 / 114 = 0
    16'b01101000_01110011 : OUT <= 0;  //104 / 115 = 0
    16'b01101000_01110100 : OUT <= 0;  //104 / 116 = 0
    16'b01101000_01110101 : OUT <= 0;  //104 / 117 = 0
    16'b01101000_01110110 : OUT <= 0;  //104 / 118 = 0
    16'b01101000_01110111 : OUT <= 0;  //104 / 119 = 0
    16'b01101000_01111000 : OUT <= 0;  //104 / 120 = 0
    16'b01101000_01111001 : OUT <= 0;  //104 / 121 = 0
    16'b01101000_01111010 : OUT <= 0;  //104 / 122 = 0
    16'b01101000_01111011 : OUT <= 0;  //104 / 123 = 0
    16'b01101000_01111100 : OUT <= 0;  //104 / 124 = 0
    16'b01101000_01111101 : OUT <= 0;  //104 / 125 = 0
    16'b01101000_01111110 : OUT <= 0;  //104 / 126 = 0
    16'b01101000_01111111 : OUT <= 0;  //104 / 127 = 0
    16'b01101000_10000000 : OUT <= 0;  //104 / 128 = 0
    16'b01101000_10000001 : OUT <= 0;  //104 / 129 = 0
    16'b01101000_10000010 : OUT <= 0;  //104 / 130 = 0
    16'b01101000_10000011 : OUT <= 0;  //104 / 131 = 0
    16'b01101000_10000100 : OUT <= 0;  //104 / 132 = 0
    16'b01101000_10000101 : OUT <= 0;  //104 / 133 = 0
    16'b01101000_10000110 : OUT <= 0;  //104 / 134 = 0
    16'b01101000_10000111 : OUT <= 0;  //104 / 135 = 0
    16'b01101000_10001000 : OUT <= 0;  //104 / 136 = 0
    16'b01101000_10001001 : OUT <= 0;  //104 / 137 = 0
    16'b01101000_10001010 : OUT <= 0;  //104 / 138 = 0
    16'b01101000_10001011 : OUT <= 0;  //104 / 139 = 0
    16'b01101000_10001100 : OUT <= 0;  //104 / 140 = 0
    16'b01101000_10001101 : OUT <= 0;  //104 / 141 = 0
    16'b01101000_10001110 : OUT <= 0;  //104 / 142 = 0
    16'b01101000_10001111 : OUT <= 0;  //104 / 143 = 0
    16'b01101000_10010000 : OUT <= 0;  //104 / 144 = 0
    16'b01101000_10010001 : OUT <= 0;  //104 / 145 = 0
    16'b01101000_10010010 : OUT <= 0;  //104 / 146 = 0
    16'b01101000_10010011 : OUT <= 0;  //104 / 147 = 0
    16'b01101000_10010100 : OUT <= 0;  //104 / 148 = 0
    16'b01101000_10010101 : OUT <= 0;  //104 / 149 = 0
    16'b01101000_10010110 : OUT <= 0;  //104 / 150 = 0
    16'b01101000_10010111 : OUT <= 0;  //104 / 151 = 0
    16'b01101000_10011000 : OUT <= 0;  //104 / 152 = 0
    16'b01101000_10011001 : OUT <= 0;  //104 / 153 = 0
    16'b01101000_10011010 : OUT <= 0;  //104 / 154 = 0
    16'b01101000_10011011 : OUT <= 0;  //104 / 155 = 0
    16'b01101000_10011100 : OUT <= 0;  //104 / 156 = 0
    16'b01101000_10011101 : OUT <= 0;  //104 / 157 = 0
    16'b01101000_10011110 : OUT <= 0;  //104 / 158 = 0
    16'b01101000_10011111 : OUT <= 0;  //104 / 159 = 0
    16'b01101000_10100000 : OUT <= 0;  //104 / 160 = 0
    16'b01101000_10100001 : OUT <= 0;  //104 / 161 = 0
    16'b01101000_10100010 : OUT <= 0;  //104 / 162 = 0
    16'b01101000_10100011 : OUT <= 0;  //104 / 163 = 0
    16'b01101000_10100100 : OUT <= 0;  //104 / 164 = 0
    16'b01101000_10100101 : OUT <= 0;  //104 / 165 = 0
    16'b01101000_10100110 : OUT <= 0;  //104 / 166 = 0
    16'b01101000_10100111 : OUT <= 0;  //104 / 167 = 0
    16'b01101000_10101000 : OUT <= 0;  //104 / 168 = 0
    16'b01101000_10101001 : OUT <= 0;  //104 / 169 = 0
    16'b01101000_10101010 : OUT <= 0;  //104 / 170 = 0
    16'b01101000_10101011 : OUT <= 0;  //104 / 171 = 0
    16'b01101000_10101100 : OUT <= 0;  //104 / 172 = 0
    16'b01101000_10101101 : OUT <= 0;  //104 / 173 = 0
    16'b01101000_10101110 : OUT <= 0;  //104 / 174 = 0
    16'b01101000_10101111 : OUT <= 0;  //104 / 175 = 0
    16'b01101000_10110000 : OUT <= 0;  //104 / 176 = 0
    16'b01101000_10110001 : OUT <= 0;  //104 / 177 = 0
    16'b01101000_10110010 : OUT <= 0;  //104 / 178 = 0
    16'b01101000_10110011 : OUT <= 0;  //104 / 179 = 0
    16'b01101000_10110100 : OUT <= 0;  //104 / 180 = 0
    16'b01101000_10110101 : OUT <= 0;  //104 / 181 = 0
    16'b01101000_10110110 : OUT <= 0;  //104 / 182 = 0
    16'b01101000_10110111 : OUT <= 0;  //104 / 183 = 0
    16'b01101000_10111000 : OUT <= 0;  //104 / 184 = 0
    16'b01101000_10111001 : OUT <= 0;  //104 / 185 = 0
    16'b01101000_10111010 : OUT <= 0;  //104 / 186 = 0
    16'b01101000_10111011 : OUT <= 0;  //104 / 187 = 0
    16'b01101000_10111100 : OUT <= 0;  //104 / 188 = 0
    16'b01101000_10111101 : OUT <= 0;  //104 / 189 = 0
    16'b01101000_10111110 : OUT <= 0;  //104 / 190 = 0
    16'b01101000_10111111 : OUT <= 0;  //104 / 191 = 0
    16'b01101000_11000000 : OUT <= 0;  //104 / 192 = 0
    16'b01101000_11000001 : OUT <= 0;  //104 / 193 = 0
    16'b01101000_11000010 : OUT <= 0;  //104 / 194 = 0
    16'b01101000_11000011 : OUT <= 0;  //104 / 195 = 0
    16'b01101000_11000100 : OUT <= 0;  //104 / 196 = 0
    16'b01101000_11000101 : OUT <= 0;  //104 / 197 = 0
    16'b01101000_11000110 : OUT <= 0;  //104 / 198 = 0
    16'b01101000_11000111 : OUT <= 0;  //104 / 199 = 0
    16'b01101000_11001000 : OUT <= 0;  //104 / 200 = 0
    16'b01101000_11001001 : OUT <= 0;  //104 / 201 = 0
    16'b01101000_11001010 : OUT <= 0;  //104 / 202 = 0
    16'b01101000_11001011 : OUT <= 0;  //104 / 203 = 0
    16'b01101000_11001100 : OUT <= 0;  //104 / 204 = 0
    16'b01101000_11001101 : OUT <= 0;  //104 / 205 = 0
    16'b01101000_11001110 : OUT <= 0;  //104 / 206 = 0
    16'b01101000_11001111 : OUT <= 0;  //104 / 207 = 0
    16'b01101000_11010000 : OUT <= 0;  //104 / 208 = 0
    16'b01101000_11010001 : OUT <= 0;  //104 / 209 = 0
    16'b01101000_11010010 : OUT <= 0;  //104 / 210 = 0
    16'b01101000_11010011 : OUT <= 0;  //104 / 211 = 0
    16'b01101000_11010100 : OUT <= 0;  //104 / 212 = 0
    16'b01101000_11010101 : OUT <= 0;  //104 / 213 = 0
    16'b01101000_11010110 : OUT <= 0;  //104 / 214 = 0
    16'b01101000_11010111 : OUT <= 0;  //104 / 215 = 0
    16'b01101000_11011000 : OUT <= 0;  //104 / 216 = 0
    16'b01101000_11011001 : OUT <= 0;  //104 / 217 = 0
    16'b01101000_11011010 : OUT <= 0;  //104 / 218 = 0
    16'b01101000_11011011 : OUT <= 0;  //104 / 219 = 0
    16'b01101000_11011100 : OUT <= 0;  //104 / 220 = 0
    16'b01101000_11011101 : OUT <= 0;  //104 / 221 = 0
    16'b01101000_11011110 : OUT <= 0;  //104 / 222 = 0
    16'b01101000_11011111 : OUT <= 0;  //104 / 223 = 0
    16'b01101000_11100000 : OUT <= 0;  //104 / 224 = 0
    16'b01101000_11100001 : OUT <= 0;  //104 / 225 = 0
    16'b01101000_11100010 : OUT <= 0;  //104 / 226 = 0
    16'b01101000_11100011 : OUT <= 0;  //104 / 227 = 0
    16'b01101000_11100100 : OUT <= 0;  //104 / 228 = 0
    16'b01101000_11100101 : OUT <= 0;  //104 / 229 = 0
    16'b01101000_11100110 : OUT <= 0;  //104 / 230 = 0
    16'b01101000_11100111 : OUT <= 0;  //104 / 231 = 0
    16'b01101000_11101000 : OUT <= 0;  //104 / 232 = 0
    16'b01101000_11101001 : OUT <= 0;  //104 / 233 = 0
    16'b01101000_11101010 : OUT <= 0;  //104 / 234 = 0
    16'b01101000_11101011 : OUT <= 0;  //104 / 235 = 0
    16'b01101000_11101100 : OUT <= 0;  //104 / 236 = 0
    16'b01101000_11101101 : OUT <= 0;  //104 / 237 = 0
    16'b01101000_11101110 : OUT <= 0;  //104 / 238 = 0
    16'b01101000_11101111 : OUT <= 0;  //104 / 239 = 0
    16'b01101000_11110000 : OUT <= 0;  //104 / 240 = 0
    16'b01101000_11110001 : OUT <= 0;  //104 / 241 = 0
    16'b01101000_11110010 : OUT <= 0;  //104 / 242 = 0
    16'b01101000_11110011 : OUT <= 0;  //104 / 243 = 0
    16'b01101000_11110100 : OUT <= 0;  //104 / 244 = 0
    16'b01101000_11110101 : OUT <= 0;  //104 / 245 = 0
    16'b01101000_11110110 : OUT <= 0;  //104 / 246 = 0
    16'b01101000_11110111 : OUT <= 0;  //104 / 247 = 0
    16'b01101000_11111000 : OUT <= 0;  //104 / 248 = 0
    16'b01101000_11111001 : OUT <= 0;  //104 / 249 = 0
    16'b01101000_11111010 : OUT <= 0;  //104 / 250 = 0
    16'b01101000_11111011 : OUT <= 0;  //104 / 251 = 0
    16'b01101000_11111100 : OUT <= 0;  //104 / 252 = 0
    16'b01101000_11111101 : OUT <= 0;  //104 / 253 = 0
    16'b01101000_11111110 : OUT <= 0;  //104 / 254 = 0
    16'b01101000_11111111 : OUT <= 0;  //104 / 255 = 0
    16'b01101001_00000000 : OUT <= 0;  //105 / 0 = 0
    16'b01101001_00000001 : OUT <= 105;  //105 / 1 = 105
    16'b01101001_00000010 : OUT <= 52;  //105 / 2 = 52
    16'b01101001_00000011 : OUT <= 35;  //105 / 3 = 35
    16'b01101001_00000100 : OUT <= 26;  //105 / 4 = 26
    16'b01101001_00000101 : OUT <= 21;  //105 / 5 = 21
    16'b01101001_00000110 : OUT <= 17;  //105 / 6 = 17
    16'b01101001_00000111 : OUT <= 15;  //105 / 7 = 15
    16'b01101001_00001000 : OUT <= 13;  //105 / 8 = 13
    16'b01101001_00001001 : OUT <= 11;  //105 / 9 = 11
    16'b01101001_00001010 : OUT <= 10;  //105 / 10 = 10
    16'b01101001_00001011 : OUT <= 9;  //105 / 11 = 9
    16'b01101001_00001100 : OUT <= 8;  //105 / 12 = 8
    16'b01101001_00001101 : OUT <= 8;  //105 / 13 = 8
    16'b01101001_00001110 : OUT <= 7;  //105 / 14 = 7
    16'b01101001_00001111 : OUT <= 7;  //105 / 15 = 7
    16'b01101001_00010000 : OUT <= 6;  //105 / 16 = 6
    16'b01101001_00010001 : OUT <= 6;  //105 / 17 = 6
    16'b01101001_00010010 : OUT <= 5;  //105 / 18 = 5
    16'b01101001_00010011 : OUT <= 5;  //105 / 19 = 5
    16'b01101001_00010100 : OUT <= 5;  //105 / 20 = 5
    16'b01101001_00010101 : OUT <= 5;  //105 / 21 = 5
    16'b01101001_00010110 : OUT <= 4;  //105 / 22 = 4
    16'b01101001_00010111 : OUT <= 4;  //105 / 23 = 4
    16'b01101001_00011000 : OUT <= 4;  //105 / 24 = 4
    16'b01101001_00011001 : OUT <= 4;  //105 / 25 = 4
    16'b01101001_00011010 : OUT <= 4;  //105 / 26 = 4
    16'b01101001_00011011 : OUT <= 3;  //105 / 27 = 3
    16'b01101001_00011100 : OUT <= 3;  //105 / 28 = 3
    16'b01101001_00011101 : OUT <= 3;  //105 / 29 = 3
    16'b01101001_00011110 : OUT <= 3;  //105 / 30 = 3
    16'b01101001_00011111 : OUT <= 3;  //105 / 31 = 3
    16'b01101001_00100000 : OUT <= 3;  //105 / 32 = 3
    16'b01101001_00100001 : OUT <= 3;  //105 / 33 = 3
    16'b01101001_00100010 : OUT <= 3;  //105 / 34 = 3
    16'b01101001_00100011 : OUT <= 3;  //105 / 35 = 3
    16'b01101001_00100100 : OUT <= 2;  //105 / 36 = 2
    16'b01101001_00100101 : OUT <= 2;  //105 / 37 = 2
    16'b01101001_00100110 : OUT <= 2;  //105 / 38 = 2
    16'b01101001_00100111 : OUT <= 2;  //105 / 39 = 2
    16'b01101001_00101000 : OUT <= 2;  //105 / 40 = 2
    16'b01101001_00101001 : OUT <= 2;  //105 / 41 = 2
    16'b01101001_00101010 : OUT <= 2;  //105 / 42 = 2
    16'b01101001_00101011 : OUT <= 2;  //105 / 43 = 2
    16'b01101001_00101100 : OUT <= 2;  //105 / 44 = 2
    16'b01101001_00101101 : OUT <= 2;  //105 / 45 = 2
    16'b01101001_00101110 : OUT <= 2;  //105 / 46 = 2
    16'b01101001_00101111 : OUT <= 2;  //105 / 47 = 2
    16'b01101001_00110000 : OUT <= 2;  //105 / 48 = 2
    16'b01101001_00110001 : OUT <= 2;  //105 / 49 = 2
    16'b01101001_00110010 : OUT <= 2;  //105 / 50 = 2
    16'b01101001_00110011 : OUT <= 2;  //105 / 51 = 2
    16'b01101001_00110100 : OUT <= 2;  //105 / 52 = 2
    16'b01101001_00110101 : OUT <= 1;  //105 / 53 = 1
    16'b01101001_00110110 : OUT <= 1;  //105 / 54 = 1
    16'b01101001_00110111 : OUT <= 1;  //105 / 55 = 1
    16'b01101001_00111000 : OUT <= 1;  //105 / 56 = 1
    16'b01101001_00111001 : OUT <= 1;  //105 / 57 = 1
    16'b01101001_00111010 : OUT <= 1;  //105 / 58 = 1
    16'b01101001_00111011 : OUT <= 1;  //105 / 59 = 1
    16'b01101001_00111100 : OUT <= 1;  //105 / 60 = 1
    16'b01101001_00111101 : OUT <= 1;  //105 / 61 = 1
    16'b01101001_00111110 : OUT <= 1;  //105 / 62 = 1
    16'b01101001_00111111 : OUT <= 1;  //105 / 63 = 1
    16'b01101001_01000000 : OUT <= 1;  //105 / 64 = 1
    16'b01101001_01000001 : OUT <= 1;  //105 / 65 = 1
    16'b01101001_01000010 : OUT <= 1;  //105 / 66 = 1
    16'b01101001_01000011 : OUT <= 1;  //105 / 67 = 1
    16'b01101001_01000100 : OUT <= 1;  //105 / 68 = 1
    16'b01101001_01000101 : OUT <= 1;  //105 / 69 = 1
    16'b01101001_01000110 : OUT <= 1;  //105 / 70 = 1
    16'b01101001_01000111 : OUT <= 1;  //105 / 71 = 1
    16'b01101001_01001000 : OUT <= 1;  //105 / 72 = 1
    16'b01101001_01001001 : OUT <= 1;  //105 / 73 = 1
    16'b01101001_01001010 : OUT <= 1;  //105 / 74 = 1
    16'b01101001_01001011 : OUT <= 1;  //105 / 75 = 1
    16'b01101001_01001100 : OUT <= 1;  //105 / 76 = 1
    16'b01101001_01001101 : OUT <= 1;  //105 / 77 = 1
    16'b01101001_01001110 : OUT <= 1;  //105 / 78 = 1
    16'b01101001_01001111 : OUT <= 1;  //105 / 79 = 1
    16'b01101001_01010000 : OUT <= 1;  //105 / 80 = 1
    16'b01101001_01010001 : OUT <= 1;  //105 / 81 = 1
    16'b01101001_01010010 : OUT <= 1;  //105 / 82 = 1
    16'b01101001_01010011 : OUT <= 1;  //105 / 83 = 1
    16'b01101001_01010100 : OUT <= 1;  //105 / 84 = 1
    16'b01101001_01010101 : OUT <= 1;  //105 / 85 = 1
    16'b01101001_01010110 : OUT <= 1;  //105 / 86 = 1
    16'b01101001_01010111 : OUT <= 1;  //105 / 87 = 1
    16'b01101001_01011000 : OUT <= 1;  //105 / 88 = 1
    16'b01101001_01011001 : OUT <= 1;  //105 / 89 = 1
    16'b01101001_01011010 : OUT <= 1;  //105 / 90 = 1
    16'b01101001_01011011 : OUT <= 1;  //105 / 91 = 1
    16'b01101001_01011100 : OUT <= 1;  //105 / 92 = 1
    16'b01101001_01011101 : OUT <= 1;  //105 / 93 = 1
    16'b01101001_01011110 : OUT <= 1;  //105 / 94 = 1
    16'b01101001_01011111 : OUT <= 1;  //105 / 95 = 1
    16'b01101001_01100000 : OUT <= 1;  //105 / 96 = 1
    16'b01101001_01100001 : OUT <= 1;  //105 / 97 = 1
    16'b01101001_01100010 : OUT <= 1;  //105 / 98 = 1
    16'b01101001_01100011 : OUT <= 1;  //105 / 99 = 1
    16'b01101001_01100100 : OUT <= 1;  //105 / 100 = 1
    16'b01101001_01100101 : OUT <= 1;  //105 / 101 = 1
    16'b01101001_01100110 : OUT <= 1;  //105 / 102 = 1
    16'b01101001_01100111 : OUT <= 1;  //105 / 103 = 1
    16'b01101001_01101000 : OUT <= 1;  //105 / 104 = 1
    16'b01101001_01101001 : OUT <= 1;  //105 / 105 = 1
    16'b01101001_01101010 : OUT <= 0;  //105 / 106 = 0
    16'b01101001_01101011 : OUT <= 0;  //105 / 107 = 0
    16'b01101001_01101100 : OUT <= 0;  //105 / 108 = 0
    16'b01101001_01101101 : OUT <= 0;  //105 / 109 = 0
    16'b01101001_01101110 : OUT <= 0;  //105 / 110 = 0
    16'b01101001_01101111 : OUT <= 0;  //105 / 111 = 0
    16'b01101001_01110000 : OUT <= 0;  //105 / 112 = 0
    16'b01101001_01110001 : OUT <= 0;  //105 / 113 = 0
    16'b01101001_01110010 : OUT <= 0;  //105 / 114 = 0
    16'b01101001_01110011 : OUT <= 0;  //105 / 115 = 0
    16'b01101001_01110100 : OUT <= 0;  //105 / 116 = 0
    16'b01101001_01110101 : OUT <= 0;  //105 / 117 = 0
    16'b01101001_01110110 : OUT <= 0;  //105 / 118 = 0
    16'b01101001_01110111 : OUT <= 0;  //105 / 119 = 0
    16'b01101001_01111000 : OUT <= 0;  //105 / 120 = 0
    16'b01101001_01111001 : OUT <= 0;  //105 / 121 = 0
    16'b01101001_01111010 : OUT <= 0;  //105 / 122 = 0
    16'b01101001_01111011 : OUT <= 0;  //105 / 123 = 0
    16'b01101001_01111100 : OUT <= 0;  //105 / 124 = 0
    16'b01101001_01111101 : OUT <= 0;  //105 / 125 = 0
    16'b01101001_01111110 : OUT <= 0;  //105 / 126 = 0
    16'b01101001_01111111 : OUT <= 0;  //105 / 127 = 0
    16'b01101001_10000000 : OUT <= 0;  //105 / 128 = 0
    16'b01101001_10000001 : OUT <= 0;  //105 / 129 = 0
    16'b01101001_10000010 : OUT <= 0;  //105 / 130 = 0
    16'b01101001_10000011 : OUT <= 0;  //105 / 131 = 0
    16'b01101001_10000100 : OUT <= 0;  //105 / 132 = 0
    16'b01101001_10000101 : OUT <= 0;  //105 / 133 = 0
    16'b01101001_10000110 : OUT <= 0;  //105 / 134 = 0
    16'b01101001_10000111 : OUT <= 0;  //105 / 135 = 0
    16'b01101001_10001000 : OUT <= 0;  //105 / 136 = 0
    16'b01101001_10001001 : OUT <= 0;  //105 / 137 = 0
    16'b01101001_10001010 : OUT <= 0;  //105 / 138 = 0
    16'b01101001_10001011 : OUT <= 0;  //105 / 139 = 0
    16'b01101001_10001100 : OUT <= 0;  //105 / 140 = 0
    16'b01101001_10001101 : OUT <= 0;  //105 / 141 = 0
    16'b01101001_10001110 : OUT <= 0;  //105 / 142 = 0
    16'b01101001_10001111 : OUT <= 0;  //105 / 143 = 0
    16'b01101001_10010000 : OUT <= 0;  //105 / 144 = 0
    16'b01101001_10010001 : OUT <= 0;  //105 / 145 = 0
    16'b01101001_10010010 : OUT <= 0;  //105 / 146 = 0
    16'b01101001_10010011 : OUT <= 0;  //105 / 147 = 0
    16'b01101001_10010100 : OUT <= 0;  //105 / 148 = 0
    16'b01101001_10010101 : OUT <= 0;  //105 / 149 = 0
    16'b01101001_10010110 : OUT <= 0;  //105 / 150 = 0
    16'b01101001_10010111 : OUT <= 0;  //105 / 151 = 0
    16'b01101001_10011000 : OUT <= 0;  //105 / 152 = 0
    16'b01101001_10011001 : OUT <= 0;  //105 / 153 = 0
    16'b01101001_10011010 : OUT <= 0;  //105 / 154 = 0
    16'b01101001_10011011 : OUT <= 0;  //105 / 155 = 0
    16'b01101001_10011100 : OUT <= 0;  //105 / 156 = 0
    16'b01101001_10011101 : OUT <= 0;  //105 / 157 = 0
    16'b01101001_10011110 : OUT <= 0;  //105 / 158 = 0
    16'b01101001_10011111 : OUT <= 0;  //105 / 159 = 0
    16'b01101001_10100000 : OUT <= 0;  //105 / 160 = 0
    16'b01101001_10100001 : OUT <= 0;  //105 / 161 = 0
    16'b01101001_10100010 : OUT <= 0;  //105 / 162 = 0
    16'b01101001_10100011 : OUT <= 0;  //105 / 163 = 0
    16'b01101001_10100100 : OUT <= 0;  //105 / 164 = 0
    16'b01101001_10100101 : OUT <= 0;  //105 / 165 = 0
    16'b01101001_10100110 : OUT <= 0;  //105 / 166 = 0
    16'b01101001_10100111 : OUT <= 0;  //105 / 167 = 0
    16'b01101001_10101000 : OUT <= 0;  //105 / 168 = 0
    16'b01101001_10101001 : OUT <= 0;  //105 / 169 = 0
    16'b01101001_10101010 : OUT <= 0;  //105 / 170 = 0
    16'b01101001_10101011 : OUT <= 0;  //105 / 171 = 0
    16'b01101001_10101100 : OUT <= 0;  //105 / 172 = 0
    16'b01101001_10101101 : OUT <= 0;  //105 / 173 = 0
    16'b01101001_10101110 : OUT <= 0;  //105 / 174 = 0
    16'b01101001_10101111 : OUT <= 0;  //105 / 175 = 0
    16'b01101001_10110000 : OUT <= 0;  //105 / 176 = 0
    16'b01101001_10110001 : OUT <= 0;  //105 / 177 = 0
    16'b01101001_10110010 : OUT <= 0;  //105 / 178 = 0
    16'b01101001_10110011 : OUT <= 0;  //105 / 179 = 0
    16'b01101001_10110100 : OUT <= 0;  //105 / 180 = 0
    16'b01101001_10110101 : OUT <= 0;  //105 / 181 = 0
    16'b01101001_10110110 : OUT <= 0;  //105 / 182 = 0
    16'b01101001_10110111 : OUT <= 0;  //105 / 183 = 0
    16'b01101001_10111000 : OUT <= 0;  //105 / 184 = 0
    16'b01101001_10111001 : OUT <= 0;  //105 / 185 = 0
    16'b01101001_10111010 : OUT <= 0;  //105 / 186 = 0
    16'b01101001_10111011 : OUT <= 0;  //105 / 187 = 0
    16'b01101001_10111100 : OUT <= 0;  //105 / 188 = 0
    16'b01101001_10111101 : OUT <= 0;  //105 / 189 = 0
    16'b01101001_10111110 : OUT <= 0;  //105 / 190 = 0
    16'b01101001_10111111 : OUT <= 0;  //105 / 191 = 0
    16'b01101001_11000000 : OUT <= 0;  //105 / 192 = 0
    16'b01101001_11000001 : OUT <= 0;  //105 / 193 = 0
    16'b01101001_11000010 : OUT <= 0;  //105 / 194 = 0
    16'b01101001_11000011 : OUT <= 0;  //105 / 195 = 0
    16'b01101001_11000100 : OUT <= 0;  //105 / 196 = 0
    16'b01101001_11000101 : OUT <= 0;  //105 / 197 = 0
    16'b01101001_11000110 : OUT <= 0;  //105 / 198 = 0
    16'b01101001_11000111 : OUT <= 0;  //105 / 199 = 0
    16'b01101001_11001000 : OUT <= 0;  //105 / 200 = 0
    16'b01101001_11001001 : OUT <= 0;  //105 / 201 = 0
    16'b01101001_11001010 : OUT <= 0;  //105 / 202 = 0
    16'b01101001_11001011 : OUT <= 0;  //105 / 203 = 0
    16'b01101001_11001100 : OUT <= 0;  //105 / 204 = 0
    16'b01101001_11001101 : OUT <= 0;  //105 / 205 = 0
    16'b01101001_11001110 : OUT <= 0;  //105 / 206 = 0
    16'b01101001_11001111 : OUT <= 0;  //105 / 207 = 0
    16'b01101001_11010000 : OUT <= 0;  //105 / 208 = 0
    16'b01101001_11010001 : OUT <= 0;  //105 / 209 = 0
    16'b01101001_11010010 : OUT <= 0;  //105 / 210 = 0
    16'b01101001_11010011 : OUT <= 0;  //105 / 211 = 0
    16'b01101001_11010100 : OUT <= 0;  //105 / 212 = 0
    16'b01101001_11010101 : OUT <= 0;  //105 / 213 = 0
    16'b01101001_11010110 : OUT <= 0;  //105 / 214 = 0
    16'b01101001_11010111 : OUT <= 0;  //105 / 215 = 0
    16'b01101001_11011000 : OUT <= 0;  //105 / 216 = 0
    16'b01101001_11011001 : OUT <= 0;  //105 / 217 = 0
    16'b01101001_11011010 : OUT <= 0;  //105 / 218 = 0
    16'b01101001_11011011 : OUT <= 0;  //105 / 219 = 0
    16'b01101001_11011100 : OUT <= 0;  //105 / 220 = 0
    16'b01101001_11011101 : OUT <= 0;  //105 / 221 = 0
    16'b01101001_11011110 : OUT <= 0;  //105 / 222 = 0
    16'b01101001_11011111 : OUT <= 0;  //105 / 223 = 0
    16'b01101001_11100000 : OUT <= 0;  //105 / 224 = 0
    16'b01101001_11100001 : OUT <= 0;  //105 / 225 = 0
    16'b01101001_11100010 : OUT <= 0;  //105 / 226 = 0
    16'b01101001_11100011 : OUT <= 0;  //105 / 227 = 0
    16'b01101001_11100100 : OUT <= 0;  //105 / 228 = 0
    16'b01101001_11100101 : OUT <= 0;  //105 / 229 = 0
    16'b01101001_11100110 : OUT <= 0;  //105 / 230 = 0
    16'b01101001_11100111 : OUT <= 0;  //105 / 231 = 0
    16'b01101001_11101000 : OUT <= 0;  //105 / 232 = 0
    16'b01101001_11101001 : OUT <= 0;  //105 / 233 = 0
    16'b01101001_11101010 : OUT <= 0;  //105 / 234 = 0
    16'b01101001_11101011 : OUT <= 0;  //105 / 235 = 0
    16'b01101001_11101100 : OUT <= 0;  //105 / 236 = 0
    16'b01101001_11101101 : OUT <= 0;  //105 / 237 = 0
    16'b01101001_11101110 : OUT <= 0;  //105 / 238 = 0
    16'b01101001_11101111 : OUT <= 0;  //105 / 239 = 0
    16'b01101001_11110000 : OUT <= 0;  //105 / 240 = 0
    16'b01101001_11110001 : OUT <= 0;  //105 / 241 = 0
    16'b01101001_11110010 : OUT <= 0;  //105 / 242 = 0
    16'b01101001_11110011 : OUT <= 0;  //105 / 243 = 0
    16'b01101001_11110100 : OUT <= 0;  //105 / 244 = 0
    16'b01101001_11110101 : OUT <= 0;  //105 / 245 = 0
    16'b01101001_11110110 : OUT <= 0;  //105 / 246 = 0
    16'b01101001_11110111 : OUT <= 0;  //105 / 247 = 0
    16'b01101001_11111000 : OUT <= 0;  //105 / 248 = 0
    16'b01101001_11111001 : OUT <= 0;  //105 / 249 = 0
    16'b01101001_11111010 : OUT <= 0;  //105 / 250 = 0
    16'b01101001_11111011 : OUT <= 0;  //105 / 251 = 0
    16'b01101001_11111100 : OUT <= 0;  //105 / 252 = 0
    16'b01101001_11111101 : OUT <= 0;  //105 / 253 = 0
    16'b01101001_11111110 : OUT <= 0;  //105 / 254 = 0
    16'b01101001_11111111 : OUT <= 0;  //105 / 255 = 0
    16'b01101010_00000000 : OUT <= 0;  //106 / 0 = 0
    16'b01101010_00000001 : OUT <= 106;  //106 / 1 = 106
    16'b01101010_00000010 : OUT <= 53;  //106 / 2 = 53
    16'b01101010_00000011 : OUT <= 35;  //106 / 3 = 35
    16'b01101010_00000100 : OUT <= 26;  //106 / 4 = 26
    16'b01101010_00000101 : OUT <= 21;  //106 / 5 = 21
    16'b01101010_00000110 : OUT <= 17;  //106 / 6 = 17
    16'b01101010_00000111 : OUT <= 15;  //106 / 7 = 15
    16'b01101010_00001000 : OUT <= 13;  //106 / 8 = 13
    16'b01101010_00001001 : OUT <= 11;  //106 / 9 = 11
    16'b01101010_00001010 : OUT <= 10;  //106 / 10 = 10
    16'b01101010_00001011 : OUT <= 9;  //106 / 11 = 9
    16'b01101010_00001100 : OUT <= 8;  //106 / 12 = 8
    16'b01101010_00001101 : OUT <= 8;  //106 / 13 = 8
    16'b01101010_00001110 : OUT <= 7;  //106 / 14 = 7
    16'b01101010_00001111 : OUT <= 7;  //106 / 15 = 7
    16'b01101010_00010000 : OUT <= 6;  //106 / 16 = 6
    16'b01101010_00010001 : OUT <= 6;  //106 / 17 = 6
    16'b01101010_00010010 : OUT <= 5;  //106 / 18 = 5
    16'b01101010_00010011 : OUT <= 5;  //106 / 19 = 5
    16'b01101010_00010100 : OUT <= 5;  //106 / 20 = 5
    16'b01101010_00010101 : OUT <= 5;  //106 / 21 = 5
    16'b01101010_00010110 : OUT <= 4;  //106 / 22 = 4
    16'b01101010_00010111 : OUT <= 4;  //106 / 23 = 4
    16'b01101010_00011000 : OUT <= 4;  //106 / 24 = 4
    16'b01101010_00011001 : OUT <= 4;  //106 / 25 = 4
    16'b01101010_00011010 : OUT <= 4;  //106 / 26 = 4
    16'b01101010_00011011 : OUT <= 3;  //106 / 27 = 3
    16'b01101010_00011100 : OUT <= 3;  //106 / 28 = 3
    16'b01101010_00011101 : OUT <= 3;  //106 / 29 = 3
    16'b01101010_00011110 : OUT <= 3;  //106 / 30 = 3
    16'b01101010_00011111 : OUT <= 3;  //106 / 31 = 3
    16'b01101010_00100000 : OUT <= 3;  //106 / 32 = 3
    16'b01101010_00100001 : OUT <= 3;  //106 / 33 = 3
    16'b01101010_00100010 : OUT <= 3;  //106 / 34 = 3
    16'b01101010_00100011 : OUT <= 3;  //106 / 35 = 3
    16'b01101010_00100100 : OUT <= 2;  //106 / 36 = 2
    16'b01101010_00100101 : OUT <= 2;  //106 / 37 = 2
    16'b01101010_00100110 : OUT <= 2;  //106 / 38 = 2
    16'b01101010_00100111 : OUT <= 2;  //106 / 39 = 2
    16'b01101010_00101000 : OUT <= 2;  //106 / 40 = 2
    16'b01101010_00101001 : OUT <= 2;  //106 / 41 = 2
    16'b01101010_00101010 : OUT <= 2;  //106 / 42 = 2
    16'b01101010_00101011 : OUT <= 2;  //106 / 43 = 2
    16'b01101010_00101100 : OUT <= 2;  //106 / 44 = 2
    16'b01101010_00101101 : OUT <= 2;  //106 / 45 = 2
    16'b01101010_00101110 : OUT <= 2;  //106 / 46 = 2
    16'b01101010_00101111 : OUT <= 2;  //106 / 47 = 2
    16'b01101010_00110000 : OUT <= 2;  //106 / 48 = 2
    16'b01101010_00110001 : OUT <= 2;  //106 / 49 = 2
    16'b01101010_00110010 : OUT <= 2;  //106 / 50 = 2
    16'b01101010_00110011 : OUT <= 2;  //106 / 51 = 2
    16'b01101010_00110100 : OUT <= 2;  //106 / 52 = 2
    16'b01101010_00110101 : OUT <= 2;  //106 / 53 = 2
    16'b01101010_00110110 : OUT <= 1;  //106 / 54 = 1
    16'b01101010_00110111 : OUT <= 1;  //106 / 55 = 1
    16'b01101010_00111000 : OUT <= 1;  //106 / 56 = 1
    16'b01101010_00111001 : OUT <= 1;  //106 / 57 = 1
    16'b01101010_00111010 : OUT <= 1;  //106 / 58 = 1
    16'b01101010_00111011 : OUT <= 1;  //106 / 59 = 1
    16'b01101010_00111100 : OUT <= 1;  //106 / 60 = 1
    16'b01101010_00111101 : OUT <= 1;  //106 / 61 = 1
    16'b01101010_00111110 : OUT <= 1;  //106 / 62 = 1
    16'b01101010_00111111 : OUT <= 1;  //106 / 63 = 1
    16'b01101010_01000000 : OUT <= 1;  //106 / 64 = 1
    16'b01101010_01000001 : OUT <= 1;  //106 / 65 = 1
    16'b01101010_01000010 : OUT <= 1;  //106 / 66 = 1
    16'b01101010_01000011 : OUT <= 1;  //106 / 67 = 1
    16'b01101010_01000100 : OUT <= 1;  //106 / 68 = 1
    16'b01101010_01000101 : OUT <= 1;  //106 / 69 = 1
    16'b01101010_01000110 : OUT <= 1;  //106 / 70 = 1
    16'b01101010_01000111 : OUT <= 1;  //106 / 71 = 1
    16'b01101010_01001000 : OUT <= 1;  //106 / 72 = 1
    16'b01101010_01001001 : OUT <= 1;  //106 / 73 = 1
    16'b01101010_01001010 : OUT <= 1;  //106 / 74 = 1
    16'b01101010_01001011 : OUT <= 1;  //106 / 75 = 1
    16'b01101010_01001100 : OUT <= 1;  //106 / 76 = 1
    16'b01101010_01001101 : OUT <= 1;  //106 / 77 = 1
    16'b01101010_01001110 : OUT <= 1;  //106 / 78 = 1
    16'b01101010_01001111 : OUT <= 1;  //106 / 79 = 1
    16'b01101010_01010000 : OUT <= 1;  //106 / 80 = 1
    16'b01101010_01010001 : OUT <= 1;  //106 / 81 = 1
    16'b01101010_01010010 : OUT <= 1;  //106 / 82 = 1
    16'b01101010_01010011 : OUT <= 1;  //106 / 83 = 1
    16'b01101010_01010100 : OUT <= 1;  //106 / 84 = 1
    16'b01101010_01010101 : OUT <= 1;  //106 / 85 = 1
    16'b01101010_01010110 : OUT <= 1;  //106 / 86 = 1
    16'b01101010_01010111 : OUT <= 1;  //106 / 87 = 1
    16'b01101010_01011000 : OUT <= 1;  //106 / 88 = 1
    16'b01101010_01011001 : OUT <= 1;  //106 / 89 = 1
    16'b01101010_01011010 : OUT <= 1;  //106 / 90 = 1
    16'b01101010_01011011 : OUT <= 1;  //106 / 91 = 1
    16'b01101010_01011100 : OUT <= 1;  //106 / 92 = 1
    16'b01101010_01011101 : OUT <= 1;  //106 / 93 = 1
    16'b01101010_01011110 : OUT <= 1;  //106 / 94 = 1
    16'b01101010_01011111 : OUT <= 1;  //106 / 95 = 1
    16'b01101010_01100000 : OUT <= 1;  //106 / 96 = 1
    16'b01101010_01100001 : OUT <= 1;  //106 / 97 = 1
    16'b01101010_01100010 : OUT <= 1;  //106 / 98 = 1
    16'b01101010_01100011 : OUT <= 1;  //106 / 99 = 1
    16'b01101010_01100100 : OUT <= 1;  //106 / 100 = 1
    16'b01101010_01100101 : OUT <= 1;  //106 / 101 = 1
    16'b01101010_01100110 : OUT <= 1;  //106 / 102 = 1
    16'b01101010_01100111 : OUT <= 1;  //106 / 103 = 1
    16'b01101010_01101000 : OUT <= 1;  //106 / 104 = 1
    16'b01101010_01101001 : OUT <= 1;  //106 / 105 = 1
    16'b01101010_01101010 : OUT <= 1;  //106 / 106 = 1
    16'b01101010_01101011 : OUT <= 0;  //106 / 107 = 0
    16'b01101010_01101100 : OUT <= 0;  //106 / 108 = 0
    16'b01101010_01101101 : OUT <= 0;  //106 / 109 = 0
    16'b01101010_01101110 : OUT <= 0;  //106 / 110 = 0
    16'b01101010_01101111 : OUT <= 0;  //106 / 111 = 0
    16'b01101010_01110000 : OUT <= 0;  //106 / 112 = 0
    16'b01101010_01110001 : OUT <= 0;  //106 / 113 = 0
    16'b01101010_01110010 : OUT <= 0;  //106 / 114 = 0
    16'b01101010_01110011 : OUT <= 0;  //106 / 115 = 0
    16'b01101010_01110100 : OUT <= 0;  //106 / 116 = 0
    16'b01101010_01110101 : OUT <= 0;  //106 / 117 = 0
    16'b01101010_01110110 : OUT <= 0;  //106 / 118 = 0
    16'b01101010_01110111 : OUT <= 0;  //106 / 119 = 0
    16'b01101010_01111000 : OUT <= 0;  //106 / 120 = 0
    16'b01101010_01111001 : OUT <= 0;  //106 / 121 = 0
    16'b01101010_01111010 : OUT <= 0;  //106 / 122 = 0
    16'b01101010_01111011 : OUT <= 0;  //106 / 123 = 0
    16'b01101010_01111100 : OUT <= 0;  //106 / 124 = 0
    16'b01101010_01111101 : OUT <= 0;  //106 / 125 = 0
    16'b01101010_01111110 : OUT <= 0;  //106 / 126 = 0
    16'b01101010_01111111 : OUT <= 0;  //106 / 127 = 0
    16'b01101010_10000000 : OUT <= 0;  //106 / 128 = 0
    16'b01101010_10000001 : OUT <= 0;  //106 / 129 = 0
    16'b01101010_10000010 : OUT <= 0;  //106 / 130 = 0
    16'b01101010_10000011 : OUT <= 0;  //106 / 131 = 0
    16'b01101010_10000100 : OUT <= 0;  //106 / 132 = 0
    16'b01101010_10000101 : OUT <= 0;  //106 / 133 = 0
    16'b01101010_10000110 : OUT <= 0;  //106 / 134 = 0
    16'b01101010_10000111 : OUT <= 0;  //106 / 135 = 0
    16'b01101010_10001000 : OUT <= 0;  //106 / 136 = 0
    16'b01101010_10001001 : OUT <= 0;  //106 / 137 = 0
    16'b01101010_10001010 : OUT <= 0;  //106 / 138 = 0
    16'b01101010_10001011 : OUT <= 0;  //106 / 139 = 0
    16'b01101010_10001100 : OUT <= 0;  //106 / 140 = 0
    16'b01101010_10001101 : OUT <= 0;  //106 / 141 = 0
    16'b01101010_10001110 : OUT <= 0;  //106 / 142 = 0
    16'b01101010_10001111 : OUT <= 0;  //106 / 143 = 0
    16'b01101010_10010000 : OUT <= 0;  //106 / 144 = 0
    16'b01101010_10010001 : OUT <= 0;  //106 / 145 = 0
    16'b01101010_10010010 : OUT <= 0;  //106 / 146 = 0
    16'b01101010_10010011 : OUT <= 0;  //106 / 147 = 0
    16'b01101010_10010100 : OUT <= 0;  //106 / 148 = 0
    16'b01101010_10010101 : OUT <= 0;  //106 / 149 = 0
    16'b01101010_10010110 : OUT <= 0;  //106 / 150 = 0
    16'b01101010_10010111 : OUT <= 0;  //106 / 151 = 0
    16'b01101010_10011000 : OUT <= 0;  //106 / 152 = 0
    16'b01101010_10011001 : OUT <= 0;  //106 / 153 = 0
    16'b01101010_10011010 : OUT <= 0;  //106 / 154 = 0
    16'b01101010_10011011 : OUT <= 0;  //106 / 155 = 0
    16'b01101010_10011100 : OUT <= 0;  //106 / 156 = 0
    16'b01101010_10011101 : OUT <= 0;  //106 / 157 = 0
    16'b01101010_10011110 : OUT <= 0;  //106 / 158 = 0
    16'b01101010_10011111 : OUT <= 0;  //106 / 159 = 0
    16'b01101010_10100000 : OUT <= 0;  //106 / 160 = 0
    16'b01101010_10100001 : OUT <= 0;  //106 / 161 = 0
    16'b01101010_10100010 : OUT <= 0;  //106 / 162 = 0
    16'b01101010_10100011 : OUT <= 0;  //106 / 163 = 0
    16'b01101010_10100100 : OUT <= 0;  //106 / 164 = 0
    16'b01101010_10100101 : OUT <= 0;  //106 / 165 = 0
    16'b01101010_10100110 : OUT <= 0;  //106 / 166 = 0
    16'b01101010_10100111 : OUT <= 0;  //106 / 167 = 0
    16'b01101010_10101000 : OUT <= 0;  //106 / 168 = 0
    16'b01101010_10101001 : OUT <= 0;  //106 / 169 = 0
    16'b01101010_10101010 : OUT <= 0;  //106 / 170 = 0
    16'b01101010_10101011 : OUT <= 0;  //106 / 171 = 0
    16'b01101010_10101100 : OUT <= 0;  //106 / 172 = 0
    16'b01101010_10101101 : OUT <= 0;  //106 / 173 = 0
    16'b01101010_10101110 : OUT <= 0;  //106 / 174 = 0
    16'b01101010_10101111 : OUT <= 0;  //106 / 175 = 0
    16'b01101010_10110000 : OUT <= 0;  //106 / 176 = 0
    16'b01101010_10110001 : OUT <= 0;  //106 / 177 = 0
    16'b01101010_10110010 : OUT <= 0;  //106 / 178 = 0
    16'b01101010_10110011 : OUT <= 0;  //106 / 179 = 0
    16'b01101010_10110100 : OUT <= 0;  //106 / 180 = 0
    16'b01101010_10110101 : OUT <= 0;  //106 / 181 = 0
    16'b01101010_10110110 : OUT <= 0;  //106 / 182 = 0
    16'b01101010_10110111 : OUT <= 0;  //106 / 183 = 0
    16'b01101010_10111000 : OUT <= 0;  //106 / 184 = 0
    16'b01101010_10111001 : OUT <= 0;  //106 / 185 = 0
    16'b01101010_10111010 : OUT <= 0;  //106 / 186 = 0
    16'b01101010_10111011 : OUT <= 0;  //106 / 187 = 0
    16'b01101010_10111100 : OUT <= 0;  //106 / 188 = 0
    16'b01101010_10111101 : OUT <= 0;  //106 / 189 = 0
    16'b01101010_10111110 : OUT <= 0;  //106 / 190 = 0
    16'b01101010_10111111 : OUT <= 0;  //106 / 191 = 0
    16'b01101010_11000000 : OUT <= 0;  //106 / 192 = 0
    16'b01101010_11000001 : OUT <= 0;  //106 / 193 = 0
    16'b01101010_11000010 : OUT <= 0;  //106 / 194 = 0
    16'b01101010_11000011 : OUT <= 0;  //106 / 195 = 0
    16'b01101010_11000100 : OUT <= 0;  //106 / 196 = 0
    16'b01101010_11000101 : OUT <= 0;  //106 / 197 = 0
    16'b01101010_11000110 : OUT <= 0;  //106 / 198 = 0
    16'b01101010_11000111 : OUT <= 0;  //106 / 199 = 0
    16'b01101010_11001000 : OUT <= 0;  //106 / 200 = 0
    16'b01101010_11001001 : OUT <= 0;  //106 / 201 = 0
    16'b01101010_11001010 : OUT <= 0;  //106 / 202 = 0
    16'b01101010_11001011 : OUT <= 0;  //106 / 203 = 0
    16'b01101010_11001100 : OUT <= 0;  //106 / 204 = 0
    16'b01101010_11001101 : OUT <= 0;  //106 / 205 = 0
    16'b01101010_11001110 : OUT <= 0;  //106 / 206 = 0
    16'b01101010_11001111 : OUT <= 0;  //106 / 207 = 0
    16'b01101010_11010000 : OUT <= 0;  //106 / 208 = 0
    16'b01101010_11010001 : OUT <= 0;  //106 / 209 = 0
    16'b01101010_11010010 : OUT <= 0;  //106 / 210 = 0
    16'b01101010_11010011 : OUT <= 0;  //106 / 211 = 0
    16'b01101010_11010100 : OUT <= 0;  //106 / 212 = 0
    16'b01101010_11010101 : OUT <= 0;  //106 / 213 = 0
    16'b01101010_11010110 : OUT <= 0;  //106 / 214 = 0
    16'b01101010_11010111 : OUT <= 0;  //106 / 215 = 0
    16'b01101010_11011000 : OUT <= 0;  //106 / 216 = 0
    16'b01101010_11011001 : OUT <= 0;  //106 / 217 = 0
    16'b01101010_11011010 : OUT <= 0;  //106 / 218 = 0
    16'b01101010_11011011 : OUT <= 0;  //106 / 219 = 0
    16'b01101010_11011100 : OUT <= 0;  //106 / 220 = 0
    16'b01101010_11011101 : OUT <= 0;  //106 / 221 = 0
    16'b01101010_11011110 : OUT <= 0;  //106 / 222 = 0
    16'b01101010_11011111 : OUT <= 0;  //106 / 223 = 0
    16'b01101010_11100000 : OUT <= 0;  //106 / 224 = 0
    16'b01101010_11100001 : OUT <= 0;  //106 / 225 = 0
    16'b01101010_11100010 : OUT <= 0;  //106 / 226 = 0
    16'b01101010_11100011 : OUT <= 0;  //106 / 227 = 0
    16'b01101010_11100100 : OUT <= 0;  //106 / 228 = 0
    16'b01101010_11100101 : OUT <= 0;  //106 / 229 = 0
    16'b01101010_11100110 : OUT <= 0;  //106 / 230 = 0
    16'b01101010_11100111 : OUT <= 0;  //106 / 231 = 0
    16'b01101010_11101000 : OUT <= 0;  //106 / 232 = 0
    16'b01101010_11101001 : OUT <= 0;  //106 / 233 = 0
    16'b01101010_11101010 : OUT <= 0;  //106 / 234 = 0
    16'b01101010_11101011 : OUT <= 0;  //106 / 235 = 0
    16'b01101010_11101100 : OUT <= 0;  //106 / 236 = 0
    16'b01101010_11101101 : OUT <= 0;  //106 / 237 = 0
    16'b01101010_11101110 : OUT <= 0;  //106 / 238 = 0
    16'b01101010_11101111 : OUT <= 0;  //106 / 239 = 0
    16'b01101010_11110000 : OUT <= 0;  //106 / 240 = 0
    16'b01101010_11110001 : OUT <= 0;  //106 / 241 = 0
    16'b01101010_11110010 : OUT <= 0;  //106 / 242 = 0
    16'b01101010_11110011 : OUT <= 0;  //106 / 243 = 0
    16'b01101010_11110100 : OUT <= 0;  //106 / 244 = 0
    16'b01101010_11110101 : OUT <= 0;  //106 / 245 = 0
    16'b01101010_11110110 : OUT <= 0;  //106 / 246 = 0
    16'b01101010_11110111 : OUT <= 0;  //106 / 247 = 0
    16'b01101010_11111000 : OUT <= 0;  //106 / 248 = 0
    16'b01101010_11111001 : OUT <= 0;  //106 / 249 = 0
    16'b01101010_11111010 : OUT <= 0;  //106 / 250 = 0
    16'b01101010_11111011 : OUT <= 0;  //106 / 251 = 0
    16'b01101010_11111100 : OUT <= 0;  //106 / 252 = 0
    16'b01101010_11111101 : OUT <= 0;  //106 / 253 = 0
    16'b01101010_11111110 : OUT <= 0;  //106 / 254 = 0
    16'b01101010_11111111 : OUT <= 0;  //106 / 255 = 0
    16'b01101011_00000000 : OUT <= 0;  //107 / 0 = 0
    16'b01101011_00000001 : OUT <= 107;  //107 / 1 = 107
    16'b01101011_00000010 : OUT <= 53;  //107 / 2 = 53
    16'b01101011_00000011 : OUT <= 35;  //107 / 3 = 35
    16'b01101011_00000100 : OUT <= 26;  //107 / 4 = 26
    16'b01101011_00000101 : OUT <= 21;  //107 / 5 = 21
    16'b01101011_00000110 : OUT <= 17;  //107 / 6 = 17
    16'b01101011_00000111 : OUT <= 15;  //107 / 7 = 15
    16'b01101011_00001000 : OUT <= 13;  //107 / 8 = 13
    16'b01101011_00001001 : OUT <= 11;  //107 / 9 = 11
    16'b01101011_00001010 : OUT <= 10;  //107 / 10 = 10
    16'b01101011_00001011 : OUT <= 9;  //107 / 11 = 9
    16'b01101011_00001100 : OUT <= 8;  //107 / 12 = 8
    16'b01101011_00001101 : OUT <= 8;  //107 / 13 = 8
    16'b01101011_00001110 : OUT <= 7;  //107 / 14 = 7
    16'b01101011_00001111 : OUT <= 7;  //107 / 15 = 7
    16'b01101011_00010000 : OUT <= 6;  //107 / 16 = 6
    16'b01101011_00010001 : OUT <= 6;  //107 / 17 = 6
    16'b01101011_00010010 : OUT <= 5;  //107 / 18 = 5
    16'b01101011_00010011 : OUT <= 5;  //107 / 19 = 5
    16'b01101011_00010100 : OUT <= 5;  //107 / 20 = 5
    16'b01101011_00010101 : OUT <= 5;  //107 / 21 = 5
    16'b01101011_00010110 : OUT <= 4;  //107 / 22 = 4
    16'b01101011_00010111 : OUT <= 4;  //107 / 23 = 4
    16'b01101011_00011000 : OUT <= 4;  //107 / 24 = 4
    16'b01101011_00011001 : OUT <= 4;  //107 / 25 = 4
    16'b01101011_00011010 : OUT <= 4;  //107 / 26 = 4
    16'b01101011_00011011 : OUT <= 3;  //107 / 27 = 3
    16'b01101011_00011100 : OUT <= 3;  //107 / 28 = 3
    16'b01101011_00011101 : OUT <= 3;  //107 / 29 = 3
    16'b01101011_00011110 : OUT <= 3;  //107 / 30 = 3
    16'b01101011_00011111 : OUT <= 3;  //107 / 31 = 3
    16'b01101011_00100000 : OUT <= 3;  //107 / 32 = 3
    16'b01101011_00100001 : OUT <= 3;  //107 / 33 = 3
    16'b01101011_00100010 : OUT <= 3;  //107 / 34 = 3
    16'b01101011_00100011 : OUT <= 3;  //107 / 35 = 3
    16'b01101011_00100100 : OUT <= 2;  //107 / 36 = 2
    16'b01101011_00100101 : OUT <= 2;  //107 / 37 = 2
    16'b01101011_00100110 : OUT <= 2;  //107 / 38 = 2
    16'b01101011_00100111 : OUT <= 2;  //107 / 39 = 2
    16'b01101011_00101000 : OUT <= 2;  //107 / 40 = 2
    16'b01101011_00101001 : OUT <= 2;  //107 / 41 = 2
    16'b01101011_00101010 : OUT <= 2;  //107 / 42 = 2
    16'b01101011_00101011 : OUT <= 2;  //107 / 43 = 2
    16'b01101011_00101100 : OUT <= 2;  //107 / 44 = 2
    16'b01101011_00101101 : OUT <= 2;  //107 / 45 = 2
    16'b01101011_00101110 : OUT <= 2;  //107 / 46 = 2
    16'b01101011_00101111 : OUT <= 2;  //107 / 47 = 2
    16'b01101011_00110000 : OUT <= 2;  //107 / 48 = 2
    16'b01101011_00110001 : OUT <= 2;  //107 / 49 = 2
    16'b01101011_00110010 : OUT <= 2;  //107 / 50 = 2
    16'b01101011_00110011 : OUT <= 2;  //107 / 51 = 2
    16'b01101011_00110100 : OUT <= 2;  //107 / 52 = 2
    16'b01101011_00110101 : OUT <= 2;  //107 / 53 = 2
    16'b01101011_00110110 : OUT <= 1;  //107 / 54 = 1
    16'b01101011_00110111 : OUT <= 1;  //107 / 55 = 1
    16'b01101011_00111000 : OUT <= 1;  //107 / 56 = 1
    16'b01101011_00111001 : OUT <= 1;  //107 / 57 = 1
    16'b01101011_00111010 : OUT <= 1;  //107 / 58 = 1
    16'b01101011_00111011 : OUT <= 1;  //107 / 59 = 1
    16'b01101011_00111100 : OUT <= 1;  //107 / 60 = 1
    16'b01101011_00111101 : OUT <= 1;  //107 / 61 = 1
    16'b01101011_00111110 : OUT <= 1;  //107 / 62 = 1
    16'b01101011_00111111 : OUT <= 1;  //107 / 63 = 1
    16'b01101011_01000000 : OUT <= 1;  //107 / 64 = 1
    16'b01101011_01000001 : OUT <= 1;  //107 / 65 = 1
    16'b01101011_01000010 : OUT <= 1;  //107 / 66 = 1
    16'b01101011_01000011 : OUT <= 1;  //107 / 67 = 1
    16'b01101011_01000100 : OUT <= 1;  //107 / 68 = 1
    16'b01101011_01000101 : OUT <= 1;  //107 / 69 = 1
    16'b01101011_01000110 : OUT <= 1;  //107 / 70 = 1
    16'b01101011_01000111 : OUT <= 1;  //107 / 71 = 1
    16'b01101011_01001000 : OUT <= 1;  //107 / 72 = 1
    16'b01101011_01001001 : OUT <= 1;  //107 / 73 = 1
    16'b01101011_01001010 : OUT <= 1;  //107 / 74 = 1
    16'b01101011_01001011 : OUT <= 1;  //107 / 75 = 1
    16'b01101011_01001100 : OUT <= 1;  //107 / 76 = 1
    16'b01101011_01001101 : OUT <= 1;  //107 / 77 = 1
    16'b01101011_01001110 : OUT <= 1;  //107 / 78 = 1
    16'b01101011_01001111 : OUT <= 1;  //107 / 79 = 1
    16'b01101011_01010000 : OUT <= 1;  //107 / 80 = 1
    16'b01101011_01010001 : OUT <= 1;  //107 / 81 = 1
    16'b01101011_01010010 : OUT <= 1;  //107 / 82 = 1
    16'b01101011_01010011 : OUT <= 1;  //107 / 83 = 1
    16'b01101011_01010100 : OUT <= 1;  //107 / 84 = 1
    16'b01101011_01010101 : OUT <= 1;  //107 / 85 = 1
    16'b01101011_01010110 : OUT <= 1;  //107 / 86 = 1
    16'b01101011_01010111 : OUT <= 1;  //107 / 87 = 1
    16'b01101011_01011000 : OUT <= 1;  //107 / 88 = 1
    16'b01101011_01011001 : OUT <= 1;  //107 / 89 = 1
    16'b01101011_01011010 : OUT <= 1;  //107 / 90 = 1
    16'b01101011_01011011 : OUT <= 1;  //107 / 91 = 1
    16'b01101011_01011100 : OUT <= 1;  //107 / 92 = 1
    16'b01101011_01011101 : OUT <= 1;  //107 / 93 = 1
    16'b01101011_01011110 : OUT <= 1;  //107 / 94 = 1
    16'b01101011_01011111 : OUT <= 1;  //107 / 95 = 1
    16'b01101011_01100000 : OUT <= 1;  //107 / 96 = 1
    16'b01101011_01100001 : OUT <= 1;  //107 / 97 = 1
    16'b01101011_01100010 : OUT <= 1;  //107 / 98 = 1
    16'b01101011_01100011 : OUT <= 1;  //107 / 99 = 1
    16'b01101011_01100100 : OUT <= 1;  //107 / 100 = 1
    16'b01101011_01100101 : OUT <= 1;  //107 / 101 = 1
    16'b01101011_01100110 : OUT <= 1;  //107 / 102 = 1
    16'b01101011_01100111 : OUT <= 1;  //107 / 103 = 1
    16'b01101011_01101000 : OUT <= 1;  //107 / 104 = 1
    16'b01101011_01101001 : OUT <= 1;  //107 / 105 = 1
    16'b01101011_01101010 : OUT <= 1;  //107 / 106 = 1
    16'b01101011_01101011 : OUT <= 1;  //107 / 107 = 1
    16'b01101011_01101100 : OUT <= 0;  //107 / 108 = 0
    16'b01101011_01101101 : OUT <= 0;  //107 / 109 = 0
    16'b01101011_01101110 : OUT <= 0;  //107 / 110 = 0
    16'b01101011_01101111 : OUT <= 0;  //107 / 111 = 0
    16'b01101011_01110000 : OUT <= 0;  //107 / 112 = 0
    16'b01101011_01110001 : OUT <= 0;  //107 / 113 = 0
    16'b01101011_01110010 : OUT <= 0;  //107 / 114 = 0
    16'b01101011_01110011 : OUT <= 0;  //107 / 115 = 0
    16'b01101011_01110100 : OUT <= 0;  //107 / 116 = 0
    16'b01101011_01110101 : OUT <= 0;  //107 / 117 = 0
    16'b01101011_01110110 : OUT <= 0;  //107 / 118 = 0
    16'b01101011_01110111 : OUT <= 0;  //107 / 119 = 0
    16'b01101011_01111000 : OUT <= 0;  //107 / 120 = 0
    16'b01101011_01111001 : OUT <= 0;  //107 / 121 = 0
    16'b01101011_01111010 : OUT <= 0;  //107 / 122 = 0
    16'b01101011_01111011 : OUT <= 0;  //107 / 123 = 0
    16'b01101011_01111100 : OUT <= 0;  //107 / 124 = 0
    16'b01101011_01111101 : OUT <= 0;  //107 / 125 = 0
    16'b01101011_01111110 : OUT <= 0;  //107 / 126 = 0
    16'b01101011_01111111 : OUT <= 0;  //107 / 127 = 0
    16'b01101011_10000000 : OUT <= 0;  //107 / 128 = 0
    16'b01101011_10000001 : OUT <= 0;  //107 / 129 = 0
    16'b01101011_10000010 : OUT <= 0;  //107 / 130 = 0
    16'b01101011_10000011 : OUT <= 0;  //107 / 131 = 0
    16'b01101011_10000100 : OUT <= 0;  //107 / 132 = 0
    16'b01101011_10000101 : OUT <= 0;  //107 / 133 = 0
    16'b01101011_10000110 : OUT <= 0;  //107 / 134 = 0
    16'b01101011_10000111 : OUT <= 0;  //107 / 135 = 0
    16'b01101011_10001000 : OUT <= 0;  //107 / 136 = 0
    16'b01101011_10001001 : OUT <= 0;  //107 / 137 = 0
    16'b01101011_10001010 : OUT <= 0;  //107 / 138 = 0
    16'b01101011_10001011 : OUT <= 0;  //107 / 139 = 0
    16'b01101011_10001100 : OUT <= 0;  //107 / 140 = 0
    16'b01101011_10001101 : OUT <= 0;  //107 / 141 = 0
    16'b01101011_10001110 : OUT <= 0;  //107 / 142 = 0
    16'b01101011_10001111 : OUT <= 0;  //107 / 143 = 0
    16'b01101011_10010000 : OUT <= 0;  //107 / 144 = 0
    16'b01101011_10010001 : OUT <= 0;  //107 / 145 = 0
    16'b01101011_10010010 : OUT <= 0;  //107 / 146 = 0
    16'b01101011_10010011 : OUT <= 0;  //107 / 147 = 0
    16'b01101011_10010100 : OUT <= 0;  //107 / 148 = 0
    16'b01101011_10010101 : OUT <= 0;  //107 / 149 = 0
    16'b01101011_10010110 : OUT <= 0;  //107 / 150 = 0
    16'b01101011_10010111 : OUT <= 0;  //107 / 151 = 0
    16'b01101011_10011000 : OUT <= 0;  //107 / 152 = 0
    16'b01101011_10011001 : OUT <= 0;  //107 / 153 = 0
    16'b01101011_10011010 : OUT <= 0;  //107 / 154 = 0
    16'b01101011_10011011 : OUT <= 0;  //107 / 155 = 0
    16'b01101011_10011100 : OUT <= 0;  //107 / 156 = 0
    16'b01101011_10011101 : OUT <= 0;  //107 / 157 = 0
    16'b01101011_10011110 : OUT <= 0;  //107 / 158 = 0
    16'b01101011_10011111 : OUT <= 0;  //107 / 159 = 0
    16'b01101011_10100000 : OUT <= 0;  //107 / 160 = 0
    16'b01101011_10100001 : OUT <= 0;  //107 / 161 = 0
    16'b01101011_10100010 : OUT <= 0;  //107 / 162 = 0
    16'b01101011_10100011 : OUT <= 0;  //107 / 163 = 0
    16'b01101011_10100100 : OUT <= 0;  //107 / 164 = 0
    16'b01101011_10100101 : OUT <= 0;  //107 / 165 = 0
    16'b01101011_10100110 : OUT <= 0;  //107 / 166 = 0
    16'b01101011_10100111 : OUT <= 0;  //107 / 167 = 0
    16'b01101011_10101000 : OUT <= 0;  //107 / 168 = 0
    16'b01101011_10101001 : OUT <= 0;  //107 / 169 = 0
    16'b01101011_10101010 : OUT <= 0;  //107 / 170 = 0
    16'b01101011_10101011 : OUT <= 0;  //107 / 171 = 0
    16'b01101011_10101100 : OUT <= 0;  //107 / 172 = 0
    16'b01101011_10101101 : OUT <= 0;  //107 / 173 = 0
    16'b01101011_10101110 : OUT <= 0;  //107 / 174 = 0
    16'b01101011_10101111 : OUT <= 0;  //107 / 175 = 0
    16'b01101011_10110000 : OUT <= 0;  //107 / 176 = 0
    16'b01101011_10110001 : OUT <= 0;  //107 / 177 = 0
    16'b01101011_10110010 : OUT <= 0;  //107 / 178 = 0
    16'b01101011_10110011 : OUT <= 0;  //107 / 179 = 0
    16'b01101011_10110100 : OUT <= 0;  //107 / 180 = 0
    16'b01101011_10110101 : OUT <= 0;  //107 / 181 = 0
    16'b01101011_10110110 : OUT <= 0;  //107 / 182 = 0
    16'b01101011_10110111 : OUT <= 0;  //107 / 183 = 0
    16'b01101011_10111000 : OUT <= 0;  //107 / 184 = 0
    16'b01101011_10111001 : OUT <= 0;  //107 / 185 = 0
    16'b01101011_10111010 : OUT <= 0;  //107 / 186 = 0
    16'b01101011_10111011 : OUT <= 0;  //107 / 187 = 0
    16'b01101011_10111100 : OUT <= 0;  //107 / 188 = 0
    16'b01101011_10111101 : OUT <= 0;  //107 / 189 = 0
    16'b01101011_10111110 : OUT <= 0;  //107 / 190 = 0
    16'b01101011_10111111 : OUT <= 0;  //107 / 191 = 0
    16'b01101011_11000000 : OUT <= 0;  //107 / 192 = 0
    16'b01101011_11000001 : OUT <= 0;  //107 / 193 = 0
    16'b01101011_11000010 : OUT <= 0;  //107 / 194 = 0
    16'b01101011_11000011 : OUT <= 0;  //107 / 195 = 0
    16'b01101011_11000100 : OUT <= 0;  //107 / 196 = 0
    16'b01101011_11000101 : OUT <= 0;  //107 / 197 = 0
    16'b01101011_11000110 : OUT <= 0;  //107 / 198 = 0
    16'b01101011_11000111 : OUT <= 0;  //107 / 199 = 0
    16'b01101011_11001000 : OUT <= 0;  //107 / 200 = 0
    16'b01101011_11001001 : OUT <= 0;  //107 / 201 = 0
    16'b01101011_11001010 : OUT <= 0;  //107 / 202 = 0
    16'b01101011_11001011 : OUT <= 0;  //107 / 203 = 0
    16'b01101011_11001100 : OUT <= 0;  //107 / 204 = 0
    16'b01101011_11001101 : OUT <= 0;  //107 / 205 = 0
    16'b01101011_11001110 : OUT <= 0;  //107 / 206 = 0
    16'b01101011_11001111 : OUT <= 0;  //107 / 207 = 0
    16'b01101011_11010000 : OUT <= 0;  //107 / 208 = 0
    16'b01101011_11010001 : OUT <= 0;  //107 / 209 = 0
    16'b01101011_11010010 : OUT <= 0;  //107 / 210 = 0
    16'b01101011_11010011 : OUT <= 0;  //107 / 211 = 0
    16'b01101011_11010100 : OUT <= 0;  //107 / 212 = 0
    16'b01101011_11010101 : OUT <= 0;  //107 / 213 = 0
    16'b01101011_11010110 : OUT <= 0;  //107 / 214 = 0
    16'b01101011_11010111 : OUT <= 0;  //107 / 215 = 0
    16'b01101011_11011000 : OUT <= 0;  //107 / 216 = 0
    16'b01101011_11011001 : OUT <= 0;  //107 / 217 = 0
    16'b01101011_11011010 : OUT <= 0;  //107 / 218 = 0
    16'b01101011_11011011 : OUT <= 0;  //107 / 219 = 0
    16'b01101011_11011100 : OUT <= 0;  //107 / 220 = 0
    16'b01101011_11011101 : OUT <= 0;  //107 / 221 = 0
    16'b01101011_11011110 : OUT <= 0;  //107 / 222 = 0
    16'b01101011_11011111 : OUT <= 0;  //107 / 223 = 0
    16'b01101011_11100000 : OUT <= 0;  //107 / 224 = 0
    16'b01101011_11100001 : OUT <= 0;  //107 / 225 = 0
    16'b01101011_11100010 : OUT <= 0;  //107 / 226 = 0
    16'b01101011_11100011 : OUT <= 0;  //107 / 227 = 0
    16'b01101011_11100100 : OUT <= 0;  //107 / 228 = 0
    16'b01101011_11100101 : OUT <= 0;  //107 / 229 = 0
    16'b01101011_11100110 : OUT <= 0;  //107 / 230 = 0
    16'b01101011_11100111 : OUT <= 0;  //107 / 231 = 0
    16'b01101011_11101000 : OUT <= 0;  //107 / 232 = 0
    16'b01101011_11101001 : OUT <= 0;  //107 / 233 = 0
    16'b01101011_11101010 : OUT <= 0;  //107 / 234 = 0
    16'b01101011_11101011 : OUT <= 0;  //107 / 235 = 0
    16'b01101011_11101100 : OUT <= 0;  //107 / 236 = 0
    16'b01101011_11101101 : OUT <= 0;  //107 / 237 = 0
    16'b01101011_11101110 : OUT <= 0;  //107 / 238 = 0
    16'b01101011_11101111 : OUT <= 0;  //107 / 239 = 0
    16'b01101011_11110000 : OUT <= 0;  //107 / 240 = 0
    16'b01101011_11110001 : OUT <= 0;  //107 / 241 = 0
    16'b01101011_11110010 : OUT <= 0;  //107 / 242 = 0
    16'b01101011_11110011 : OUT <= 0;  //107 / 243 = 0
    16'b01101011_11110100 : OUT <= 0;  //107 / 244 = 0
    16'b01101011_11110101 : OUT <= 0;  //107 / 245 = 0
    16'b01101011_11110110 : OUT <= 0;  //107 / 246 = 0
    16'b01101011_11110111 : OUT <= 0;  //107 / 247 = 0
    16'b01101011_11111000 : OUT <= 0;  //107 / 248 = 0
    16'b01101011_11111001 : OUT <= 0;  //107 / 249 = 0
    16'b01101011_11111010 : OUT <= 0;  //107 / 250 = 0
    16'b01101011_11111011 : OUT <= 0;  //107 / 251 = 0
    16'b01101011_11111100 : OUT <= 0;  //107 / 252 = 0
    16'b01101011_11111101 : OUT <= 0;  //107 / 253 = 0
    16'b01101011_11111110 : OUT <= 0;  //107 / 254 = 0
    16'b01101011_11111111 : OUT <= 0;  //107 / 255 = 0
    16'b01101100_00000000 : OUT <= 0;  //108 / 0 = 0
    16'b01101100_00000001 : OUT <= 108;  //108 / 1 = 108
    16'b01101100_00000010 : OUT <= 54;  //108 / 2 = 54
    16'b01101100_00000011 : OUT <= 36;  //108 / 3 = 36
    16'b01101100_00000100 : OUT <= 27;  //108 / 4 = 27
    16'b01101100_00000101 : OUT <= 21;  //108 / 5 = 21
    16'b01101100_00000110 : OUT <= 18;  //108 / 6 = 18
    16'b01101100_00000111 : OUT <= 15;  //108 / 7 = 15
    16'b01101100_00001000 : OUT <= 13;  //108 / 8 = 13
    16'b01101100_00001001 : OUT <= 12;  //108 / 9 = 12
    16'b01101100_00001010 : OUT <= 10;  //108 / 10 = 10
    16'b01101100_00001011 : OUT <= 9;  //108 / 11 = 9
    16'b01101100_00001100 : OUT <= 9;  //108 / 12 = 9
    16'b01101100_00001101 : OUT <= 8;  //108 / 13 = 8
    16'b01101100_00001110 : OUT <= 7;  //108 / 14 = 7
    16'b01101100_00001111 : OUT <= 7;  //108 / 15 = 7
    16'b01101100_00010000 : OUT <= 6;  //108 / 16 = 6
    16'b01101100_00010001 : OUT <= 6;  //108 / 17 = 6
    16'b01101100_00010010 : OUT <= 6;  //108 / 18 = 6
    16'b01101100_00010011 : OUT <= 5;  //108 / 19 = 5
    16'b01101100_00010100 : OUT <= 5;  //108 / 20 = 5
    16'b01101100_00010101 : OUT <= 5;  //108 / 21 = 5
    16'b01101100_00010110 : OUT <= 4;  //108 / 22 = 4
    16'b01101100_00010111 : OUT <= 4;  //108 / 23 = 4
    16'b01101100_00011000 : OUT <= 4;  //108 / 24 = 4
    16'b01101100_00011001 : OUT <= 4;  //108 / 25 = 4
    16'b01101100_00011010 : OUT <= 4;  //108 / 26 = 4
    16'b01101100_00011011 : OUT <= 4;  //108 / 27 = 4
    16'b01101100_00011100 : OUT <= 3;  //108 / 28 = 3
    16'b01101100_00011101 : OUT <= 3;  //108 / 29 = 3
    16'b01101100_00011110 : OUT <= 3;  //108 / 30 = 3
    16'b01101100_00011111 : OUT <= 3;  //108 / 31 = 3
    16'b01101100_00100000 : OUT <= 3;  //108 / 32 = 3
    16'b01101100_00100001 : OUT <= 3;  //108 / 33 = 3
    16'b01101100_00100010 : OUT <= 3;  //108 / 34 = 3
    16'b01101100_00100011 : OUT <= 3;  //108 / 35 = 3
    16'b01101100_00100100 : OUT <= 3;  //108 / 36 = 3
    16'b01101100_00100101 : OUT <= 2;  //108 / 37 = 2
    16'b01101100_00100110 : OUT <= 2;  //108 / 38 = 2
    16'b01101100_00100111 : OUT <= 2;  //108 / 39 = 2
    16'b01101100_00101000 : OUT <= 2;  //108 / 40 = 2
    16'b01101100_00101001 : OUT <= 2;  //108 / 41 = 2
    16'b01101100_00101010 : OUT <= 2;  //108 / 42 = 2
    16'b01101100_00101011 : OUT <= 2;  //108 / 43 = 2
    16'b01101100_00101100 : OUT <= 2;  //108 / 44 = 2
    16'b01101100_00101101 : OUT <= 2;  //108 / 45 = 2
    16'b01101100_00101110 : OUT <= 2;  //108 / 46 = 2
    16'b01101100_00101111 : OUT <= 2;  //108 / 47 = 2
    16'b01101100_00110000 : OUT <= 2;  //108 / 48 = 2
    16'b01101100_00110001 : OUT <= 2;  //108 / 49 = 2
    16'b01101100_00110010 : OUT <= 2;  //108 / 50 = 2
    16'b01101100_00110011 : OUT <= 2;  //108 / 51 = 2
    16'b01101100_00110100 : OUT <= 2;  //108 / 52 = 2
    16'b01101100_00110101 : OUT <= 2;  //108 / 53 = 2
    16'b01101100_00110110 : OUT <= 2;  //108 / 54 = 2
    16'b01101100_00110111 : OUT <= 1;  //108 / 55 = 1
    16'b01101100_00111000 : OUT <= 1;  //108 / 56 = 1
    16'b01101100_00111001 : OUT <= 1;  //108 / 57 = 1
    16'b01101100_00111010 : OUT <= 1;  //108 / 58 = 1
    16'b01101100_00111011 : OUT <= 1;  //108 / 59 = 1
    16'b01101100_00111100 : OUT <= 1;  //108 / 60 = 1
    16'b01101100_00111101 : OUT <= 1;  //108 / 61 = 1
    16'b01101100_00111110 : OUT <= 1;  //108 / 62 = 1
    16'b01101100_00111111 : OUT <= 1;  //108 / 63 = 1
    16'b01101100_01000000 : OUT <= 1;  //108 / 64 = 1
    16'b01101100_01000001 : OUT <= 1;  //108 / 65 = 1
    16'b01101100_01000010 : OUT <= 1;  //108 / 66 = 1
    16'b01101100_01000011 : OUT <= 1;  //108 / 67 = 1
    16'b01101100_01000100 : OUT <= 1;  //108 / 68 = 1
    16'b01101100_01000101 : OUT <= 1;  //108 / 69 = 1
    16'b01101100_01000110 : OUT <= 1;  //108 / 70 = 1
    16'b01101100_01000111 : OUT <= 1;  //108 / 71 = 1
    16'b01101100_01001000 : OUT <= 1;  //108 / 72 = 1
    16'b01101100_01001001 : OUT <= 1;  //108 / 73 = 1
    16'b01101100_01001010 : OUT <= 1;  //108 / 74 = 1
    16'b01101100_01001011 : OUT <= 1;  //108 / 75 = 1
    16'b01101100_01001100 : OUT <= 1;  //108 / 76 = 1
    16'b01101100_01001101 : OUT <= 1;  //108 / 77 = 1
    16'b01101100_01001110 : OUT <= 1;  //108 / 78 = 1
    16'b01101100_01001111 : OUT <= 1;  //108 / 79 = 1
    16'b01101100_01010000 : OUT <= 1;  //108 / 80 = 1
    16'b01101100_01010001 : OUT <= 1;  //108 / 81 = 1
    16'b01101100_01010010 : OUT <= 1;  //108 / 82 = 1
    16'b01101100_01010011 : OUT <= 1;  //108 / 83 = 1
    16'b01101100_01010100 : OUT <= 1;  //108 / 84 = 1
    16'b01101100_01010101 : OUT <= 1;  //108 / 85 = 1
    16'b01101100_01010110 : OUT <= 1;  //108 / 86 = 1
    16'b01101100_01010111 : OUT <= 1;  //108 / 87 = 1
    16'b01101100_01011000 : OUT <= 1;  //108 / 88 = 1
    16'b01101100_01011001 : OUT <= 1;  //108 / 89 = 1
    16'b01101100_01011010 : OUT <= 1;  //108 / 90 = 1
    16'b01101100_01011011 : OUT <= 1;  //108 / 91 = 1
    16'b01101100_01011100 : OUT <= 1;  //108 / 92 = 1
    16'b01101100_01011101 : OUT <= 1;  //108 / 93 = 1
    16'b01101100_01011110 : OUT <= 1;  //108 / 94 = 1
    16'b01101100_01011111 : OUT <= 1;  //108 / 95 = 1
    16'b01101100_01100000 : OUT <= 1;  //108 / 96 = 1
    16'b01101100_01100001 : OUT <= 1;  //108 / 97 = 1
    16'b01101100_01100010 : OUT <= 1;  //108 / 98 = 1
    16'b01101100_01100011 : OUT <= 1;  //108 / 99 = 1
    16'b01101100_01100100 : OUT <= 1;  //108 / 100 = 1
    16'b01101100_01100101 : OUT <= 1;  //108 / 101 = 1
    16'b01101100_01100110 : OUT <= 1;  //108 / 102 = 1
    16'b01101100_01100111 : OUT <= 1;  //108 / 103 = 1
    16'b01101100_01101000 : OUT <= 1;  //108 / 104 = 1
    16'b01101100_01101001 : OUT <= 1;  //108 / 105 = 1
    16'b01101100_01101010 : OUT <= 1;  //108 / 106 = 1
    16'b01101100_01101011 : OUT <= 1;  //108 / 107 = 1
    16'b01101100_01101100 : OUT <= 1;  //108 / 108 = 1
    16'b01101100_01101101 : OUT <= 0;  //108 / 109 = 0
    16'b01101100_01101110 : OUT <= 0;  //108 / 110 = 0
    16'b01101100_01101111 : OUT <= 0;  //108 / 111 = 0
    16'b01101100_01110000 : OUT <= 0;  //108 / 112 = 0
    16'b01101100_01110001 : OUT <= 0;  //108 / 113 = 0
    16'b01101100_01110010 : OUT <= 0;  //108 / 114 = 0
    16'b01101100_01110011 : OUT <= 0;  //108 / 115 = 0
    16'b01101100_01110100 : OUT <= 0;  //108 / 116 = 0
    16'b01101100_01110101 : OUT <= 0;  //108 / 117 = 0
    16'b01101100_01110110 : OUT <= 0;  //108 / 118 = 0
    16'b01101100_01110111 : OUT <= 0;  //108 / 119 = 0
    16'b01101100_01111000 : OUT <= 0;  //108 / 120 = 0
    16'b01101100_01111001 : OUT <= 0;  //108 / 121 = 0
    16'b01101100_01111010 : OUT <= 0;  //108 / 122 = 0
    16'b01101100_01111011 : OUT <= 0;  //108 / 123 = 0
    16'b01101100_01111100 : OUT <= 0;  //108 / 124 = 0
    16'b01101100_01111101 : OUT <= 0;  //108 / 125 = 0
    16'b01101100_01111110 : OUT <= 0;  //108 / 126 = 0
    16'b01101100_01111111 : OUT <= 0;  //108 / 127 = 0
    16'b01101100_10000000 : OUT <= 0;  //108 / 128 = 0
    16'b01101100_10000001 : OUT <= 0;  //108 / 129 = 0
    16'b01101100_10000010 : OUT <= 0;  //108 / 130 = 0
    16'b01101100_10000011 : OUT <= 0;  //108 / 131 = 0
    16'b01101100_10000100 : OUT <= 0;  //108 / 132 = 0
    16'b01101100_10000101 : OUT <= 0;  //108 / 133 = 0
    16'b01101100_10000110 : OUT <= 0;  //108 / 134 = 0
    16'b01101100_10000111 : OUT <= 0;  //108 / 135 = 0
    16'b01101100_10001000 : OUT <= 0;  //108 / 136 = 0
    16'b01101100_10001001 : OUT <= 0;  //108 / 137 = 0
    16'b01101100_10001010 : OUT <= 0;  //108 / 138 = 0
    16'b01101100_10001011 : OUT <= 0;  //108 / 139 = 0
    16'b01101100_10001100 : OUT <= 0;  //108 / 140 = 0
    16'b01101100_10001101 : OUT <= 0;  //108 / 141 = 0
    16'b01101100_10001110 : OUT <= 0;  //108 / 142 = 0
    16'b01101100_10001111 : OUT <= 0;  //108 / 143 = 0
    16'b01101100_10010000 : OUT <= 0;  //108 / 144 = 0
    16'b01101100_10010001 : OUT <= 0;  //108 / 145 = 0
    16'b01101100_10010010 : OUT <= 0;  //108 / 146 = 0
    16'b01101100_10010011 : OUT <= 0;  //108 / 147 = 0
    16'b01101100_10010100 : OUT <= 0;  //108 / 148 = 0
    16'b01101100_10010101 : OUT <= 0;  //108 / 149 = 0
    16'b01101100_10010110 : OUT <= 0;  //108 / 150 = 0
    16'b01101100_10010111 : OUT <= 0;  //108 / 151 = 0
    16'b01101100_10011000 : OUT <= 0;  //108 / 152 = 0
    16'b01101100_10011001 : OUT <= 0;  //108 / 153 = 0
    16'b01101100_10011010 : OUT <= 0;  //108 / 154 = 0
    16'b01101100_10011011 : OUT <= 0;  //108 / 155 = 0
    16'b01101100_10011100 : OUT <= 0;  //108 / 156 = 0
    16'b01101100_10011101 : OUT <= 0;  //108 / 157 = 0
    16'b01101100_10011110 : OUT <= 0;  //108 / 158 = 0
    16'b01101100_10011111 : OUT <= 0;  //108 / 159 = 0
    16'b01101100_10100000 : OUT <= 0;  //108 / 160 = 0
    16'b01101100_10100001 : OUT <= 0;  //108 / 161 = 0
    16'b01101100_10100010 : OUT <= 0;  //108 / 162 = 0
    16'b01101100_10100011 : OUT <= 0;  //108 / 163 = 0
    16'b01101100_10100100 : OUT <= 0;  //108 / 164 = 0
    16'b01101100_10100101 : OUT <= 0;  //108 / 165 = 0
    16'b01101100_10100110 : OUT <= 0;  //108 / 166 = 0
    16'b01101100_10100111 : OUT <= 0;  //108 / 167 = 0
    16'b01101100_10101000 : OUT <= 0;  //108 / 168 = 0
    16'b01101100_10101001 : OUT <= 0;  //108 / 169 = 0
    16'b01101100_10101010 : OUT <= 0;  //108 / 170 = 0
    16'b01101100_10101011 : OUT <= 0;  //108 / 171 = 0
    16'b01101100_10101100 : OUT <= 0;  //108 / 172 = 0
    16'b01101100_10101101 : OUT <= 0;  //108 / 173 = 0
    16'b01101100_10101110 : OUT <= 0;  //108 / 174 = 0
    16'b01101100_10101111 : OUT <= 0;  //108 / 175 = 0
    16'b01101100_10110000 : OUT <= 0;  //108 / 176 = 0
    16'b01101100_10110001 : OUT <= 0;  //108 / 177 = 0
    16'b01101100_10110010 : OUT <= 0;  //108 / 178 = 0
    16'b01101100_10110011 : OUT <= 0;  //108 / 179 = 0
    16'b01101100_10110100 : OUT <= 0;  //108 / 180 = 0
    16'b01101100_10110101 : OUT <= 0;  //108 / 181 = 0
    16'b01101100_10110110 : OUT <= 0;  //108 / 182 = 0
    16'b01101100_10110111 : OUT <= 0;  //108 / 183 = 0
    16'b01101100_10111000 : OUT <= 0;  //108 / 184 = 0
    16'b01101100_10111001 : OUT <= 0;  //108 / 185 = 0
    16'b01101100_10111010 : OUT <= 0;  //108 / 186 = 0
    16'b01101100_10111011 : OUT <= 0;  //108 / 187 = 0
    16'b01101100_10111100 : OUT <= 0;  //108 / 188 = 0
    16'b01101100_10111101 : OUT <= 0;  //108 / 189 = 0
    16'b01101100_10111110 : OUT <= 0;  //108 / 190 = 0
    16'b01101100_10111111 : OUT <= 0;  //108 / 191 = 0
    16'b01101100_11000000 : OUT <= 0;  //108 / 192 = 0
    16'b01101100_11000001 : OUT <= 0;  //108 / 193 = 0
    16'b01101100_11000010 : OUT <= 0;  //108 / 194 = 0
    16'b01101100_11000011 : OUT <= 0;  //108 / 195 = 0
    16'b01101100_11000100 : OUT <= 0;  //108 / 196 = 0
    16'b01101100_11000101 : OUT <= 0;  //108 / 197 = 0
    16'b01101100_11000110 : OUT <= 0;  //108 / 198 = 0
    16'b01101100_11000111 : OUT <= 0;  //108 / 199 = 0
    16'b01101100_11001000 : OUT <= 0;  //108 / 200 = 0
    16'b01101100_11001001 : OUT <= 0;  //108 / 201 = 0
    16'b01101100_11001010 : OUT <= 0;  //108 / 202 = 0
    16'b01101100_11001011 : OUT <= 0;  //108 / 203 = 0
    16'b01101100_11001100 : OUT <= 0;  //108 / 204 = 0
    16'b01101100_11001101 : OUT <= 0;  //108 / 205 = 0
    16'b01101100_11001110 : OUT <= 0;  //108 / 206 = 0
    16'b01101100_11001111 : OUT <= 0;  //108 / 207 = 0
    16'b01101100_11010000 : OUT <= 0;  //108 / 208 = 0
    16'b01101100_11010001 : OUT <= 0;  //108 / 209 = 0
    16'b01101100_11010010 : OUT <= 0;  //108 / 210 = 0
    16'b01101100_11010011 : OUT <= 0;  //108 / 211 = 0
    16'b01101100_11010100 : OUT <= 0;  //108 / 212 = 0
    16'b01101100_11010101 : OUT <= 0;  //108 / 213 = 0
    16'b01101100_11010110 : OUT <= 0;  //108 / 214 = 0
    16'b01101100_11010111 : OUT <= 0;  //108 / 215 = 0
    16'b01101100_11011000 : OUT <= 0;  //108 / 216 = 0
    16'b01101100_11011001 : OUT <= 0;  //108 / 217 = 0
    16'b01101100_11011010 : OUT <= 0;  //108 / 218 = 0
    16'b01101100_11011011 : OUT <= 0;  //108 / 219 = 0
    16'b01101100_11011100 : OUT <= 0;  //108 / 220 = 0
    16'b01101100_11011101 : OUT <= 0;  //108 / 221 = 0
    16'b01101100_11011110 : OUT <= 0;  //108 / 222 = 0
    16'b01101100_11011111 : OUT <= 0;  //108 / 223 = 0
    16'b01101100_11100000 : OUT <= 0;  //108 / 224 = 0
    16'b01101100_11100001 : OUT <= 0;  //108 / 225 = 0
    16'b01101100_11100010 : OUT <= 0;  //108 / 226 = 0
    16'b01101100_11100011 : OUT <= 0;  //108 / 227 = 0
    16'b01101100_11100100 : OUT <= 0;  //108 / 228 = 0
    16'b01101100_11100101 : OUT <= 0;  //108 / 229 = 0
    16'b01101100_11100110 : OUT <= 0;  //108 / 230 = 0
    16'b01101100_11100111 : OUT <= 0;  //108 / 231 = 0
    16'b01101100_11101000 : OUT <= 0;  //108 / 232 = 0
    16'b01101100_11101001 : OUT <= 0;  //108 / 233 = 0
    16'b01101100_11101010 : OUT <= 0;  //108 / 234 = 0
    16'b01101100_11101011 : OUT <= 0;  //108 / 235 = 0
    16'b01101100_11101100 : OUT <= 0;  //108 / 236 = 0
    16'b01101100_11101101 : OUT <= 0;  //108 / 237 = 0
    16'b01101100_11101110 : OUT <= 0;  //108 / 238 = 0
    16'b01101100_11101111 : OUT <= 0;  //108 / 239 = 0
    16'b01101100_11110000 : OUT <= 0;  //108 / 240 = 0
    16'b01101100_11110001 : OUT <= 0;  //108 / 241 = 0
    16'b01101100_11110010 : OUT <= 0;  //108 / 242 = 0
    16'b01101100_11110011 : OUT <= 0;  //108 / 243 = 0
    16'b01101100_11110100 : OUT <= 0;  //108 / 244 = 0
    16'b01101100_11110101 : OUT <= 0;  //108 / 245 = 0
    16'b01101100_11110110 : OUT <= 0;  //108 / 246 = 0
    16'b01101100_11110111 : OUT <= 0;  //108 / 247 = 0
    16'b01101100_11111000 : OUT <= 0;  //108 / 248 = 0
    16'b01101100_11111001 : OUT <= 0;  //108 / 249 = 0
    16'b01101100_11111010 : OUT <= 0;  //108 / 250 = 0
    16'b01101100_11111011 : OUT <= 0;  //108 / 251 = 0
    16'b01101100_11111100 : OUT <= 0;  //108 / 252 = 0
    16'b01101100_11111101 : OUT <= 0;  //108 / 253 = 0
    16'b01101100_11111110 : OUT <= 0;  //108 / 254 = 0
    16'b01101100_11111111 : OUT <= 0;  //108 / 255 = 0
    16'b01101101_00000000 : OUT <= 0;  //109 / 0 = 0
    16'b01101101_00000001 : OUT <= 109;  //109 / 1 = 109
    16'b01101101_00000010 : OUT <= 54;  //109 / 2 = 54
    16'b01101101_00000011 : OUT <= 36;  //109 / 3 = 36
    16'b01101101_00000100 : OUT <= 27;  //109 / 4 = 27
    16'b01101101_00000101 : OUT <= 21;  //109 / 5 = 21
    16'b01101101_00000110 : OUT <= 18;  //109 / 6 = 18
    16'b01101101_00000111 : OUT <= 15;  //109 / 7 = 15
    16'b01101101_00001000 : OUT <= 13;  //109 / 8 = 13
    16'b01101101_00001001 : OUT <= 12;  //109 / 9 = 12
    16'b01101101_00001010 : OUT <= 10;  //109 / 10 = 10
    16'b01101101_00001011 : OUT <= 9;  //109 / 11 = 9
    16'b01101101_00001100 : OUT <= 9;  //109 / 12 = 9
    16'b01101101_00001101 : OUT <= 8;  //109 / 13 = 8
    16'b01101101_00001110 : OUT <= 7;  //109 / 14 = 7
    16'b01101101_00001111 : OUT <= 7;  //109 / 15 = 7
    16'b01101101_00010000 : OUT <= 6;  //109 / 16 = 6
    16'b01101101_00010001 : OUT <= 6;  //109 / 17 = 6
    16'b01101101_00010010 : OUT <= 6;  //109 / 18 = 6
    16'b01101101_00010011 : OUT <= 5;  //109 / 19 = 5
    16'b01101101_00010100 : OUT <= 5;  //109 / 20 = 5
    16'b01101101_00010101 : OUT <= 5;  //109 / 21 = 5
    16'b01101101_00010110 : OUT <= 4;  //109 / 22 = 4
    16'b01101101_00010111 : OUT <= 4;  //109 / 23 = 4
    16'b01101101_00011000 : OUT <= 4;  //109 / 24 = 4
    16'b01101101_00011001 : OUT <= 4;  //109 / 25 = 4
    16'b01101101_00011010 : OUT <= 4;  //109 / 26 = 4
    16'b01101101_00011011 : OUT <= 4;  //109 / 27 = 4
    16'b01101101_00011100 : OUT <= 3;  //109 / 28 = 3
    16'b01101101_00011101 : OUT <= 3;  //109 / 29 = 3
    16'b01101101_00011110 : OUT <= 3;  //109 / 30 = 3
    16'b01101101_00011111 : OUT <= 3;  //109 / 31 = 3
    16'b01101101_00100000 : OUT <= 3;  //109 / 32 = 3
    16'b01101101_00100001 : OUT <= 3;  //109 / 33 = 3
    16'b01101101_00100010 : OUT <= 3;  //109 / 34 = 3
    16'b01101101_00100011 : OUT <= 3;  //109 / 35 = 3
    16'b01101101_00100100 : OUT <= 3;  //109 / 36 = 3
    16'b01101101_00100101 : OUT <= 2;  //109 / 37 = 2
    16'b01101101_00100110 : OUT <= 2;  //109 / 38 = 2
    16'b01101101_00100111 : OUT <= 2;  //109 / 39 = 2
    16'b01101101_00101000 : OUT <= 2;  //109 / 40 = 2
    16'b01101101_00101001 : OUT <= 2;  //109 / 41 = 2
    16'b01101101_00101010 : OUT <= 2;  //109 / 42 = 2
    16'b01101101_00101011 : OUT <= 2;  //109 / 43 = 2
    16'b01101101_00101100 : OUT <= 2;  //109 / 44 = 2
    16'b01101101_00101101 : OUT <= 2;  //109 / 45 = 2
    16'b01101101_00101110 : OUT <= 2;  //109 / 46 = 2
    16'b01101101_00101111 : OUT <= 2;  //109 / 47 = 2
    16'b01101101_00110000 : OUT <= 2;  //109 / 48 = 2
    16'b01101101_00110001 : OUT <= 2;  //109 / 49 = 2
    16'b01101101_00110010 : OUT <= 2;  //109 / 50 = 2
    16'b01101101_00110011 : OUT <= 2;  //109 / 51 = 2
    16'b01101101_00110100 : OUT <= 2;  //109 / 52 = 2
    16'b01101101_00110101 : OUT <= 2;  //109 / 53 = 2
    16'b01101101_00110110 : OUT <= 2;  //109 / 54 = 2
    16'b01101101_00110111 : OUT <= 1;  //109 / 55 = 1
    16'b01101101_00111000 : OUT <= 1;  //109 / 56 = 1
    16'b01101101_00111001 : OUT <= 1;  //109 / 57 = 1
    16'b01101101_00111010 : OUT <= 1;  //109 / 58 = 1
    16'b01101101_00111011 : OUT <= 1;  //109 / 59 = 1
    16'b01101101_00111100 : OUT <= 1;  //109 / 60 = 1
    16'b01101101_00111101 : OUT <= 1;  //109 / 61 = 1
    16'b01101101_00111110 : OUT <= 1;  //109 / 62 = 1
    16'b01101101_00111111 : OUT <= 1;  //109 / 63 = 1
    16'b01101101_01000000 : OUT <= 1;  //109 / 64 = 1
    16'b01101101_01000001 : OUT <= 1;  //109 / 65 = 1
    16'b01101101_01000010 : OUT <= 1;  //109 / 66 = 1
    16'b01101101_01000011 : OUT <= 1;  //109 / 67 = 1
    16'b01101101_01000100 : OUT <= 1;  //109 / 68 = 1
    16'b01101101_01000101 : OUT <= 1;  //109 / 69 = 1
    16'b01101101_01000110 : OUT <= 1;  //109 / 70 = 1
    16'b01101101_01000111 : OUT <= 1;  //109 / 71 = 1
    16'b01101101_01001000 : OUT <= 1;  //109 / 72 = 1
    16'b01101101_01001001 : OUT <= 1;  //109 / 73 = 1
    16'b01101101_01001010 : OUT <= 1;  //109 / 74 = 1
    16'b01101101_01001011 : OUT <= 1;  //109 / 75 = 1
    16'b01101101_01001100 : OUT <= 1;  //109 / 76 = 1
    16'b01101101_01001101 : OUT <= 1;  //109 / 77 = 1
    16'b01101101_01001110 : OUT <= 1;  //109 / 78 = 1
    16'b01101101_01001111 : OUT <= 1;  //109 / 79 = 1
    16'b01101101_01010000 : OUT <= 1;  //109 / 80 = 1
    16'b01101101_01010001 : OUT <= 1;  //109 / 81 = 1
    16'b01101101_01010010 : OUT <= 1;  //109 / 82 = 1
    16'b01101101_01010011 : OUT <= 1;  //109 / 83 = 1
    16'b01101101_01010100 : OUT <= 1;  //109 / 84 = 1
    16'b01101101_01010101 : OUT <= 1;  //109 / 85 = 1
    16'b01101101_01010110 : OUT <= 1;  //109 / 86 = 1
    16'b01101101_01010111 : OUT <= 1;  //109 / 87 = 1
    16'b01101101_01011000 : OUT <= 1;  //109 / 88 = 1
    16'b01101101_01011001 : OUT <= 1;  //109 / 89 = 1
    16'b01101101_01011010 : OUT <= 1;  //109 / 90 = 1
    16'b01101101_01011011 : OUT <= 1;  //109 / 91 = 1
    16'b01101101_01011100 : OUT <= 1;  //109 / 92 = 1
    16'b01101101_01011101 : OUT <= 1;  //109 / 93 = 1
    16'b01101101_01011110 : OUT <= 1;  //109 / 94 = 1
    16'b01101101_01011111 : OUT <= 1;  //109 / 95 = 1
    16'b01101101_01100000 : OUT <= 1;  //109 / 96 = 1
    16'b01101101_01100001 : OUT <= 1;  //109 / 97 = 1
    16'b01101101_01100010 : OUT <= 1;  //109 / 98 = 1
    16'b01101101_01100011 : OUT <= 1;  //109 / 99 = 1
    16'b01101101_01100100 : OUT <= 1;  //109 / 100 = 1
    16'b01101101_01100101 : OUT <= 1;  //109 / 101 = 1
    16'b01101101_01100110 : OUT <= 1;  //109 / 102 = 1
    16'b01101101_01100111 : OUT <= 1;  //109 / 103 = 1
    16'b01101101_01101000 : OUT <= 1;  //109 / 104 = 1
    16'b01101101_01101001 : OUT <= 1;  //109 / 105 = 1
    16'b01101101_01101010 : OUT <= 1;  //109 / 106 = 1
    16'b01101101_01101011 : OUT <= 1;  //109 / 107 = 1
    16'b01101101_01101100 : OUT <= 1;  //109 / 108 = 1
    16'b01101101_01101101 : OUT <= 1;  //109 / 109 = 1
    16'b01101101_01101110 : OUT <= 0;  //109 / 110 = 0
    16'b01101101_01101111 : OUT <= 0;  //109 / 111 = 0
    16'b01101101_01110000 : OUT <= 0;  //109 / 112 = 0
    16'b01101101_01110001 : OUT <= 0;  //109 / 113 = 0
    16'b01101101_01110010 : OUT <= 0;  //109 / 114 = 0
    16'b01101101_01110011 : OUT <= 0;  //109 / 115 = 0
    16'b01101101_01110100 : OUT <= 0;  //109 / 116 = 0
    16'b01101101_01110101 : OUT <= 0;  //109 / 117 = 0
    16'b01101101_01110110 : OUT <= 0;  //109 / 118 = 0
    16'b01101101_01110111 : OUT <= 0;  //109 / 119 = 0
    16'b01101101_01111000 : OUT <= 0;  //109 / 120 = 0
    16'b01101101_01111001 : OUT <= 0;  //109 / 121 = 0
    16'b01101101_01111010 : OUT <= 0;  //109 / 122 = 0
    16'b01101101_01111011 : OUT <= 0;  //109 / 123 = 0
    16'b01101101_01111100 : OUT <= 0;  //109 / 124 = 0
    16'b01101101_01111101 : OUT <= 0;  //109 / 125 = 0
    16'b01101101_01111110 : OUT <= 0;  //109 / 126 = 0
    16'b01101101_01111111 : OUT <= 0;  //109 / 127 = 0
    16'b01101101_10000000 : OUT <= 0;  //109 / 128 = 0
    16'b01101101_10000001 : OUT <= 0;  //109 / 129 = 0
    16'b01101101_10000010 : OUT <= 0;  //109 / 130 = 0
    16'b01101101_10000011 : OUT <= 0;  //109 / 131 = 0
    16'b01101101_10000100 : OUT <= 0;  //109 / 132 = 0
    16'b01101101_10000101 : OUT <= 0;  //109 / 133 = 0
    16'b01101101_10000110 : OUT <= 0;  //109 / 134 = 0
    16'b01101101_10000111 : OUT <= 0;  //109 / 135 = 0
    16'b01101101_10001000 : OUT <= 0;  //109 / 136 = 0
    16'b01101101_10001001 : OUT <= 0;  //109 / 137 = 0
    16'b01101101_10001010 : OUT <= 0;  //109 / 138 = 0
    16'b01101101_10001011 : OUT <= 0;  //109 / 139 = 0
    16'b01101101_10001100 : OUT <= 0;  //109 / 140 = 0
    16'b01101101_10001101 : OUT <= 0;  //109 / 141 = 0
    16'b01101101_10001110 : OUT <= 0;  //109 / 142 = 0
    16'b01101101_10001111 : OUT <= 0;  //109 / 143 = 0
    16'b01101101_10010000 : OUT <= 0;  //109 / 144 = 0
    16'b01101101_10010001 : OUT <= 0;  //109 / 145 = 0
    16'b01101101_10010010 : OUT <= 0;  //109 / 146 = 0
    16'b01101101_10010011 : OUT <= 0;  //109 / 147 = 0
    16'b01101101_10010100 : OUT <= 0;  //109 / 148 = 0
    16'b01101101_10010101 : OUT <= 0;  //109 / 149 = 0
    16'b01101101_10010110 : OUT <= 0;  //109 / 150 = 0
    16'b01101101_10010111 : OUT <= 0;  //109 / 151 = 0
    16'b01101101_10011000 : OUT <= 0;  //109 / 152 = 0
    16'b01101101_10011001 : OUT <= 0;  //109 / 153 = 0
    16'b01101101_10011010 : OUT <= 0;  //109 / 154 = 0
    16'b01101101_10011011 : OUT <= 0;  //109 / 155 = 0
    16'b01101101_10011100 : OUT <= 0;  //109 / 156 = 0
    16'b01101101_10011101 : OUT <= 0;  //109 / 157 = 0
    16'b01101101_10011110 : OUT <= 0;  //109 / 158 = 0
    16'b01101101_10011111 : OUT <= 0;  //109 / 159 = 0
    16'b01101101_10100000 : OUT <= 0;  //109 / 160 = 0
    16'b01101101_10100001 : OUT <= 0;  //109 / 161 = 0
    16'b01101101_10100010 : OUT <= 0;  //109 / 162 = 0
    16'b01101101_10100011 : OUT <= 0;  //109 / 163 = 0
    16'b01101101_10100100 : OUT <= 0;  //109 / 164 = 0
    16'b01101101_10100101 : OUT <= 0;  //109 / 165 = 0
    16'b01101101_10100110 : OUT <= 0;  //109 / 166 = 0
    16'b01101101_10100111 : OUT <= 0;  //109 / 167 = 0
    16'b01101101_10101000 : OUT <= 0;  //109 / 168 = 0
    16'b01101101_10101001 : OUT <= 0;  //109 / 169 = 0
    16'b01101101_10101010 : OUT <= 0;  //109 / 170 = 0
    16'b01101101_10101011 : OUT <= 0;  //109 / 171 = 0
    16'b01101101_10101100 : OUT <= 0;  //109 / 172 = 0
    16'b01101101_10101101 : OUT <= 0;  //109 / 173 = 0
    16'b01101101_10101110 : OUT <= 0;  //109 / 174 = 0
    16'b01101101_10101111 : OUT <= 0;  //109 / 175 = 0
    16'b01101101_10110000 : OUT <= 0;  //109 / 176 = 0
    16'b01101101_10110001 : OUT <= 0;  //109 / 177 = 0
    16'b01101101_10110010 : OUT <= 0;  //109 / 178 = 0
    16'b01101101_10110011 : OUT <= 0;  //109 / 179 = 0
    16'b01101101_10110100 : OUT <= 0;  //109 / 180 = 0
    16'b01101101_10110101 : OUT <= 0;  //109 / 181 = 0
    16'b01101101_10110110 : OUT <= 0;  //109 / 182 = 0
    16'b01101101_10110111 : OUT <= 0;  //109 / 183 = 0
    16'b01101101_10111000 : OUT <= 0;  //109 / 184 = 0
    16'b01101101_10111001 : OUT <= 0;  //109 / 185 = 0
    16'b01101101_10111010 : OUT <= 0;  //109 / 186 = 0
    16'b01101101_10111011 : OUT <= 0;  //109 / 187 = 0
    16'b01101101_10111100 : OUT <= 0;  //109 / 188 = 0
    16'b01101101_10111101 : OUT <= 0;  //109 / 189 = 0
    16'b01101101_10111110 : OUT <= 0;  //109 / 190 = 0
    16'b01101101_10111111 : OUT <= 0;  //109 / 191 = 0
    16'b01101101_11000000 : OUT <= 0;  //109 / 192 = 0
    16'b01101101_11000001 : OUT <= 0;  //109 / 193 = 0
    16'b01101101_11000010 : OUT <= 0;  //109 / 194 = 0
    16'b01101101_11000011 : OUT <= 0;  //109 / 195 = 0
    16'b01101101_11000100 : OUT <= 0;  //109 / 196 = 0
    16'b01101101_11000101 : OUT <= 0;  //109 / 197 = 0
    16'b01101101_11000110 : OUT <= 0;  //109 / 198 = 0
    16'b01101101_11000111 : OUT <= 0;  //109 / 199 = 0
    16'b01101101_11001000 : OUT <= 0;  //109 / 200 = 0
    16'b01101101_11001001 : OUT <= 0;  //109 / 201 = 0
    16'b01101101_11001010 : OUT <= 0;  //109 / 202 = 0
    16'b01101101_11001011 : OUT <= 0;  //109 / 203 = 0
    16'b01101101_11001100 : OUT <= 0;  //109 / 204 = 0
    16'b01101101_11001101 : OUT <= 0;  //109 / 205 = 0
    16'b01101101_11001110 : OUT <= 0;  //109 / 206 = 0
    16'b01101101_11001111 : OUT <= 0;  //109 / 207 = 0
    16'b01101101_11010000 : OUT <= 0;  //109 / 208 = 0
    16'b01101101_11010001 : OUT <= 0;  //109 / 209 = 0
    16'b01101101_11010010 : OUT <= 0;  //109 / 210 = 0
    16'b01101101_11010011 : OUT <= 0;  //109 / 211 = 0
    16'b01101101_11010100 : OUT <= 0;  //109 / 212 = 0
    16'b01101101_11010101 : OUT <= 0;  //109 / 213 = 0
    16'b01101101_11010110 : OUT <= 0;  //109 / 214 = 0
    16'b01101101_11010111 : OUT <= 0;  //109 / 215 = 0
    16'b01101101_11011000 : OUT <= 0;  //109 / 216 = 0
    16'b01101101_11011001 : OUT <= 0;  //109 / 217 = 0
    16'b01101101_11011010 : OUT <= 0;  //109 / 218 = 0
    16'b01101101_11011011 : OUT <= 0;  //109 / 219 = 0
    16'b01101101_11011100 : OUT <= 0;  //109 / 220 = 0
    16'b01101101_11011101 : OUT <= 0;  //109 / 221 = 0
    16'b01101101_11011110 : OUT <= 0;  //109 / 222 = 0
    16'b01101101_11011111 : OUT <= 0;  //109 / 223 = 0
    16'b01101101_11100000 : OUT <= 0;  //109 / 224 = 0
    16'b01101101_11100001 : OUT <= 0;  //109 / 225 = 0
    16'b01101101_11100010 : OUT <= 0;  //109 / 226 = 0
    16'b01101101_11100011 : OUT <= 0;  //109 / 227 = 0
    16'b01101101_11100100 : OUT <= 0;  //109 / 228 = 0
    16'b01101101_11100101 : OUT <= 0;  //109 / 229 = 0
    16'b01101101_11100110 : OUT <= 0;  //109 / 230 = 0
    16'b01101101_11100111 : OUT <= 0;  //109 / 231 = 0
    16'b01101101_11101000 : OUT <= 0;  //109 / 232 = 0
    16'b01101101_11101001 : OUT <= 0;  //109 / 233 = 0
    16'b01101101_11101010 : OUT <= 0;  //109 / 234 = 0
    16'b01101101_11101011 : OUT <= 0;  //109 / 235 = 0
    16'b01101101_11101100 : OUT <= 0;  //109 / 236 = 0
    16'b01101101_11101101 : OUT <= 0;  //109 / 237 = 0
    16'b01101101_11101110 : OUT <= 0;  //109 / 238 = 0
    16'b01101101_11101111 : OUT <= 0;  //109 / 239 = 0
    16'b01101101_11110000 : OUT <= 0;  //109 / 240 = 0
    16'b01101101_11110001 : OUT <= 0;  //109 / 241 = 0
    16'b01101101_11110010 : OUT <= 0;  //109 / 242 = 0
    16'b01101101_11110011 : OUT <= 0;  //109 / 243 = 0
    16'b01101101_11110100 : OUT <= 0;  //109 / 244 = 0
    16'b01101101_11110101 : OUT <= 0;  //109 / 245 = 0
    16'b01101101_11110110 : OUT <= 0;  //109 / 246 = 0
    16'b01101101_11110111 : OUT <= 0;  //109 / 247 = 0
    16'b01101101_11111000 : OUT <= 0;  //109 / 248 = 0
    16'b01101101_11111001 : OUT <= 0;  //109 / 249 = 0
    16'b01101101_11111010 : OUT <= 0;  //109 / 250 = 0
    16'b01101101_11111011 : OUT <= 0;  //109 / 251 = 0
    16'b01101101_11111100 : OUT <= 0;  //109 / 252 = 0
    16'b01101101_11111101 : OUT <= 0;  //109 / 253 = 0
    16'b01101101_11111110 : OUT <= 0;  //109 / 254 = 0
    16'b01101101_11111111 : OUT <= 0;  //109 / 255 = 0
    16'b01101110_00000000 : OUT <= 0;  //110 / 0 = 0
    16'b01101110_00000001 : OUT <= 110;  //110 / 1 = 110
    16'b01101110_00000010 : OUT <= 55;  //110 / 2 = 55
    16'b01101110_00000011 : OUT <= 36;  //110 / 3 = 36
    16'b01101110_00000100 : OUT <= 27;  //110 / 4 = 27
    16'b01101110_00000101 : OUT <= 22;  //110 / 5 = 22
    16'b01101110_00000110 : OUT <= 18;  //110 / 6 = 18
    16'b01101110_00000111 : OUT <= 15;  //110 / 7 = 15
    16'b01101110_00001000 : OUT <= 13;  //110 / 8 = 13
    16'b01101110_00001001 : OUT <= 12;  //110 / 9 = 12
    16'b01101110_00001010 : OUT <= 11;  //110 / 10 = 11
    16'b01101110_00001011 : OUT <= 10;  //110 / 11 = 10
    16'b01101110_00001100 : OUT <= 9;  //110 / 12 = 9
    16'b01101110_00001101 : OUT <= 8;  //110 / 13 = 8
    16'b01101110_00001110 : OUT <= 7;  //110 / 14 = 7
    16'b01101110_00001111 : OUT <= 7;  //110 / 15 = 7
    16'b01101110_00010000 : OUT <= 6;  //110 / 16 = 6
    16'b01101110_00010001 : OUT <= 6;  //110 / 17 = 6
    16'b01101110_00010010 : OUT <= 6;  //110 / 18 = 6
    16'b01101110_00010011 : OUT <= 5;  //110 / 19 = 5
    16'b01101110_00010100 : OUT <= 5;  //110 / 20 = 5
    16'b01101110_00010101 : OUT <= 5;  //110 / 21 = 5
    16'b01101110_00010110 : OUT <= 5;  //110 / 22 = 5
    16'b01101110_00010111 : OUT <= 4;  //110 / 23 = 4
    16'b01101110_00011000 : OUT <= 4;  //110 / 24 = 4
    16'b01101110_00011001 : OUT <= 4;  //110 / 25 = 4
    16'b01101110_00011010 : OUT <= 4;  //110 / 26 = 4
    16'b01101110_00011011 : OUT <= 4;  //110 / 27 = 4
    16'b01101110_00011100 : OUT <= 3;  //110 / 28 = 3
    16'b01101110_00011101 : OUT <= 3;  //110 / 29 = 3
    16'b01101110_00011110 : OUT <= 3;  //110 / 30 = 3
    16'b01101110_00011111 : OUT <= 3;  //110 / 31 = 3
    16'b01101110_00100000 : OUT <= 3;  //110 / 32 = 3
    16'b01101110_00100001 : OUT <= 3;  //110 / 33 = 3
    16'b01101110_00100010 : OUT <= 3;  //110 / 34 = 3
    16'b01101110_00100011 : OUT <= 3;  //110 / 35 = 3
    16'b01101110_00100100 : OUT <= 3;  //110 / 36 = 3
    16'b01101110_00100101 : OUT <= 2;  //110 / 37 = 2
    16'b01101110_00100110 : OUT <= 2;  //110 / 38 = 2
    16'b01101110_00100111 : OUT <= 2;  //110 / 39 = 2
    16'b01101110_00101000 : OUT <= 2;  //110 / 40 = 2
    16'b01101110_00101001 : OUT <= 2;  //110 / 41 = 2
    16'b01101110_00101010 : OUT <= 2;  //110 / 42 = 2
    16'b01101110_00101011 : OUT <= 2;  //110 / 43 = 2
    16'b01101110_00101100 : OUT <= 2;  //110 / 44 = 2
    16'b01101110_00101101 : OUT <= 2;  //110 / 45 = 2
    16'b01101110_00101110 : OUT <= 2;  //110 / 46 = 2
    16'b01101110_00101111 : OUT <= 2;  //110 / 47 = 2
    16'b01101110_00110000 : OUT <= 2;  //110 / 48 = 2
    16'b01101110_00110001 : OUT <= 2;  //110 / 49 = 2
    16'b01101110_00110010 : OUT <= 2;  //110 / 50 = 2
    16'b01101110_00110011 : OUT <= 2;  //110 / 51 = 2
    16'b01101110_00110100 : OUT <= 2;  //110 / 52 = 2
    16'b01101110_00110101 : OUT <= 2;  //110 / 53 = 2
    16'b01101110_00110110 : OUT <= 2;  //110 / 54 = 2
    16'b01101110_00110111 : OUT <= 2;  //110 / 55 = 2
    16'b01101110_00111000 : OUT <= 1;  //110 / 56 = 1
    16'b01101110_00111001 : OUT <= 1;  //110 / 57 = 1
    16'b01101110_00111010 : OUT <= 1;  //110 / 58 = 1
    16'b01101110_00111011 : OUT <= 1;  //110 / 59 = 1
    16'b01101110_00111100 : OUT <= 1;  //110 / 60 = 1
    16'b01101110_00111101 : OUT <= 1;  //110 / 61 = 1
    16'b01101110_00111110 : OUT <= 1;  //110 / 62 = 1
    16'b01101110_00111111 : OUT <= 1;  //110 / 63 = 1
    16'b01101110_01000000 : OUT <= 1;  //110 / 64 = 1
    16'b01101110_01000001 : OUT <= 1;  //110 / 65 = 1
    16'b01101110_01000010 : OUT <= 1;  //110 / 66 = 1
    16'b01101110_01000011 : OUT <= 1;  //110 / 67 = 1
    16'b01101110_01000100 : OUT <= 1;  //110 / 68 = 1
    16'b01101110_01000101 : OUT <= 1;  //110 / 69 = 1
    16'b01101110_01000110 : OUT <= 1;  //110 / 70 = 1
    16'b01101110_01000111 : OUT <= 1;  //110 / 71 = 1
    16'b01101110_01001000 : OUT <= 1;  //110 / 72 = 1
    16'b01101110_01001001 : OUT <= 1;  //110 / 73 = 1
    16'b01101110_01001010 : OUT <= 1;  //110 / 74 = 1
    16'b01101110_01001011 : OUT <= 1;  //110 / 75 = 1
    16'b01101110_01001100 : OUT <= 1;  //110 / 76 = 1
    16'b01101110_01001101 : OUT <= 1;  //110 / 77 = 1
    16'b01101110_01001110 : OUT <= 1;  //110 / 78 = 1
    16'b01101110_01001111 : OUT <= 1;  //110 / 79 = 1
    16'b01101110_01010000 : OUT <= 1;  //110 / 80 = 1
    16'b01101110_01010001 : OUT <= 1;  //110 / 81 = 1
    16'b01101110_01010010 : OUT <= 1;  //110 / 82 = 1
    16'b01101110_01010011 : OUT <= 1;  //110 / 83 = 1
    16'b01101110_01010100 : OUT <= 1;  //110 / 84 = 1
    16'b01101110_01010101 : OUT <= 1;  //110 / 85 = 1
    16'b01101110_01010110 : OUT <= 1;  //110 / 86 = 1
    16'b01101110_01010111 : OUT <= 1;  //110 / 87 = 1
    16'b01101110_01011000 : OUT <= 1;  //110 / 88 = 1
    16'b01101110_01011001 : OUT <= 1;  //110 / 89 = 1
    16'b01101110_01011010 : OUT <= 1;  //110 / 90 = 1
    16'b01101110_01011011 : OUT <= 1;  //110 / 91 = 1
    16'b01101110_01011100 : OUT <= 1;  //110 / 92 = 1
    16'b01101110_01011101 : OUT <= 1;  //110 / 93 = 1
    16'b01101110_01011110 : OUT <= 1;  //110 / 94 = 1
    16'b01101110_01011111 : OUT <= 1;  //110 / 95 = 1
    16'b01101110_01100000 : OUT <= 1;  //110 / 96 = 1
    16'b01101110_01100001 : OUT <= 1;  //110 / 97 = 1
    16'b01101110_01100010 : OUT <= 1;  //110 / 98 = 1
    16'b01101110_01100011 : OUT <= 1;  //110 / 99 = 1
    16'b01101110_01100100 : OUT <= 1;  //110 / 100 = 1
    16'b01101110_01100101 : OUT <= 1;  //110 / 101 = 1
    16'b01101110_01100110 : OUT <= 1;  //110 / 102 = 1
    16'b01101110_01100111 : OUT <= 1;  //110 / 103 = 1
    16'b01101110_01101000 : OUT <= 1;  //110 / 104 = 1
    16'b01101110_01101001 : OUT <= 1;  //110 / 105 = 1
    16'b01101110_01101010 : OUT <= 1;  //110 / 106 = 1
    16'b01101110_01101011 : OUT <= 1;  //110 / 107 = 1
    16'b01101110_01101100 : OUT <= 1;  //110 / 108 = 1
    16'b01101110_01101101 : OUT <= 1;  //110 / 109 = 1
    16'b01101110_01101110 : OUT <= 1;  //110 / 110 = 1
    16'b01101110_01101111 : OUT <= 0;  //110 / 111 = 0
    16'b01101110_01110000 : OUT <= 0;  //110 / 112 = 0
    16'b01101110_01110001 : OUT <= 0;  //110 / 113 = 0
    16'b01101110_01110010 : OUT <= 0;  //110 / 114 = 0
    16'b01101110_01110011 : OUT <= 0;  //110 / 115 = 0
    16'b01101110_01110100 : OUT <= 0;  //110 / 116 = 0
    16'b01101110_01110101 : OUT <= 0;  //110 / 117 = 0
    16'b01101110_01110110 : OUT <= 0;  //110 / 118 = 0
    16'b01101110_01110111 : OUT <= 0;  //110 / 119 = 0
    16'b01101110_01111000 : OUT <= 0;  //110 / 120 = 0
    16'b01101110_01111001 : OUT <= 0;  //110 / 121 = 0
    16'b01101110_01111010 : OUT <= 0;  //110 / 122 = 0
    16'b01101110_01111011 : OUT <= 0;  //110 / 123 = 0
    16'b01101110_01111100 : OUT <= 0;  //110 / 124 = 0
    16'b01101110_01111101 : OUT <= 0;  //110 / 125 = 0
    16'b01101110_01111110 : OUT <= 0;  //110 / 126 = 0
    16'b01101110_01111111 : OUT <= 0;  //110 / 127 = 0
    16'b01101110_10000000 : OUT <= 0;  //110 / 128 = 0
    16'b01101110_10000001 : OUT <= 0;  //110 / 129 = 0
    16'b01101110_10000010 : OUT <= 0;  //110 / 130 = 0
    16'b01101110_10000011 : OUT <= 0;  //110 / 131 = 0
    16'b01101110_10000100 : OUT <= 0;  //110 / 132 = 0
    16'b01101110_10000101 : OUT <= 0;  //110 / 133 = 0
    16'b01101110_10000110 : OUT <= 0;  //110 / 134 = 0
    16'b01101110_10000111 : OUT <= 0;  //110 / 135 = 0
    16'b01101110_10001000 : OUT <= 0;  //110 / 136 = 0
    16'b01101110_10001001 : OUT <= 0;  //110 / 137 = 0
    16'b01101110_10001010 : OUT <= 0;  //110 / 138 = 0
    16'b01101110_10001011 : OUT <= 0;  //110 / 139 = 0
    16'b01101110_10001100 : OUT <= 0;  //110 / 140 = 0
    16'b01101110_10001101 : OUT <= 0;  //110 / 141 = 0
    16'b01101110_10001110 : OUT <= 0;  //110 / 142 = 0
    16'b01101110_10001111 : OUT <= 0;  //110 / 143 = 0
    16'b01101110_10010000 : OUT <= 0;  //110 / 144 = 0
    16'b01101110_10010001 : OUT <= 0;  //110 / 145 = 0
    16'b01101110_10010010 : OUT <= 0;  //110 / 146 = 0
    16'b01101110_10010011 : OUT <= 0;  //110 / 147 = 0
    16'b01101110_10010100 : OUT <= 0;  //110 / 148 = 0
    16'b01101110_10010101 : OUT <= 0;  //110 / 149 = 0
    16'b01101110_10010110 : OUT <= 0;  //110 / 150 = 0
    16'b01101110_10010111 : OUT <= 0;  //110 / 151 = 0
    16'b01101110_10011000 : OUT <= 0;  //110 / 152 = 0
    16'b01101110_10011001 : OUT <= 0;  //110 / 153 = 0
    16'b01101110_10011010 : OUT <= 0;  //110 / 154 = 0
    16'b01101110_10011011 : OUT <= 0;  //110 / 155 = 0
    16'b01101110_10011100 : OUT <= 0;  //110 / 156 = 0
    16'b01101110_10011101 : OUT <= 0;  //110 / 157 = 0
    16'b01101110_10011110 : OUT <= 0;  //110 / 158 = 0
    16'b01101110_10011111 : OUT <= 0;  //110 / 159 = 0
    16'b01101110_10100000 : OUT <= 0;  //110 / 160 = 0
    16'b01101110_10100001 : OUT <= 0;  //110 / 161 = 0
    16'b01101110_10100010 : OUT <= 0;  //110 / 162 = 0
    16'b01101110_10100011 : OUT <= 0;  //110 / 163 = 0
    16'b01101110_10100100 : OUT <= 0;  //110 / 164 = 0
    16'b01101110_10100101 : OUT <= 0;  //110 / 165 = 0
    16'b01101110_10100110 : OUT <= 0;  //110 / 166 = 0
    16'b01101110_10100111 : OUT <= 0;  //110 / 167 = 0
    16'b01101110_10101000 : OUT <= 0;  //110 / 168 = 0
    16'b01101110_10101001 : OUT <= 0;  //110 / 169 = 0
    16'b01101110_10101010 : OUT <= 0;  //110 / 170 = 0
    16'b01101110_10101011 : OUT <= 0;  //110 / 171 = 0
    16'b01101110_10101100 : OUT <= 0;  //110 / 172 = 0
    16'b01101110_10101101 : OUT <= 0;  //110 / 173 = 0
    16'b01101110_10101110 : OUT <= 0;  //110 / 174 = 0
    16'b01101110_10101111 : OUT <= 0;  //110 / 175 = 0
    16'b01101110_10110000 : OUT <= 0;  //110 / 176 = 0
    16'b01101110_10110001 : OUT <= 0;  //110 / 177 = 0
    16'b01101110_10110010 : OUT <= 0;  //110 / 178 = 0
    16'b01101110_10110011 : OUT <= 0;  //110 / 179 = 0
    16'b01101110_10110100 : OUT <= 0;  //110 / 180 = 0
    16'b01101110_10110101 : OUT <= 0;  //110 / 181 = 0
    16'b01101110_10110110 : OUT <= 0;  //110 / 182 = 0
    16'b01101110_10110111 : OUT <= 0;  //110 / 183 = 0
    16'b01101110_10111000 : OUT <= 0;  //110 / 184 = 0
    16'b01101110_10111001 : OUT <= 0;  //110 / 185 = 0
    16'b01101110_10111010 : OUT <= 0;  //110 / 186 = 0
    16'b01101110_10111011 : OUT <= 0;  //110 / 187 = 0
    16'b01101110_10111100 : OUT <= 0;  //110 / 188 = 0
    16'b01101110_10111101 : OUT <= 0;  //110 / 189 = 0
    16'b01101110_10111110 : OUT <= 0;  //110 / 190 = 0
    16'b01101110_10111111 : OUT <= 0;  //110 / 191 = 0
    16'b01101110_11000000 : OUT <= 0;  //110 / 192 = 0
    16'b01101110_11000001 : OUT <= 0;  //110 / 193 = 0
    16'b01101110_11000010 : OUT <= 0;  //110 / 194 = 0
    16'b01101110_11000011 : OUT <= 0;  //110 / 195 = 0
    16'b01101110_11000100 : OUT <= 0;  //110 / 196 = 0
    16'b01101110_11000101 : OUT <= 0;  //110 / 197 = 0
    16'b01101110_11000110 : OUT <= 0;  //110 / 198 = 0
    16'b01101110_11000111 : OUT <= 0;  //110 / 199 = 0
    16'b01101110_11001000 : OUT <= 0;  //110 / 200 = 0
    16'b01101110_11001001 : OUT <= 0;  //110 / 201 = 0
    16'b01101110_11001010 : OUT <= 0;  //110 / 202 = 0
    16'b01101110_11001011 : OUT <= 0;  //110 / 203 = 0
    16'b01101110_11001100 : OUT <= 0;  //110 / 204 = 0
    16'b01101110_11001101 : OUT <= 0;  //110 / 205 = 0
    16'b01101110_11001110 : OUT <= 0;  //110 / 206 = 0
    16'b01101110_11001111 : OUT <= 0;  //110 / 207 = 0
    16'b01101110_11010000 : OUT <= 0;  //110 / 208 = 0
    16'b01101110_11010001 : OUT <= 0;  //110 / 209 = 0
    16'b01101110_11010010 : OUT <= 0;  //110 / 210 = 0
    16'b01101110_11010011 : OUT <= 0;  //110 / 211 = 0
    16'b01101110_11010100 : OUT <= 0;  //110 / 212 = 0
    16'b01101110_11010101 : OUT <= 0;  //110 / 213 = 0
    16'b01101110_11010110 : OUT <= 0;  //110 / 214 = 0
    16'b01101110_11010111 : OUT <= 0;  //110 / 215 = 0
    16'b01101110_11011000 : OUT <= 0;  //110 / 216 = 0
    16'b01101110_11011001 : OUT <= 0;  //110 / 217 = 0
    16'b01101110_11011010 : OUT <= 0;  //110 / 218 = 0
    16'b01101110_11011011 : OUT <= 0;  //110 / 219 = 0
    16'b01101110_11011100 : OUT <= 0;  //110 / 220 = 0
    16'b01101110_11011101 : OUT <= 0;  //110 / 221 = 0
    16'b01101110_11011110 : OUT <= 0;  //110 / 222 = 0
    16'b01101110_11011111 : OUT <= 0;  //110 / 223 = 0
    16'b01101110_11100000 : OUT <= 0;  //110 / 224 = 0
    16'b01101110_11100001 : OUT <= 0;  //110 / 225 = 0
    16'b01101110_11100010 : OUT <= 0;  //110 / 226 = 0
    16'b01101110_11100011 : OUT <= 0;  //110 / 227 = 0
    16'b01101110_11100100 : OUT <= 0;  //110 / 228 = 0
    16'b01101110_11100101 : OUT <= 0;  //110 / 229 = 0
    16'b01101110_11100110 : OUT <= 0;  //110 / 230 = 0
    16'b01101110_11100111 : OUT <= 0;  //110 / 231 = 0
    16'b01101110_11101000 : OUT <= 0;  //110 / 232 = 0
    16'b01101110_11101001 : OUT <= 0;  //110 / 233 = 0
    16'b01101110_11101010 : OUT <= 0;  //110 / 234 = 0
    16'b01101110_11101011 : OUT <= 0;  //110 / 235 = 0
    16'b01101110_11101100 : OUT <= 0;  //110 / 236 = 0
    16'b01101110_11101101 : OUT <= 0;  //110 / 237 = 0
    16'b01101110_11101110 : OUT <= 0;  //110 / 238 = 0
    16'b01101110_11101111 : OUT <= 0;  //110 / 239 = 0
    16'b01101110_11110000 : OUT <= 0;  //110 / 240 = 0
    16'b01101110_11110001 : OUT <= 0;  //110 / 241 = 0
    16'b01101110_11110010 : OUT <= 0;  //110 / 242 = 0
    16'b01101110_11110011 : OUT <= 0;  //110 / 243 = 0
    16'b01101110_11110100 : OUT <= 0;  //110 / 244 = 0
    16'b01101110_11110101 : OUT <= 0;  //110 / 245 = 0
    16'b01101110_11110110 : OUT <= 0;  //110 / 246 = 0
    16'b01101110_11110111 : OUT <= 0;  //110 / 247 = 0
    16'b01101110_11111000 : OUT <= 0;  //110 / 248 = 0
    16'b01101110_11111001 : OUT <= 0;  //110 / 249 = 0
    16'b01101110_11111010 : OUT <= 0;  //110 / 250 = 0
    16'b01101110_11111011 : OUT <= 0;  //110 / 251 = 0
    16'b01101110_11111100 : OUT <= 0;  //110 / 252 = 0
    16'b01101110_11111101 : OUT <= 0;  //110 / 253 = 0
    16'b01101110_11111110 : OUT <= 0;  //110 / 254 = 0
    16'b01101110_11111111 : OUT <= 0;  //110 / 255 = 0
    16'b01101111_00000000 : OUT <= 0;  //111 / 0 = 0
    16'b01101111_00000001 : OUT <= 111;  //111 / 1 = 111
    16'b01101111_00000010 : OUT <= 55;  //111 / 2 = 55
    16'b01101111_00000011 : OUT <= 37;  //111 / 3 = 37
    16'b01101111_00000100 : OUT <= 27;  //111 / 4 = 27
    16'b01101111_00000101 : OUT <= 22;  //111 / 5 = 22
    16'b01101111_00000110 : OUT <= 18;  //111 / 6 = 18
    16'b01101111_00000111 : OUT <= 15;  //111 / 7 = 15
    16'b01101111_00001000 : OUT <= 13;  //111 / 8 = 13
    16'b01101111_00001001 : OUT <= 12;  //111 / 9 = 12
    16'b01101111_00001010 : OUT <= 11;  //111 / 10 = 11
    16'b01101111_00001011 : OUT <= 10;  //111 / 11 = 10
    16'b01101111_00001100 : OUT <= 9;  //111 / 12 = 9
    16'b01101111_00001101 : OUT <= 8;  //111 / 13 = 8
    16'b01101111_00001110 : OUT <= 7;  //111 / 14 = 7
    16'b01101111_00001111 : OUT <= 7;  //111 / 15 = 7
    16'b01101111_00010000 : OUT <= 6;  //111 / 16 = 6
    16'b01101111_00010001 : OUT <= 6;  //111 / 17 = 6
    16'b01101111_00010010 : OUT <= 6;  //111 / 18 = 6
    16'b01101111_00010011 : OUT <= 5;  //111 / 19 = 5
    16'b01101111_00010100 : OUT <= 5;  //111 / 20 = 5
    16'b01101111_00010101 : OUT <= 5;  //111 / 21 = 5
    16'b01101111_00010110 : OUT <= 5;  //111 / 22 = 5
    16'b01101111_00010111 : OUT <= 4;  //111 / 23 = 4
    16'b01101111_00011000 : OUT <= 4;  //111 / 24 = 4
    16'b01101111_00011001 : OUT <= 4;  //111 / 25 = 4
    16'b01101111_00011010 : OUT <= 4;  //111 / 26 = 4
    16'b01101111_00011011 : OUT <= 4;  //111 / 27 = 4
    16'b01101111_00011100 : OUT <= 3;  //111 / 28 = 3
    16'b01101111_00011101 : OUT <= 3;  //111 / 29 = 3
    16'b01101111_00011110 : OUT <= 3;  //111 / 30 = 3
    16'b01101111_00011111 : OUT <= 3;  //111 / 31 = 3
    16'b01101111_00100000 : OUT <= 3;  //111 / 32 = 3
    16'b01101111_00100001 : OUT <= 3;  //111 / 33 = 3
    16'b01101111_00100010 : OUT <= 3;  //111 / 34 = 3
    16'b01101111_00100011 : OUT <= 3;  //111 / 35 = 3
    16'b01101111_00100100 : OUT <= 3;  //111 / 36 = 3
    16'b01101111_00100101 : OUT <= 3;  //111 / 37 = 3
    16'b01101111_00100110 : OUT <= 2;  //111 / 38 = 2
    16'b01101111_00100111 : OUT <= 2;  //111 / 39 = 2
    16'b01101111_00101000 : OUT <= 2;  //111 / 40 = 2
    16'b01101111_00101001 : OUT <= 2;  //111 / 41 = 2
    16'b01101111_00101010 : OUT <= 2;  //111 / 42 = 2
    16'b01101111_00101011 : OUT <= 2;  //111 / 43 = 2
    16'b01101111_00101100 : OUT <= 2;  //111 / 44 = 2
    16'b01101111_00101101 : OUT <= 2;  //111 / 45 = 2
    16'b01101111_00101110 : OUT <= 2;  //111 / 46 = 2
    16'b01101111_00101111 : OUT <= 2;  //111 / 47 = 2
    16'b01101111_00110000 : OUT <= 2;  //111 / 48 = 2
    16'b01101111_00110001 : OUT <= 2;  //111 / 49 = 2
    16'b01101111_00110010 : OUT <= 2;  //111 / 50 = 2
    16'b01101111_00110011 : OUT <= 2;  //111 / 51 = 2
    16'b01101111_00110100 : OUT <= 2;  //111 / 52 = 2
    16'b01101111_00110101 : OUT <= 2;  //111 / 53 = 2
    16'b01101111_00110110 : OUT <= 2;  //111 / 54 = 2
    16'b01101111_00110111 : OUT <= 2;  //111 / 55 = 2
    16'b01101111_00111000 : OUT <= 1;  //111 / 56 = 1
    16'b01101111_00111001 : OUT <= 1;  //111 / 57 = 1
    16'b01101111_00111010 : OUT <= 1;  //111 / 58 = 1
    16'b01101111_00111011 : OUT <= 1;  //111 / 59 = 1
    16'b01101111_00111100 : OUT <= 1;  //111 / 60 = 1
    16'b01101111_00111101 : OUT <= 1;  //111 / 61 = 1
    16'b01101111_00111110 : OUT <= 1;  //111 / 62 = 1
    16'b01101111_00111111 : OUT <= 1;  //111 / 63 = 1
    16'b01101111_01000000 : OUT <= 1;  //111 / 64 = 1
    16'b01101111_01000001 : OUT <= 1;  //111 / 65 = 1
    16'b01101111_01000010 : OUT <= 1;  //111 / 66 = 1
    16'b01101111_01000011 : OUT <= 1;  //111 / 67 = 1
    16'b01101111_01000100 : OUT <= 1;  //111 / 68 = 1
    16'b01101111_01000101 : OUT <= 1;  //111 / 69 = 1
    16'b01101111_01000110 : OUT <= 1;  //111 / 70 = 1
    16'b01101111_01000111 : OUT <= 1;  //111 / 71 = 1
    16'b01101111_01001000 : OUT <= 1;  //111 / 72 = 1
    16'b01101111_01001001 : OUT <= 1;  //111 / 73 = 1
    16'b01101111_01001010 : OUT <= 1;  //111 / 74 = 1
    16'b01101111_01001011 : OUT <= 1;  //111 / 75 = 1
    16'b01101111_01001100 : OUT <= 1;  //111 / 76 = 1
    16'b01101111_01001101 : OUT <= 1;  //111 / 77 = 1
    16'b01101111_01001110 : OUT <= 1;  //111 / 78 = 1
    16'b01101111_01001111 : OUT <= 1;  //111 / 79 = 1
    16'b01101111_01010000 : OUT <= 1;  //111 / 80 = 1
    16'b01101111_01010001 : OUT <= 1;  //111 / 81 = 1
    16'b01101111_01010010 : OUT <= 1;  //111 / 82 = 1
    16'b01101111_01010011 : OUT <= 1;  //111 / 83 = 1
    16'b01101111_01010100 : OUT <= 1;  //111 / 84 = 1
    16'b01101111_01010101 : OUT <= 1;  //111 / 85 = 1
    16'b01101111_01010110 : OUT <= 1;  //111 / 86 = 1
    16'b01101111_01010111 : OUT <= 1;  //111 / 87 = 1
    16'b01101111_01011000 : OUT <= 1;  //111 / 88 = 1
    16'b01101111_01011001 : OUT <= 1;  //111 / 89 = 1
    16'b01101111_01011010 : OUT <= 1;  //111 / 90 = 1
    16'b01101111_01011011 : OUT <= 1;  //111 / 91 = 1
    16'b01101111_01011100 : OUT <= 1;  //111 / 92 = 1
    16'b01101111_01011101 : OUT <= 1;  //111 / 93 = 1
    16'b01101111_01011110 : OUT <= 1;  //111 / 94 = 1
    16'b01101111_01011111 : OUT <= 1;  //111 / 95 = 1
    16'b01101111_01100000 : OUT <= 1;  //111 / 96 = 1
    16'b01101111_01100001 : OUT <= 1;  //111 / 97 = 1
    16'b01101111_01100010 : OUT <= 1;  //111 / 98 = 1
    16'b01101111_01100011 : OUT <= 1;  //111 / 99 = 1
    16'b01101111_01100100 : OUT <= 1;  //111 / 100 = 1
    16'b01101111_01100101 : OUT <= 1;  //111 / 101 = 1
    16'b01101111_01100110 : OUT <= 1;  //111 / 102 = 1
    16'b01101111_01100111 : OUT <= 1;  //111 / 103 = 1
    16'b01101111_01101000 : OUT <= 1;  //111 / 104 = 1
    16'b01101111_01101001 : OUT <= 1;  //111 / 105 = 1
    16'b01101111_01101010 : OUT <= 1;  //111 / 106 = 1
    16'b01101111_01101011 : OUT <= 1;  //111 / 107 = 1
    16'b01101111_01101100 : OUT <= 1;  //111 / 108 = 1
    16'b01101111_01101101 : OUT <= 1;  //111 / 109 = 1
    16'b01101111_01101110 : OUT <= 1;  //111 / 110 = 1
    16'b01101111_01101111 : OUT <= 1;  //111 / 111 = 1
    16'b01101111_01110000 : OUT <= 0;  //111 / 112 = 0
    16'b01101111_01110001 : OUT <= 0;  //111 / 113 = 0
    16'b01101111_01110010 : OUT <= 0;  //111 / 114 = 0
    16'b01101111_01110011 : OUT <= 0;  //111 / 115 = 0
    16'b01101111_01110100 : OUT <= 0;  //111 / 116 = 0
    16'b01101111_01110101 : OUT <= 0;  //111 / 117 = 0
    16'b01101111_01110110 : OUT <= 0;  //111 / 118 = 0
    16'b01101111_01110111 : OUT <= 0;  //111 / 119 = 0
    16'b01101111_01111000 : OUT <= 0;  //111 / 120 = 0
    16'b01101111_01111001 : OUT <= 0;  //111 / 121 = 0
    16'b01101111_01111010 : OUT <= 0;  //111 / 122 = 0
    16'b01101111_01111011 : OUT <= 0;  //111 / 123 = 0
    16'b01101111_01111100 : OUT <= 0;  //111 / 124 = 0
    16'b01101111_01111101 : OUT <= 0;  //111 / 125 = 0
    16'b01101111_01111110 : OUT <= 0;  //111 / 126 = 0
    16'b01101111_01111111 : OUT <= 0;  //111 / 127 = 0
    16'b01101111_10000000 : OUT <= 0;  //111 / 128 = 0
    16'b01101111_10000001 : OUT <= 0;  //111 / 129 = 0
    16'b01101111_10000010 : OUT <= 0;  //111 / 130 = 0
    16'b01101111_10000011 : OUT <= 0;  //111 / 131 = 0
    16'b01101111_10000100 : OUT <= 0;  //111 / 132 = 0
    16'b01101111_10000101 : OUT <= 0;  //111 / 133 = 0
    16'b01101111_10000110 : OUT <= 0;  //111 / 134 = 0
    16'b01101111_10000111 : OUT <= 0;  //111 / 135 = 0
    16'b01101111_10001000 : OUT <= 0;  //111 / 136 = 0
    16'b01101111_10001001 : OUT <= 0;  //111 / 137 = 0
    16'b01101111_10001010 : OUT <= 0;  //111 / 138 = 0
    16'b01101111_10001011 : OUT <= 0;  //111 / 139 = 0
    16'b01101111_10001100 : OUT <= 0;  //111 / 140 = 0
    16'b01101111_10001101 : OUT <= 0;  //111 / 141 = 0
    16'b01101111_10001110 : OUT <= 0;  //111 / 142 = 0
    16'b01101111_10001111 : OUT <= 0;  //111 / 143 = 0
    16'b01101111_10010000 : OUT <= 0;  //111 / 144 = 0
    16'b01101111_10010001 : OUT <= 0;  //111 / 145 = 0
    16'b01101111_10010010 : OUT <= 0;  //111 / 146 = 0
    16'b01101111_10010011 : OUT <= 0;  //111 / 147 = 0
    16'b01101111_10010100 : OUT <= 0;  //111 / 148 = 0
    16'b01101111_10010101 : OUT <= 0;  //111 / 149 = 0
    16'b01101111_10010110 : OUT <= 0;  //111 / 150 = 0
    16'b01101111_10010111 : OUT <= 0;  //111 / 151 = 0
    16'b01101111_10011000 : OUT <= 0;  //111 / 152 = 0
    16'b01101111_10011001 : OUT <= 0;  //111 / 153 = 0
    16'b01101111_10011010 : OUT <= 0;  //111 / 154 = 0
    16'b01101111_10011011 : OUT <= 0;  //111 / 155 = 0
    16'b01101111_10011100 : OUT <= 0;  //111 / 156 = 0
    16'b01101111_10011101 : OUT <= 0;  //111 / 157 = 0
    16'b01101111_10011110 : OUT <= 0;  //111 / 158 = 0
    16'b01101111_10011111 : OUT <= 0;  //111 / 159 = 0
    16'b01101111_10100000 : OUT <= 0;  //111 / 160 = 0
    16'b01101111_10100001 : OUT <= 0;  //111 / 161 = 0
    16'b01101111_10100010 : OUT <= 0;  //111 / 162 = 0
    16'b01101111_10100011 : OUT <= 0;  //111 / 163 = 0
    16'b01101111_10100100 : OUT <= 0;  //111 / 164 = 0
    16'b01101111_10100101 : OUT <= 0;  //111 / 165 = 0
    16'b01101111_10100110 : OUT <= 0;  //111 / 166 = 0
    16'b01101111_10100111 : OUT <= 0;  //111 / 167 = 0
    16'b01101111_10101000 : OUT <= 0;  //111 / 168 = 0
    16'b01101111_10101001 : OUT <= 0;  //111 / 169 = 0
    16'b01101111_10101010 : OUT <= 0;  //111 / 170 = 0
    16'b01101111_10101011 : OUT <= 0;  //111 / 171 = 0
    16'b01101111_10101100 : OUT <= 0;  //111 / 172 = 0
    16'b01101111_10101101 : OUT <= 0;  //111 / 173 = 0
    16'b01101111_10101110 : OUT <= 0;  //111 / 174 = 0
    16'b01101111_10101111 : OUT <= 0;  //111 / 175 = 0
    16'b01101111_10110000 : OUT <= 0;  //111 / 176 = 0
    16'b01101111_10110001 : OUT <= 0;  //111 / 177 = 0
    16'b01101111_10110010 : OUT <= 0;  //111 / 178 = 0
    16'b01101111_10110011 : OUT <= 0;  //111 / 179 = 0
    16'b01101111_10110100 : OUT <= 0;  //111 / 180 = 0
    16'b01101111_10110101 : OUT <= 0;  //111 / 181 = 0
    16'b01101111_10110110 : OUT <= 0;  //111 / 182 = 0
    16'b01101111_10110111 : OUT <= 0;  //111 / 183 = 0
    16'b01101111_10111000 : OUT <= 0;  //111 / 184 = 0
    16'b01101111_10111001 : OUT <= 0;  //111 / 185 = 0
    16'b01101111_10111010 : OUT <= 0;  //111 / 186 = 0
    16'b01101111_10111011 : OUT <= 0;  //111 / 187 = 0
    16'b01101111_10111100 : OUT <= 0;  //111 / 188 = 0
    16'b01101111_10111101 : OUT <= 0;  //111 / 189 = 0
    16'b01101111_10111110 : OUT <= 0;  //111 / 190 = 0
    16'b01101111_10111111 : OUT <= 0;  //111 / 191 = 0
    16'b01101111_11000000 : OUT <= 0;  //111 / 192 = 0
    16'b01101111_11000001 : OUT <= 0;  //111 / 193 = 0
    16'b01101111_11000010 : OUT <= 0;  //111 / 194 = 0
    16'b01101111_11000011 : OUT <= 0;  //111 / 195 = 0
    16'b01101111_11000100 : OUT <= 0;  //111 / 196 = 0
    16'b01101111_11000101 : OUT <= 0;  //111 / 197 = 0
    16'b01101111_11000110 : OUT <= 0;  //111 / 198 = 0
    16'b01101111_11000111 : OUT <= 0;  //111 / 199 = 0
    16'b01101111_11001000 : OUT <= 0;  //111 / 200 = 0
    16'b01101111_11001001 : OUT <= 0;  //111 / 201 = 0
    16'b01101111_11001010 : OUT <= 0;  //111 / 202 = 0
    16'b01101111_11001011 : OUT <= 0;  //111 / 203 = 0
    16'b01101111_11001100 : OUT <= 0;  //111 / 204 = 0
    16'b01101111_11001101 : OUT <= 0;  //111 / 205 = 0
    16'b01101111_11001110 : OUT <= 0;  //111 / 206 = 0
    16'b01101111_11001111 : OUT <= 0;  //111 / 207 = 0
    16'b01101111_11010000 : OUT <= 0;  //111 / 208 = 0
    16'b01101111_11010001 : OUT <= 0;  //111 / 209 = 0
    16'b01101111_11010010 : OUT <= 0;  //111 / 210 = 0
    16'b01101111_11010011 : OUT <= 0;  //111 / 211 = 0
    16'b01101111_11010100 : OUT <= 0;  //111 / 212 = 0
    16'b01101111_11010101 : OUT <= 0;  //111 / 213 = 0
    16'b01101111_11010110 : OUT <= 0;  //111 / 214 = 0
    16'b01101111_11010111 : OUT <= 0;  //111 / 215 = 0
    16'b01101111_11011000 : OUT <= 0;  //111 / 216 = 0
    16'b01101111_11011001 : OUT <= 0;  //111 / 217 = 0
    16'b01101111_11011010 : OUT <= 0;  //111 / 218 = 0
    16'b01101111_11011011 : OUT <= 0;  //111 / 219 = 0
    16'b01101111_11011100 : OUT <= 0;  //111 / 220 = 0
    16'b01101111_11011101 : OUT <= 0;  //111 / 221 = 0
    16'b01101111_11011110 : OUT <= 0;  //111 / 222 = 0
    16'b01101111_11011111 : OUT <= 0;  //111 / 223 = 0
    16'b01101111_11100000 : OUT <= 0;  //111 / 224 = 0
    16'b01101111_11100001 : OUT <= 0;  //111 / 225 = 0
    16'b01101111_11100010 : OUT <= 0;  //111 / 226 = 0
    16'b01101111_11100011 : OUT <= 0;  //111 / 227 = 0
    16'b01101111_11100100 : OUT <= 0;  //111 / 228 = 0
    16'b01101111_11100101 : OUT <= 0;  //111 / 229 = 0
    16'b01101111_11100110 : OUT <= 0;  //111 / 230 = 0
    16'b01101111_11100111 : OUT <= 0;  //111 / 231 = 0
    16'b01101111_11101000 : OUT <= 0;  //111 / 232 = 0
    16'b01101111_11101001 : OUT <= 0;  //111 / 233 = 0
    16'b01101111_11101010 : OUT <= 0;  //111 / 234 = 0
    16'b01101111_11101011 : OUT <= 0;  //111 / 235 = 0
    16'b01101111_11101100 : OUT <= 0;  //111 / 236 = 0
    16'b01101111_11101101 : OUT <= 0;  //111 / 237 = 0
    16'b01101111_11101110 : OUT <= 0;  //111 / 238 = 0
    16'b01101111_11101111 : OUT <= 0;  //111 / 239 = 0
    16'b01101111_11110000 : OUT <= 0;  //111 / 240 = 0
    16'b01101111_11110001 : OUT <= 0;  //111 / 241 = 0
    16'b01101111_11110010 : OUT <= 0;  //111 / 242 = 0
    16'b01101111_11110011 : OUT <= 0;  //111 / 243 = 0
    16'b01101111_11110100 : OUT <= 0;  //111 / 244 = 0
    16'b01101111_11110101 : OUT <= 0;  //111 / 245 = 0
    16'b01101111_11110110 : OUT <= 0;  //111 / 246 = 0
    16'b01101111_11110111 : OUT <= 0;  //111 / 247 = 0
    16'b01101111_11111000 : OUT <= 0;  //111 / 248 = 0
    16'b01101111_11111001 : OUT <= 0;  //111 / 249 = 0
    16'b01101111_11111010 : OUT <= 0;  //111 / 250 = 0
    16'b01101111_11111011 : OUT <= 0;  //111 / 251 = 0
    16'b01101111_11111100 : OUT <= 0;  //111 / 252 = 0
    16'b01101111_11111101 : OUT <= 0;  //111 / 253 = 0
    16'b01101111_11111110 : OUT <= 0;  //111 / 254 = 0
    16'b01101111_11111111 : OUT <= 0;  //111 / 255 = 0
    16'b01110000_00000000 : OUT <= 0;  //112 / 0 = 0
    16'b01110000_00000001 : OUT <= 112;  //112 / 1 = 112
    16'b01110000_00000010 : OUT <= 56;  //112 / 2 = 56
    16'b01110000_00000011 : OUT <= 37;  //112 / 3 = 37
    16'b01110000_00000100 : OUT <= 28;  //112 / 4 = 28
    16'b01110000_00000101 : OUT <= 22;  //112 / 5 = 22
    16'b01110000_00000110 : OUT <= 18;  //112 / 6 = 18
    16'b01110000_00000111 : OUT <= 16;  //112 / 7 = 16
    16'b01110000_00001000 : OUT <= 14;  //112 / 8 = 14
    16'b01110000_00001001 : OUT <= 12;  //112 / 9 = 12
    16'b01110000_00001010 : OUT <= 11;  //112 / 10 = 11
    16'b01110000_00001011 : OUT <= 10;  //112 / 11 = 10
    16'b01110000_00001100 : OUT <= 9;  //112 / 12 = 9
    16'b01110000_00001101 : OUT <= 8;  //112 / 13 = 8
    16'b01110000_00001110 : OUT <= 8;  //112 / 14 = 8
    16'b01110000_00001111 : OUT <= 7;  //112 / 15 = 7
    16'b01110000_00010000 : OUT <= 7;  //112 / 16 = 7
    16'b01110000_00010001 : OUT <= 6;  //112 / 17 = 6
    16'b01110000_00010010 : OUT <= 6;  //112 / 18 = 6
    16'b01110000_00010011 : OUT <= 5;  //112 / 19 = 5
    16'b01110000_00010100 : OUT <= 5;  //112 / 20 = 5
    16'b01110000_00010101 : OUT <= 5;  //112 / 21 = 5
    16'b01110000_00010110 : OUT <= 5;  //112 / 22 = 5
    16'b01110000_00010111 : OUT <= 4;  //112 / 23 = 4
    16'b01110000_00011000 : OUT <= 4;  //112 / 24 = 4
    16'b01110000_00011001 : OUT <= 4;  //112 / 25 = 4
    16'b01110000_00011010 : OUT <= 4;  //112 / 26 = 4
    16'b01110000_00011011 : OUT <= 4;  //112 / 27 = 4
    16'b01110000_00011100 : OUT <= 4;  //112 / 28 = 4
    16'b01110000_00011101 : OUT <= 3;  //112 / 29 = 3
    16'b01110000_00011110 : OUT <= 3;  //112 / 30 = 3
    16'b01110000_00011111 : OUT <= 3;  //112 / 31 = 3
    16'b01110000_00100000 : OUT <= 3;  //112 / 32 = 3
    16'b01110000_00100001 : OUT <= 3;  //112 / 33 = 3
    16'b01110000_00100010 : OUT <= 3;  //112 / 34 = 3
    16'b01110000_00100011 : OUT <= 3;  //112 / 35 = 3
    16'b01110000_00100100 : OUT <= 3;  //112 / 36 = 3
    16'b01110000_00100101 : OUT <= 3;  //112 / 37 = 3
    16'b01110000_00100110 : OUT <= 2;  //112 / 38 = 2
    16'b01110000_00100111 : OUT <= 2;  //112 / 39 = 2
    16'b01110000_00101000 : OUT <= 2;  //112 / 40 = 2
    16'b01110000_00101001 : OUT <= 2;  //112 / 41 = 2
    16'b01110000_00101010 : OUT <= 2;  //112 / 42 = 2
    16'b01110000_00101011 : OUT <= 2;  //112 / 43 = 2
    16'b01110000_00101100 : OUT <= 2;  //112 / 44 = 2
    16'b01110000_00101101 : OUT <= 2;  //112 / 45 = 2
    16'b01110000_00101110 : OUT <= 2;  //112 / 46 = 2
    16'b01110000_00101111 : OUT <= 2;  //112 / 47 = 2
    16'b01110000_00110000 : OUT <= 2;  //112 / 48 = 2
    16'b01110000_00110001 : OUT <= 2;  //112 / 49 = 2
    16'b01110000_00110010 : OUT <= 2;  //112 / 50 = 2
    16'b01110000_00110011 : OUT <= 2;  //112 / 51 = 2
    16'b01110000_00110100 : OUT <= 2;  //112 / 52 = 2
    16'b01110000_00110101 : OUT <= 2;  //112 / 53 = 2
    16'b01110000_00110110 : OUT <= 2;  //112 / 54 = 2
    16'b01110000_00110111 : OUT <= 2;  //112 / 55 = 2
    16'b01110000_00111000 : OUT <= 2;  //112 / 56 = 2
    16'b01110000_00111001 : OUT <= 1;  //112 / 57 = 1
    16'b01110000_00111010 : OUT <= 1;  //112 / 58 = 1
    16'b01110000_00111011 : OUT <= 1;  //112 / 59 = 1
    16'b01110000_00111100 : OUT <= 1;  //112 / 60 = 1
    16'b01110000_00111101 : OUT <= 1;  //112 / 61 = 1
    16'b01110000_00111110 : OUT <= 1;  //112 / 62 = 1
    16'b01110000_00111111 : OUT <= 1;  //112 / 63 = 1
    16'b01110000_01000000 : OUT <= 1;  //112 / 64 = 1
    16'b01110000_01000001 : OUT <= 1;  //112 / 65 = 1
    16'b01110000_01000010 : OUT <= 1;  //112 / 66 = 1
    16'b01110000_01000011 : OUT <= 1;  //112 / 67 = 1
    16'b01110000_01000100 : OUT <= 1;  //112 / 68 = 1
    16'b01110000_01000101 : OUT <= 1;  //112 / 69 = 1
    16'b01110000_01000110 : OUT <= 1;  //112 / 70 = 1
    16'b01110000_01000111 : OUT <= 1;  //112 / 71 = 1
    16'b01110000_01001000 : OUT <= 1;  //112 / 72 = 1
    16'b01110000_01001001 : OUT <= 1;  //112 / 73 = 1
    16'b01110000_01001010 : OUT <= 1;  //112 / 74 = 1
    16'b01110000_01001011 : OUT <= 1;  //112 / 75 = 1
    16'b01110000_01001100 : OUT <= 1;  //112 / 76 = 1
    16'b01110000_01001101 : OUT <= 1;  //112 / 77 = 1
    16'b01110000_01001110 : OUT <= 1;  //112 / 78 = 1
    16'b01110000_01001111 : OUT <= 1;  //112 / 79 = 1
    16'b01110000_01010000 : OUT <= 1;  //112 / 80 = 1
    16'b01110000_01010001 : OUT <= 1;  //112 / 81 = 1
    16'b01110000_01010010 : OUT <= 1;  //112 / 82 = 1
    16'b01110000_01010011 : OUT <= 1;  //112 / 83 = 1
    16'b01110000_01010100 : OUT <= 1;  //112 / 84 = 1
    16'b01110000_01010101 : OUT <= 1;  //112 / 85 = 1
    16'b01110000_01010110 : OUT <= 1;  //112 / 86 = 1
    16'b01110000_01010111 : OUT <= 1;  //112 / 87 = 1
    16'b01110000_01011000 : OUT <= 1;  //112 / 88 = 1
    16'b01110000_01011001 : OUT <= 1;  //112 / 89 = 1
    16'b01110000_01011010 : OUT <= 1;  //112 / 90 = 1
    16'b01110000_01011011 : OUT <= 1;  //112 / 91 = 1
    16'b01110000_01011100 : OUT <= 1;  //112 / 92 = 1
    16'b01110000_01011101 : OUT <= 1;  //112 / 93 = 1
    16'b01110000_01011110 : OUT <= 1;  //112 / 94 = 1
    16'b01110000_01011111 : OUT <= 1;  //112 / 95 = 1
    16'b01110000_01100000 : OUT <= 1;  //112 / 96 = 1
    16'b01110000_01100001 : OUT <= 1;  //112 / 97 = 1
    16'b01110000_01100010 : OUT <= 1;  //112 / 98 = 1
    16'b01110000_01100011 : OUT <= 1;  //112 / 99 = 1
    16'b01110000_01100100 : OUT <= 1;  //112 / 100 = 1
    16'b01110000_01100101 : OUT <= 1;  //112 / 101 = 1
    16'b01110000_01100110 : OUT <= 1;  //112 / 102 = 1
    16'b01110000_01100111 : OUT <= 1;  //112 / 103 = 1
    16'b01110000_01101000 : OUT <= 1;  //112 / 104 = 1
    16'b01110000_01101001 : OUT <= 1;  //112 / 105 = 1
    16'b01110000_01101010 : OUT <= 1;  //112 / 106 = 1
    16'b01110000_01101011 : OUT <= 1;  //112 / 107 = 1
    16'b01110000_01101100 : OUT <= 1;  //112 / 108 = 1
    16'b01110000_01101101 : OUT <= 1;  //112 / 109 = 1
    16'b01110000_01101110 : OUT <= 1;  //112 / 110 = 1
    16'b01110000_01101111 : OUT <= 1;  //112 / 111 = 1
    16'b01110000_01110000 : OUT <= 1;  //112 / 112 = 1
    16'b01110000_01110001 : OUT <= 0;  //112 / 113 = 0
    16'b01110000_01110010 : OUT <= 0;  //112 / 114 = 0
    16'b01110000_01110011 : OUT <= 0;  //112 / 115 = 0
    16'b01110000_01110100 : OUT <= 0;  //112 / 116 = 0
    16'b01110000_01110101 : OUT <= 0;  //112 / 117 = 0
    16'b01110000_01110110 : OUT <= 0;  //112 / 118 = 0
    16'b01110000_01110111 : OUT <= 0;  //112 / 119 = 0
    16'b01110000_01111000 : OUT <= 0;  //112 / 120 = 0
    16'b01110000_01111001 : OUT <= 0;  //112 / 121 = 0
    16'b01110000_01111010 : OUT <= 0;  //112 / 122 = 0
    16'b01110000_01111011 : OUT <= 0;  //112 / 123 = 0
    16'b01110000_01111100 : OUT <= 0;  //112 / 124 = 0
    16'b01110000_01111101 : OUT <= 0;  //112 / 125 = 0
    16'b01110000_01111110 : OUT <= 0;  //112 / 126 = 0
    16'b01110000_01111111 : OUT <= 0;  //112 / 127 = 0
    16'b01110000_10000000 : OUT <= 0;  //112 / 128 = 0
    16'b01110000_10000001 : OUT <= 0;  //112 / 129 = 0
    16'b01110000_10000010 : OUT <= 0;  //112 / 130 = 0
    16'b01110000_10000011 : OUT <= 0;  //112 / 131 = 0
    16'b01110000_10000100 : OUT <= 0;  //112 / 132 = 0
    16'b01110000_10000101 : OUT <= 0;  //112 / 133 = 0
    16'b01110000_10000110 : OUT <= 0;  //112 / 134 = 0
    16'b01110000_10000111 : OUT <= 0;  //112 / 135 = 0
    16'b01110000_10001000 : OUT <= 0;  //112 / 136 = 0
    16'b01110000_10001001 : OUT <= 0;  //112 / 137 = 0
    16'b01110000_10001010 : OUT <= 0;  //112 / 138 = 0
    16'b01110000_10001011 : OUT <= 0;  //112 / 139 = 0
    16'b01110000_10001100 : OUT <= 0;  //112 / 140 = 0
    16'b01110000_10001101 : OUT <= 0;  //112 / 141 = 0
    16'b01110000_10001110 : OUT <= 0;  //112 / 142 = 0
    16'b01110000_10001111 : OUT <= 0;  //112 / 143 = 0
    16'b01110000_10010000 : OUT <= 0;  //112 / 144 = 0
    16'b01110000_10010001 : OUT <= 0;  //112 / 145 = 0
    16'b01110000_10010010 : OUT <= 0;  //112 / 146 = 0
    16'b01110000_10010011 : OUT <= 0;  //112 / 147 = 0
    16'b01110000_10010100 : OUT <= 0;  //112 / 148 = 0
    16'b01110000_10010101 : OUT <= 0;  //112 / 149 = 0
    16'b01110000_10010110 : OUT <= 0;  //112 / 150 = 0
    16'b01110000_10010111 : OUT <= 0;  //112 / 151 = 0
    16'b01110000_10011000 : OUT <= 0;  //112 / 152 = 0
    16'b01110000_10011001 : OUT <= 0;  //112 / 153 = 0
    16'b01110000_10011010 : OUT <= 0;  //112 / 154 = 0
    16'b01110000_10011011 : OUT <= 0;  //112 / 155 = 0
    16'b01110000_10011100 : OUT <= 0;  //112 / 156 = 0
    16'b01110000_10011101 : OUT <= 0;  //112 / 157 = 0
    16'b01110000_10011110 : OUT <= 0;  //112 / 158 = 0
    16'b01110000_10011111 : OUT <= 0;  //112 / 159 = 0
    16'b01110000_10100000 : OUT <= 0;  //112 / 160 = 0
    16'b01110000_10100001 : OUT <= 0;  //112 / 161 = 0
    16'b01110000_10100010 : OUT <= 0;  //112 / 162 = 0
    16'b01110000_10100011 : OUT <= 0;  //112 / 163 = 0
    16'b01110000_10100100 : OUT <= 0;  //112 / 164 = 0
    16'b01110000_10100101 : OUT <= 0;  //112 / 165 = 0
    16'b01110000_10100110 : OUT <= 0;  //112 / 166 = 0
    16'b01110000_10100111 : OUT <= 0;  //112 / 167 = 0
    16'b01110000_10101000 : OUT <= 0;  //112 / 168 = 0
    16'b01110000_10101001 : OUT <= 0;  //112 / 169 = 0
    16'b01110000_10101010 : OUT <= 0;  //112 / 170 = 0
    16'b01110000_10101011 : OUT <= 0;  //112 / 171 = 0
    16'b01110000_10101100 : OUT <= 0;  //112 / 172 = 0
    16'b01110000_10101101 : OUT <= 0;  //112 / 173 = 0
    16'b01110000_10101110 : OUT <= 0;  //112 / 174 = 0
    16'b01110000_10101111 : OUT <= 0;  //112 / 175 = 0
    16'b01110000_10110000 : OUT <= 0;  //112 / 176 = 0
    16'b01110000_10110001 : OUT <= 0;  //112 / 177 = 0
    16'b01110000_10110010 : OUT <= 0;  //112 / 178 = 0
    16'b01110000_10110011 : OUT <= 0;  //112 / 179 = 0
    16'b01110000_10110100 : OUT <= 0;  //112 / 180 = 0
    16'b01110000_10110101 : OUT <= 0;  //112 / 181 = 0
    16'b01110000_10110110 : OUT <= 0;  //112 / 182 = 0
    16'b01110000_10110111 : OUT <= 0;  //112 / 183 = 0
    16'b01110000_10111000 : OUT <= 0;  //112 / 184 = 0
    16'b01110000_10111001 : OUT <= 0;  //112 / 185 = 0
    16'b01110000_10111010 : OUT <= 0;  //112 / 186 = 0
    16'b01110000_10111011 : OUT <= 0;  //112 / 187 = 0
    16'b01110000_10111100 : OUT <= 0;  //112 / 188 = 0
    16'b01110000_10111101 : OUT <= 0;  //112 / 189 = 0
    16'b01110000_10111110 : OUT <= 0;  //112 / 190 = 0
    16'b01110000_10111111 : OUT <= 0;  //112 / 191 = 0
    16'b01110000_11000000 : OUT <= 0;  //112 / 192 = 0
    16'b01110000_11000001 : OUT <= 0;  //112 / 193 = 0
    16'b01110000_11000010 : OUT <= 0;  //112 / 194 = 0
    16'b01110000_11000011 : OUT <= 0;  //112 / 195 = 0
    16'b01110000_11000100 : OUT <= 0;  //112 / 196 = 0
    16'b01110000_11000101 : OUT <= 0;  //112 / 197 = 0
    16'b01110000_11000110 : OUT <= 0;  //112 / 198 = 0
    16'b01110000_11000111 : OUT <= 0;  //112 / 199 = 0
    16'b01110000_11001000 : OUT <= 0;  //112 / 200 = 0
    16'b01110000_11001001 : OUT <= 0;  //112 / 201 = 0
    16'b01110000_11001010 : OUT <= 0;  //112 / 202 = 0
    16'b01110000_11001011 : OUT <= 0;  //112 / 203 = 0
    16'b01110000_11001100 : OUT <= 0;  //112 / 204 = 0
    16'b01110000_11001101 : OUT <= 0;  //112 / 205 = 0
    16'b01110000_11001110 : OUT <= 0;  //112 / 206 = 0
    16'b01110000_11001111 : OUT <= 0;  //112 / 207 = 0
    16'b01110000_11010000 : OUT <= 0;  //112 / 208 = 0
    16'b01110000_11010001 : OUT <= 0;  //112 / 209 = 0
    16'b01110000_11010010 : OUT <= 0;  //112 / 210 = 0
    16'b01110000_11010011 : OUT <= 0;  //112 / 211 = 0
    16'b01110000_11010100 : OUT <= 0;  //112 / 212 = 0
    16'b01110000_11010101 : OUT <= 0;  //112 / 213 = 0
    16'b01110000_11010110 : OUT <= 0;  //112 / 214 = 0
    16'b01110000_11010111 : OUT <= 0;  //112 / 215 = 0
    16'b01110000_11011000 : OUT <= 0;  //112 / 216 = 0
    16'b01110000_11011001 : OUT <= 0;  //112 / 217 = 0
    16'b01110000_11011010 : OUT <= 0;  //112 / 218 = 0
    16'b01110000_11011011 : OUT <= 0;  //112 / 219 = 0
    16'b01110000_11011100 : OUT <= 0;  //112 / 220 = 0
    16'b01110000_11011101 : OUT <= 0;  //112 / 221 = 0
    16'b01110000_11011110 : OUT <= 0;  //112 / 222 = 0
    16'b01110000_11011111 : OUT <= 0;  //112 / 223 = 0
    16'b01110000_11100000 : OUT <= 0;  //112 / 224 = 0
    16'b01110000_11100001 : OUT <= 0;  //112 / 225 = 0
    16'b01110000_11100010 : OUT <= 0;  //112 / 226 = 0
    16'b01110000_11100011 : OUT <= 0;  //112 / 227 = 0
    16'b01110000_11100100 : OUT <= 0;  //112 / 228 = 0
    16'b01110000_11100101 : OUT <= 0;  //112 / 229 = 0
    16'b01110000_11100110 : OUT <= 0;  //112 / 230 = 0
    16'b01110000_11100111 : OUT <= 0;  //112 / 231 = 0
    16'b01110000_11101000 : OUT <= 0;  //112 / 232 = 0
    16'b01110000_11101001 : OUT <= 0;  //112 / 233 = 0
    16'b01110000_11101010 : OUT <= 0;  //112 / 234 = 0
    16'b01110000_11101011 : OUT <= 0;  //112 / 235 = 0
    16'b01110000_11101100 : OUT <= 0;  //112 / 236 = 0
    16'b01110000_11101101 : OUT <= 0;  //112 / 237 = 0
    16'b01110000_11101110 : OUT <= 0;  //112 / 238 = 0
    16'b01110000_11101111 : OUT <= 0;  //112 / 239 = 0
    16'b01110000_11110000 : OUT <= 0;  //112 / 240 = 0
    16'b01110000_11110001 : OUT <= 0;  //112 / 241 = 0
    16'b01110000_11110010 : OUT <= 0;  //112 / 242 = 0
    16'b01110000_11110011 : OUT <= 0;  //112 / 243 = 0
    16'b01110000_11110100 : OUT <= 0;  //112 / 244 = 0
    16'b01110000_11110101 : OUT <= 0;  //112 / 245 = 0
    16'b01110000_11110110 : OUT <= 0;  //112 / 246 = 0
    16'b01110000_11110111 : OUT <= 0;  //112 / 247 = 0
    16'b01110000_11111000 : OUT <= 0;  //112 / 248 = 0
    16'b01110000_11111001 : OUT <= 0;  //112 / 249 = 0
    16'b01110000_11111010 : OUT <= 0;  //112 / 250 = 0
    16'b01110000_11111011 : OUT <= 0;  //112 / 251 = 0
    16'b01110000_11111100 : OUT <= 0;  //112 / 252 = 0
    16'b01110000_11111101 : OUT <= 0;  //112 / 253 = 0
    16'b01110000_11111110 : OUT <= 0;  //112 / 254 = 0
    16'b01110000_11111111 : OUT <= 0;  //112 / 255 = 0
    16'b01110001_00000000 : OUT <= 0;  //113 / 0 = 0
    16'b01110001_00000001 : OUT <= 113;  //113 / 1 = 113
    16'b01110001_00000010 : OUT <= 56;  //113 / 2 = 56
    16'b01110001_00000011 : OUT <= 37;  //113 / 3 = 37
    16'b01110001_00000100 : OUT <= 28;  //113 / 4 = 28
    16'b01110001_00000101 : OUT <= 22;  //113 / 5 = 22
    16'b01110001_00000110 : OUT <= 18;  //113 / 6 = 18
    16'b01110001_00000111 : OUT <= 16;  //113 / 7 = 16
    16'b01110001_00001000 : OUT <= 14;  //113 / 8 = 14
    16'b01110001_00001001 : OUT <= 12;  //113 / 9 = 12
    16'b01110001_00001010 : OUT <= 11;  //113 / 10 = 11
    16'b01110001_00001011 : OUT <= 10;  //113 / 11 = 10
    16'b01110001_00001100 : OUT <= 9;  //113 / 12 = 9
    16'b01110001_00001101 : OUT <= 8;  //113 / 13 = 8
    16'b01110001_00001110 : OUT <= 8;  //113 / 14 = 8
    16'b01110001_00001111 : OUT <= 7;  //113 / 15 = 7
    16'b01110001_00010000 : OUT <= 7;  //113 / 16 = 7
    16'b01110001_00010001 : OUT <= 6;  //113 / 17 = 6
    16'b01110001_00010010 : OUT <= 6;  //113 / 18 = 6
    16'b01110001_00010011 : OUT <= 5;  //113 / 19 = 5
    16'b01110001_00010100 : OUT <= 5;  //113 / 20 = 5
    16'b01110001_00010101 : OUT <= 5;  //113 / 21 = 5
    16'b01110001_00010110 : OUT <= 5;  //113 / 22 = 5
    16'b01110001_00010111 : OUT <= 4;  //113 / 23 = 4
    16'b01110001_00011000 : OUT <= 4;  //113 / 24 = 4
    16'b01110001_00011001 : OUT <= 4;  //113 / 25 = 4
    16'b01110001_00011010 : OUT <= 4;  //113 / 26 = 4
    16'b01110001_00011011 : OUT <= 4;  //113 / 27 = 4
    16'b01110001_00011100 : OUT <= 4;  //113 / 28 = 4
    16'b01110001_00011101 : OUT <= 3;  //113 / 29 = 3
    16'b01110001_00011110 : OUT <= 3;  //113 / 30 = 3
    16'b01110001_00011111 : OUT <= 3;  //113 / 31 = 3
    16'b01110001_00100000 : OUT <= 3;  //113 / 32 = 3
    16'b01110001_00100001 : OUT <= 3;  //113 / 33 = 3
    16'b01110001_00100010 : OUT <= 3;  //113 / 34 = 3
    16'b01110001_00100011 : OUT <= 3;  //113 / 35 = 3
    16'b01110001_00100100 : OUT <= 3;  //113 / 36 = 3
    16'b01110001_00100101 : OUT <= 3;  //113 / 37 = 3
    16'b01110001_00100110 : OUT <= 2;  //113 / 38 = 2
    16'b01110001_00100111 : OUT <= 2;  //113 / 39 = 2
    16'b01110001_00101000 : OUT <= 2;  //113 / 40 = 2
    16'b01110001_00101001 : OUT <= 2;  //113 / 41 = 2
    16'b01110001_00101010 : OUT <= 2;  //113 / 42 = 2
    16'b01110001_00101011 : OUT <= 2;  //113 / 43 = 2
    16'b01110001_00101100 : OUT <= 2;  //113 / 44 = 2
    16'b01110001_00101101 : OUT <= 2;  //113 / 45 = 2
    16'b01110001_00101110 : OUT <= 2;  //113 / 46 = 2
    16'b01110001_00101111 : OUT <= 2;  //113 / 47 = 2
    16'b01110001_00110000 : OUT <= 2;  //113 / 48 = 2
    16'b01110001_00110001 : OUT <= 2;  //113 / 49 = 2
    16'b01110001_00110010 : OUT <= 2;  //113 / 50 = 2
    16'b01110001_00110011 : OUT <= 2;  //113 / 51 = 2
    16'b01110001_00110100 : OUT <= 2;  //113 / 52 = 2
    16'b01110001_00110101 : OUT <= 2;  //113 / 53 = 2
    16'b01110001_00110110 : OUT <= 2;  //113 / 54 = 2
    16'b01110001_00110111 : OUT <= 2;  //113 / 55 = 2
    16'b01110001_00111000 : OUT <= 2;  //113 / 56 = 2
    16'b01110001_00111001 : OUT <= 1;  //113 / 57 = 1
    16'b01110001_00111010 : OUT <= 1;  //113 / 58 = 1
    16'b01110001_00111011 : OUT <= 1;  //113 / 59 = 1
    16'b01110001_00111100 : OUT <= 1;  //113 / 60 = 1
    16'b01110001_00111101 : OUT <= 1;  //113 / 61 = 1
    16'b01110001_00111110 : OUT <= 1;  //113 / 62 = 1
    16'b01110001_00111111 : OUT <= 1;  //113 / 63 = 1
    16'b01110001_01000000 : OUT <= 1;  //113 / 64 = 1
    16'b01110001_01000001 : OUT <= 1;  //113 / 65 = 1
    16'b01110001_01000010 : OUT <= 1;  //113 / 66 = 1
    16'b01110001_01000011 : OUT <= 1;  //113 / 67 = 1
    16'b01110001_01000100 : OUT <= 1;  //113 / 68 = 1
    16'b01110001_01000101 : OUT <= 1;  //113 / 69 = 1
    16'b01110001_01000110 : OUT <= 1;  //113 / 70 = 1
    16'b01110001_01000111 : OUT <= 1;  //113 / 71 = 1
    16'b01110001_01001000 : OUT <= 1;  //113 / 72 = 1
    16'b01110001_01001001 : OUT <= 1;  //113 / 73 = 1
    16'b01110001_01001010 : OUT <= 1;  //113 / 74 = 1
    16'b01110001_01001011 : OUT <= 1;  //113 / 75 = 1
    16'b01110001_01001100 : OUT <= 1;  //113 / 76 = 1
    16'b01110001_01001101 : OUT <= 1;  //113 / 77 = 1
    16'b01110001_01001110 : OUT <= 1;  //113 / 78 = 1
    16'b01110001_01001111 : OUT <= 1;  //113 / 79 = 1
    16'b01110001_01010000 : OUT <= 1;  //113 / 80 = 1
    16'b01110001_01010001 : OUT <= 1;  //113 / 81 = 1
    16'b01110001_01010010 : OUT <= 1;  //113 / 82 = 1
    16'b01110001_01010011 : OUT <= 1;  //113 / 83 = 1
    16'b01110001_01010100 : OUT <= 1;  //113 / 84 = 1
    16'b01110001_01010101 : OUT <= 1;  //113 / 85 = 1
    16'b01110001_01010110 : OUT <= 1;  //113 / 86 = 1
    16'b01110001_01010111 : OUT <= 1;  //113 / 87 = 1
    16'b01110001_01011000 : OUT <= 1;  //113 / 88 = 1
    16'b01110001_01011001 : OUT <= 1;  //113 / 89 = 1
    16'b01110001_01011010 : OUT <= 1;  //113 / 90 = 1
    16'b01110001_01011011 : OUT <= 1;  //113 / 91 = 1
    16'b01110001_01011100 : OUT <= 1;  //113 / 92 = 1
    16'b01110001_01011101 : OUT <= 1;  //113 / 93 = 1
    16'b01110001_01011110 : OUT <= 1;  //113 / 94 = 1
    16'b01110001_01011111 : OUT <= 1;  //113 / 95 = 1
    16'b01110001_01100000 : OUT <= 1;  //113 / 96 = 1
    16'b01110001_01100001 : OUT <= 1;  //113 / 97 = 1
    16'b01110001_01100010 : OUT <= 1;  //113 / 98 = 1
    16'b01110001_01100011 : OUT <= 1;  //113 / 99 = 1
    16'b01110001_01100100 : OUT <= 1;  //113 / 100 = 1
    16'b01110001_01100101 : OUT <= 1;  //113 / 101 = 1
    16'b01110001_01100110 : OUT <= 1;  //113 / 102 = 1
    16'b01110001_01100111 : OUT <= 1;  //113 / 103 = 1
    16'b01110001_01101000 : OUT <= 1;  //113 / 104 = 1
    16'b01110001_01101001 : OUT <= 1;  //113 / 105 = 1
    16'b01110001_01101010 : OUT <= 1;  //113 / 106 = 1
    16'b01110001_01101011 : OUT <= 1;  //113 / 107 = 1
    16'b01110001_01101100 : OUT <= 1;  //113 / 108 = 1
    16'b01110001_01101101 : OUT <= 1;  //113 / 109 = 1
    16'b01110001_01101110 : OUT <= 1;  //113 / 110 = 1
    16'b01110001_01101111 : OUT <= 1;  //113 / 111 = 1
    16'b01110001_01110000 : OUT <= 1;  //113 / 112 = 1
    16'b01110001_01110001 : OUT <= 1;  //113 / 113 = 1
    16'b01110001_01110010 : OUT <= 0;  //113 / 114 = 0
    16'b01110001_01110011 : OUT <= 0;  //113 / 115 = 0
    16'b01110001_01110100 : OUT <= 0;  //113 / 116 = 0
    16'b01110001_01110101 : OUT <= 0;  //113 / 117 = 0
    16'b01110001_01110110 : OUT <= 0;  //113 / 118 = 0
    16'b01110001_01110111 : OUT <= 0;  //113 / 119 = 0
    16'b01110001_01111000 : OUT <= 0;  //113 / 120 = 0
    16'b01110001_01111001 : OUT <= 0;  //113 / 121 = 0
    16'b01110001_01111010 : OUT <= 0;  //113 / 122 = 0
    16'b01110001_01111011 : OUT <= 0;  //113 / 123 = 0
    16'b01110001_01111100 : OUT <= 0;  //113 / 124 = 0
    16'b01110001_01111101 : OUT <= 0;  //113 / 125 = 0
    16'b01110001_01111110 : OUT <= 0;  //113 / 126 = 0
    16'b01110001_01111111 : OUT <= 0;  //113 / 127 = 0
    16'b01110001_10000000 : OUT <= 0;  //113 / 128 = 0
    16'b01110001_10000001 : OUT <= 0;  //113 / 129 = 0
    16'b01110001_10000010 : OUT <= 0;  //113 / 130 = 0
    16'b01110001_10000011 : OUT <= 0;  //113 / 131 = 0
    16'b01110001_10000100 : OUT <= 0;  //113 / 132 = 0
    16'b01110001_10000101 : OUT <= 0;  //113 / 133 = 0
    16'b01110001_10000110 : OUT <= 0;  //113 / 134 = 0
    16'b01110001_10000111 : OUT <= 0;  //113 / 135 = 0
    16'b01110001_10001000 : OUT <= 0;  //113 / 136 = 0
    16'b01110001_10001001 : OUT <= 0;  //113 / 137 = 0
    16'b01110001_10001010 : OUT <= 0;  //113 / 138 = 0
    16'b01110001_10001011 : OUT <= 0;  //113 / 139 = 0
    16'b01110001_10001100 : OUT <= 0;  //113 / 140 = 0
    16'b01110001_10001101 : OUT <= 0;  //113 / 141 = 0
    16'b01110001_10001110 : OUT <= 0;  //113 / 142 = 0
    16'b01110001_10001111 : OUT <= 0;  //113 / 143 = 0
    16'b01110001_10010000 : OUT <= 0;  //113 / 144 = 0
    16'b01110001_10010001 : OUT <= 0;  //113 / 145 = 0
    16'b01110001_10010010 : OUT <= 0;  //113 / 146 = 0
    16'b01110001_10010011 : OUT <= 0;  //113 / 147 = 0
    16'b01110001_10010100 : OUT <= 0;  //113 / 148 = 0
    16'b01110001_10010101 : OUT <= 0;  //113 / 149 = 0
    16'b01110001_10010110 : OUT <= 0;  //113 / 150 = 0
    16'b01110001_10010111 : OUT <= 0;  //113 / 151 = 0
    16'b01110001_10011000 : OUT <= 0;  //113 / 152 = 0
    16'b01110001_10011001 : OUT <= 0;  //113 / 153 = 0
    16'b01110001_10011010 : OUT <= 0;  //113 / 154 = 0
    16'b01110001_10011011 : OUT <= 0;  //113 / 155 = 0
    16'b01110001_10011100 : OUT <= 0;  //113 / 156 = 0
    16'b01110001_10011101 : OUT <= 0;  //113 / 157 = 0
    16'b01110001_10011110 : OUT <= 0;  //113 / 158 = 0
    16'b01110001_10011111 : OUT <= 0;  //113 / 159 = 0
    16'b01110001_10100000 : OUT <= 0;  //113 / 160 = 0
    16'b01110001_10100001 : OUT <= 0;  //113 / 161 = 0
    16'b01110001_10100010 : OUT <= 0;  //113 / 162 = 0
    16'b01110001_10100011 : OUT <= 0;  //113 / 163 = 0
    16'b01110001_10100100 : OUT <= 0;  //113 / 164 = 0
    16'b01110001_10100101 : OUT <= 0;  //113 / 165 = 0
    16'b01110001_10100110 : OUT <= 0;  //113 / 166 = 0
    16'b01110001_10100111 : OUT <= 0;  //113 / 167 = 0
    16'b01110001_10101000 : OUT <= 0;  //113 / 168 = 0
    16'b01110001_10101001 : OUT <= 0;  //113 / 169 = 0
    16'b01110001_10101010 : OUT <= 0;  //113 / 170 = 0
    16'b01110001_10101011 : OUT <= 0;  //113 / 171 = 0
    16'b01110001_10101100 : OUT <= 0;  //113 / 172 = 0
    16'b01110001_10101101 : OUT <= 0;  //113 / 173 = 0
    16'b01110001_10101110 : OUT <= 0;  //113 / 174 = 0
    16'b01110001_10101111 : OUT <= 0;  //113 / 175 = 0
    16'b01110001_10110000 : OUT <= 0;  //113 / 176 = 0
    16'b01110001_10110001 : OUT <= 0;  //113 / 177 = 0
    16'b01110001_10110010 : OUT <= 0;  //113 / 178 = 0
    16'b01110001_10110011 : OUT <= 0;  //113 / 179 = 0
    16'b01110001_10110100 : OUT <= 0;  //113 / 180 = 0
    16'b01110001_10110101 : OUT <= 0;  //113 / 181 = 0
    16'b01110001_10110110 : OUT <= 0;  //113 / 182 = 0
    16'b01110001_10110111 : OUT <= 0;  //113 / 183 = 0
    16'b01110001_10111000 : OUT <= 0;  //113 / 184 = 0
    16'b01110001_10111001 : OUT <= 0;  //113 / 185 = 0
    16'b01110001_10111010 : OUT <= 0;  //113 / 186 = 0
    16'b01110001_10111011 : OUT <= 0;  //113 / 187 = 0
    16'b01110001_10111100 : OUT <= 0;  //113 / 188 = 0
    16'b01110001_10111101 : OUT <= 0;  //113 / 189 = 0
    16'b01110001_10111110 : OUT <= 0;  //113 / 190 = 0
    16'b01110001_10111111 : OUT <= 0;  //113 / 191 = 0
    16'b01110001_11000000 : OUT <= 0;  //113 / 192 = 0
    16'b01110001_11000001 : OUT <= 0;  //113 / 193 = 0
    16'b01110001_11000010 : OUT <= 0;  //113 / 194 = 0
    16'b01110001_11000011 : OUT <= 0;  //113 / 195 = 0
    16'b01110001_11000100 : OUT <= 0;  //113 / 196 = 0
    16'b01110001_11000101 : OUT <= 0;  //113 / 197 = 0
    16'b01110001_11000110 : OUT <= 0;  //113 / 198 = 0
    16'b01110001_11000111 : OUT <= 0;  //113 / 199 = 0
    16'b01110001_11001000 : OUT <= 0;  //113 / 200 = 0
    16'b01110001_11001001 : OUT <= 0;  //113 / 201 = 0
    16'b01110001_11001010 : OUT <= 0;  //113 / 202 = 0
    16'b01110001_11001011 : OUT <= 0;  //113 / 203 = 0
    16'b01110001_11001100 : OUT <= 0;  //113 / 204 = 0
    16'b01110001_11001101 : OUT <= 0;  //113 / 205 = 0
    16'b01110001_11001110 : OUT <= 0;  //113 / 206 = 0
    16'b01110001_11001111 : OUT <= 0;  //113 / 207 = 0
    16'b01110001_11010000 : OUT <= 0;  //113 / 208 = 0
    16'b01110001_11010001 : OUT <= 0;  //113 / 209 = 0
    16'b01110001_11010010 : OUT <= 0;  //113 / 210 = 0
    16'b01110001_11010011 : OUT <= 0;  //113 / 211 = 0
    16'b01110001_11010100 : OUT <= 0;  //113 / 212 = 0
    16'b01110001_11010101 : OUT <= 0;  //113 / 213 = 0
    16'b01110001_11010110 : OUT <= 0;  //113 / 214 = 0
    16'b01110001_11010111 : OUT <= 0;  //113 / 215 = 0
    16'b01110001_11011000 : OUT <= 0;  //113 / 216 = 0
    16'b01110001_11011001 : OUT <= 0;  //113 / 217 = 0
    16'b01110001_11011010 : OUT <= 0;  //113 / 218 = 0
    16'b01110001_11011011 : OUT <= 0;  //113 / 219 = 0
    16'b01110001_11011100 : OUT <= 0;  //113 / 220 = 0
    16'b01110001_11011101 : OUT <= 0;  //113 / 221 = 0
    16'b01110001_11011110 : OUT <= 0;  //113 / 222 = 0
    16'b01110001_11011111 : OUT <= 0;  //113 / 223 = 0
    16'b01110001_11100000 : OUT <= 0;  //113 / 224 = 0
    16'b01110001_11100001 : OUT <= 0;  //113 / 225 = 0
    16'b01110001_11100010 : OUT <= 0;  //113 / 226 = 0
    16'b01110001_11100011 : OUT <= 0;  //113 / 227 = 0
    16'b01110001_11100100 : OUT <= 0;  //113 / 228 = 0
    16'b01110001_11100101 : OUT <= 0;  //113 / 229 = 0
    16'b01110001_11100110 : OUT <= 0;  //113 / 230 = 0
    16'b01110001_11100111 : OUT <= 0;  //113 / 231 = 0
    16'b01110001_11101000 : OUT <= 0;  //113 / 232 = 0
    16'b01110001_11101001 : OUT <= 0;  //113 / 233 = 0
    16'b01110001_11101010 : OUT <= 0;  //113 / 234 = 0
    16'b01110001_11101011 : OUT <= 0;  //113 / 235 = 0
    16'b01110001_11101100 : OUT <= 0;  //113 / 236 = 0
    16'b01110001_11101101 : OUT <= 0;  //113 / 237 = 0
    16'b01110001_11101110 : OUT <= 0;  //113 / 238 = 0
    16'b01110001_11101111 : OUT <= 0;  //113 / 239 = 0
    16'b01110001_11110000 : OUT <= 0;  //113 / 240 = 0
    16'b01110001_11110001 : OUT <= 0;  //113 / 241 = 0
    16'b01110001_11110010 : OUT <= 0;  //113 / 242 = 0
    16'b01110001_11110011 : OUT <= 0;  //113 / 243 = 0
    16'b01110001_11110100 : OUT <= 0;  //113 / 244 = 0
    16'b01110001_11110101 : OUT <= 0;  //113 / 245 = 0
    16'b01110001_11110110 : OUT <= 0;  //113 / 246 = 0
    16'b01110001_11110111 : OUT <= 0;  //113 / 247 = 0
    16'b01110001_11111000 : OUT <= 0;  //113 / 248 = 0
    16'b01110001_11111001 : OUT <= 0;  //113 / 249 = 0
    16'b01110001_11111010 : OUT <= 0;  //113 / 250 = 0
    16'b01110001_11111011 : OUT <= 0;  //113 / 251 = 0
    16'b01110001_11111100 : OUT <= 0;  //113 / 252 = 0
    16'b01110001_11111101 : OUT <= 0;  //113 / 253 = 0
    16'b01110001_11111110 : OUT <= 0;  //113 / 254 = 0
    16'b01110001_11111111 : OUT <= 0;  //113 / 255 = 0
    16'b01110010_00000000 : OUT <= 0;  //114 / 0 = 0
    16'b01110010_00000001 : OUT <= 114;  //114 / 1 = 114
    16'b01110010_00000010 : OUT <= 57;  //114 / 2 = 57
    16'b01110010_00000011 : OUT <= 38;  //114 / 3 = 38
    16'b01110010_00000100 : OUT <= 28;  //114 / 4 = 28
    16'b01110010_00000101 : OUT <= 22;  //114 / 5 = 22
    16'b01110010_00000110 : OUT <= 19;  //114 / 6 = 19
    16'b01110010_00000111 : OUT <= 16;  //114 / 7 = 16
    16'b01110010_00001000 : OUT <= 14;  //114 / 8 = 14
    16'b01110010_00001001 : OUT <= 12;  //114 / 9 = 12
    16'b01110010_00001010 : OUT <= 11;  //114 / 10 = 11
    16'b01110010_00001011 : OUT <= 10;  //114 / 11 = 10
    16'b01110010_00001100 : OUT <= 9;  //114 / 12 = 9
    16'b01110010_00001101 : OUT <= 8;  //114 / 13 = 8
    16'b01110010_00001110 : OUT <= 8;  //114 / 14 = 8
    16'b01110010_00001111 : OUT <= 7;  //114 / 15 = 7
    16'b01110010_00010000 : OUT <= 7;  //114 / 16 = 7
    16'b01110010_00010001 : OUT <= 6;  //114 / 17 = 6
    16'b01110010_00010010 : OUT <= 6;  //114 / 18 = 6
    16'b01110010_00010011 : OUT <= 6;  //114 / 19 = 6
    16'b01110010_00010100 : OUT <= 5;  //114 / 20 = 5
    16'b01110010_00010101 : OUT <= 5;  //114 / 21 = 5
    16'b01110010_00010110 : OUT <= 5;  //114 / 22 = 5
    16'b01110010_00010111 : OUT <= 4;  //114 / 23 = 4
    16'b01110010_00011000 : OUT <= 4;  //114 / 24 = 4
    16'b01110010_00011001 : OUT <= 4;  //114 / 25 = 4
    16'b01110010_00011010 : OUT <= 4;  //114 / 26 = 4
    16'b01110010_00011011 : OUT <= 4;  //114 / 27 = 4
    16'b01110010_00011100 : OUT <= 4;  //114 / 28 = 4
    16'b01110010_00011101 : OUT <= 3;  //114 / 29 = 3
    16'b01110010_00011110 : OUT <= 3;  //114 / 30 = 3
    16'b01110010_00011111 : OUT <= 3;  //114 / 31 = 3
    16'b01110010_00100000 : OUT <= 3;  //114 / 32 = 3
    16'b01110010_00100001 : OUT <= 3;  //114 / 33 = 3
    16'b01110010_00100010 : OUT <= 3;  //114 / 34 = 3
    16'b01110010_00100011 : OUT <= 3;  //114 / 35 = 3
    16'b01110010_00100100 : OUT <= 3;  //114 / 36 = 3
    16'b01110010_00100101 : OUT <= 3;  //114 / 37 = 3
    16'b01110010_00100110 : OUT <= 3;  //114 / 38 = 3
    16'b01110010_00100111 : OUT <= 2;  //114 / 39 = 2
    16'b01110010_00101000 : OUT <= 2;  //114 / 40 = 2
    16'b01110010_00101001 : OUT <= 2;  //114 / 41 = 2
    16'b01110010_00101010 : OUT <= 2;  //114 / 42 = 2
    16'b01110010_00101011 : OUT <= 2;  //114 / 43 = 2
    16'b01110010_00101100 : OUT <= 2;  //114 / 44 = 2
    16'b01110010_00101101 : OUT <= 2;  //114 / 45 = 2
    16'b01110010_00101110 : OUT <= 2;  //114 / 46 = 2
    16'b01110010_00101111 : OUT <= 2;  //114 / 47 = 2
    16'b01110010_00110000 : OUT <= 2;  //114 / 48 = 2
    16'b01110010_00110001 : OUT <= 2;  //114 / 49 = 2
    16'b01110010_00110010 : OUT <= 2;  //114 / 50 = 2
    16'b01110010_00110011 : OUT <= 2;  //114 / 51 = 2
    16'b01110010_00110100 : OUT <= 2;  //114 / 52 = 2
    16'b01110010_00110101 : OUT <= 2;  //114 / 53 = 2
    16'b01110010_00110110 : OUT <= 2;  //114 / 54 = 2
    16'b01110010_00110111 : OUT <= 2;  //114 / 55 = 2
    16'b01110010_00111000 : OUT <= 2;  //114 / 56 = 2
    16'b01110010_00111001 : OUT <= 2;  //114 / 57 = 2
    16'b01110010_00111010 : OUT <= 1;  //114 / 58 = 1
    16'b01110010_00111011 : OUT <= 1;  //114 / 59 = 1
    16'b01110010_00111100 : OUT <= 1;  //114 / 60 = 1
    16'b01110010_00111101 : OUT <= 1;  //114 / 61 = 1
    16'b01110010_00111110 : OUT <= 1;  //114 / 62 = 1
    16'b01110010_00111111 : OUT <= 1;  //114 / 63 = 1
    16'b01110010_01000000 : OUT <= 1;  //114 / 64 = 1
    16'b01110010_01000001 : OUT <= 1;  //114 / 65 = 1
    16'b01110010_01000010 : OUT <= 1;  //114 / 66 = 1
    16'b01110010_01000011 : OUT <= 1;  //114 / 67 = 1
    16'b01110010_01000100 : OUT <= 1;  //114 / 68 = 1
    16'b01110010_01000101 : OUT <= 1;  //114 / 69 = 1
    16'b01110010_01000110 : OUT <= 1;  //114 / 70 = 1
    16'b01110010_01000111 : OUT <= 1;  //114 / 71 = 1
    16'b01110010_01001000 : OUT <= 1;  //114 / 72 = 1
    16'b01110010_01001001 : OUT <= 1;  //114 / 73 = 1
    16'b01110010_01001010 : OUT <= 1;  //114 / 74 = 1
    16'b01110010_01001011 : OUT <= 1;  //114 / 75 = 1
    16'b01110010_01001100 : OUT <= 1;  //114 / 76 = 1
    16'b01110010_01001101 : OUT <= 1;  //114 / 77 = 1
    16'b01110010_01001110 : OUT <= 1;  //114 / 78 = 1
    16'b01110010_01001111 : OUT <= 1;  //114 / 79 = 1
    16'b01110010_01010000 : OUT <= 1;  //114 / 80 = 1
    16'b01110010_01010001 : OUT <= 1;  //114 / 81 = 1
    16'b01110010_01010010 : OUT <= 1;  //114 / 82 = 1
    16'b01110010_01010011 : OUT <= 1;  //114 / 83 = 1
    16'b01110010_01010100 : OUT <= 1;  //114 / 84 = 1
    16'b01110010_01010101 : OUT <= 1;  //114 / 85 = 1
    16'b01110010_01010110 : OUT <= 1;  //114 / 86 = 1
    16'b01110010_01010111 : OUT <= 1;  //114 / 87 = 1
    16'b01110010_01011000 : OUT <= 1;  //114 / 88 = 1
    16'b01110010_01011001 : OUT <= 1;  //114 / 89 = 1
    16'b01110010_01011010 : OUT <= 1;  //114 / 90 = 1
    16'b01110010_01011011 : OUT <= 1;  //114 / 91 = 1
    16'b01110010_01011100 : OUT <= 1;  //114 / 92 = 1
    16'b01110010_01011101 : OUT <= 1;  //114 / 93 = 1
    16'b01110010_01011110 : OUT <= 1;  //114 / 94 = 1
    16'b01110010_01011111 : OUT <= 1;  //114 / 95 = 1
    16'b01110010_01100000 : OUT <= 1;  //114 / 96 = 1
    16'b01110010_01100001 : OUT <= 1;  //114 / 97 = 1
    16'b01110010_01100010 : OUT <= 1;  //114 / 98 = 1
    16'b01110010_01100011 : OUT <= 1;  //114 / 99 = 1
    16'b01110010_01100100 : OUT <= 1;  //114 / 100 = 1
    16'b01110010_01100101 : OUT <= 1;  //114 / 101 = 1
    16'b01110010_01100110 : OUT <= 1;  //114 / 102 = 1
    16'b01110010_01100111 : OUT <= 1;  //114 / 103 = 1
    16'b01110010_01101000 : OUT <= 1;  //114 / 104 = 1
    16'b01110010_01101001 : OUT <= 1;  //114 / 105 = 1
    16'b01110010_01101010 : OUT <= 1;  //114 / 106 = 1
    16'b01110010_01101011 : OUT <= 1;  //114 / 107 = 1
    16'b01110010_01101100 : OUT <= 1;  //114 / 108 = 1
    16'b01110010_01101101 : OUT <= 1;  //114 / 109 = 1
    16'b01110010_01101110 : OUT <= 1;  //114 / 110 = 1
    16'b01110010_01101111 : OUT <= 1;  //114 / 111 = 1
    16'b01110010_01110000 : OUT <= 1;  //114 / 112 = 1
    16'b01110010_01110001 : OUT <= 1;  //114 / 113 = 1
    16'b01110010_01110010 : OUT <= 1;  //114 / 114 = 1
    16'b01110010_01110011 : OUT <= 0;  //114 / 115 = 0
    16'b01110010_01110100 : OUT <= 0;  //114 / 116 = 0
    16'b01110010_01110101 : OUT <= 0;  //114 / 117 = 0
    16'b01110010_01110110 : OUT <= 0;  //114 / 118 = 0
    16'b01110010_01110111 : OUT <= 0;  //114 / 119 = 0
    16'b01110010_01111000 : OUT <= 0;  //114 / 120 = 0
    16'b01110010_01111001 : OUT <= 0;  //114 / 121 = 0
    16'b01110010_01111010 : OUT <= 0;  //114 / 122 = 0
    16'b01110010_01111011 : OUT <= 0;  //114 / 123 = 0
    16'b01110010_01111100 : OUT <= 0;  //114 / 124 = 0
    16'b01110010_01111101 : OUT <= 0;  //114 / 125 = 0
    16'b01110010_01111110 : OUT <= 0;  //114 / 126 = 0
    16'b01110010_01111111 : OUT <= 0;  //114 / 127 = 0
    16'b01110010_10000000 : OUT <= 0;  //114 / 128 = 0
    16'b01110010_10000001 : OUT <= 0;  //114 / 129 = 0
    16'b01110010_10000010 : OUT <= 0;  //114 / 130 = 0
    16'b01110010_10000011 : OUT <= 0;  //114 / 131 = 0
    16'b01110010_10000100 : OUT <= 0;  //114 / 132 = 0
    16'b01110010_10000101 : OUT <= 0;  //114 / 133 = 0
    16'b01110010_10000110 : OUT <= 0;  //114 / 134 = 0
    16'b01110010_10000111 : OUT <= 0;  //114 / 135 = 0
    16'b01110010_10001000 : OUT <= 0;  //114 / 136 = 0
    16'b01110010_10001001 : OUT <= 0;  //114 / 137 = 0
    16'b01110010_10001010 : OUT <= 0;  //114 / 138 = 0
    16'b01110010_10001011 : OUT <= 0;  //114 / 139 = 0
    16'b01110010_10001100 : OUT <= 0;  //114 / 140 = 0
    16'b01110010_10001101 : OUT <= 0;  //114 / 141 = 0
    16'b01110010_10001110 : OUT <= 0;  //114 / 142 = 0
    16'b01110010_10001111 : OUT <= 0;  //114 / 143 = 0
    16'b01110010_10010000 : OUT <= 0;  //114 / 144 = 0
    16'b01110010_10010001 : OUT <= 0;  //114 / 145 = 0
    16'b01110010_10010010 : OUT <= 0;  //114 / 146 = 0
    16'b01110010_10010011 : OUT <= 0;  //114 / 147 = 0
    16'b01110010_10010100 : OUT <= 0;  //114 / 148 = 0
    16'b01110010_10010101 : OUT <= 0;  //114 / 149 = 0
    16'b01110010_10010110 : OUT <= 0;  //114 / 150 = 0
    16'b01110010_10010111 : OUT <= 0;  //114 / 151 = 0
    16'b01110010_10011000 : OUT <= 0;  //114 / 152 = 0
    16'b01110010_10011001 : OUT <= 0;  //114 / 153 = 0
    16'b01110010_10011010 : OUT <= 0;  //114 / 154 = 0
    16'b01110010_10011011 : OUT <= 0;  //114 / 155 = 0
    16'b01110010_10011100 : OUT <= 0;  //114 / 156 = 0
    16'b01110010_10011101 : OUT <= 0;  //114 / 157 = 0
    16'b01110010_10011110 : OUT <= 0;  //114 / 158 = 0
    16'b01110010_10011111 : OUT <= 0;  //114 / 159 = 0
    16'b01110010_10100000 : OUT <= 0;  //114 / 160 = 0
    16'b01110010_10100001 : OUT <= 0;  //114 / 161 = 0
    16'b01110010_10100010 : OUT <= 0;  //114 / 162 = 0
    16'b01110010_10100011 : OUT <= 0;  //114 / 163 = 0
    16'b01110010_10100100 : OUT <= 0;  //114 / 164 = 0
    16'b01110010_10100101 : OUT <= 0;  //114 / 165 = 0
    16'b01110010_10100110 : OUT <= 0;  //114 / 166 = 0
    16'b01110010_10100111 : OUT <= 0;  //114 / 167 = 0
    16'b01110010_10101000 : OUT <= 0;  //114 / 168 = 0
    16'b01110010_10101001 : OUT <= 0;  //114 / 169 = 0
    16'b01110010_10101010 : OUT <= 0;  //114 / 170 = 0
    16'b01110010_10101011 : OUT <= 0;  //114 / 171 = 0
    16'b01110010_10101100 : OUT <= 0;  //114 / 172 = 0
    16'b01110010_10101101 : OUT <= 0;  //114 / 173 = 0
    16'b01110010_10101110 : OUT <= 0;  //114 / 174 = 0
    16'b01110010_10101111 : OUT <= 0;  //114 / 175 = 0
    16'b01110010_10110000 : OUT <= 0;  //114 / 176 = 0
    16'b01110010_10110001 : OUT <= 0;  //114 / 177 = 0
    16'b01110010_10110010 : OUT <= 0;  //114 / 178 = 0
    16'b01110010_10110011 : OUT <= 0;  //114 / 179 = 0
    16'b01110010_10110100 : OUT <= 0;  //114 / 180 = 0
    16'b01110010_10110101 : OUT <= 0;  //114 / 181 = 0
    16'b01110010_10110110 : OUT <= 0;  //114 / 182 = 0
    16'b01110010_10110111 : OUT <= 0;  //114 / 183 = 0
    16'b01110010_10111000 : OUT <= 0;  //114 / 184 = 0
    16'b01110010_10111001 : OUT <= 0;  //114 / 185 = 0
    16'b01110010_10111010 : OUT <= 0;  //114 / 186 = 0
    16'b01110010_10111011 : OUT <= 0;  //114 / 187 = 0
    16'b01110010_10111100 : OUT <= 0;  //114 / 188 = 0
    16'b01110010_10111101 : OUT <= 0;  //114 / 189 = 0
    16'b01110010_10111110 : OUT <= 0;  //114 / 190 = 0
    16'b01110010_10111111 : OUT <= 0;  //114 / 191 = 0
    16'b01110010_11000000 : OUT <= 0;  //114 / 192 = 0
    16'b01110010_11000001 : OUT <= 0;  //114 / 193 = 0
    16'b01110010_11000010 : OUT <= 0;  //114 / 194 = 0
    16'b01110010_11000011 : OUT <= 0;  //114 / 195 = 0
    16'b01110010_11000100 : OUT <= 0;  //114 / 196 = 0
    16'b01110010_11000101 : OUT <= 0;  //114 / 197 = 0
    16'b01110010_11000110 : OUT <= 0;  //114 / 198 = 0
    16'b01110010_11000111 : OUT <= 0;  //114 / 199 = 0
    16'b01110010_11001000 : OUT <= 0;  //114 / 200 = 0
    16'b01110010_11001001 : OUT <= 0;  //114 / 201 = 0
    16'b01110010_11001010 : OUT <= 0;  //114 / 202 = 0
    16'b01110010_11001011 : OUT <= 0;  //114 / 203 = 0
    16'b01110010_11001100 : OUT <= 0;  //114 / 204 = 0
    16'b01110010_11001101 : OUT <= 0;  //114 / 205 = 0
    16'b01110010_11001110 : OUT <= 0;  //114 / 206 = 0
    16'b01110010_11001111 : OUT <= 0;  //114 / 207 = 0
    16'b01110010_11010000 : OUT <= 0;  //114 / 208 = 0
    16'b01110010_11010001 : OUT <= 0;  //114 / 209 = 0
    16'b01110010_11010010 : OUT <= 0;  //114 / 210 = 0
    16'b01110010_11010011 : OUT <= 0;  //114 / 211 = 0
    16'b01110010_11010100 : OUT <= 0;  //114 / 212 = 0
    16'b01110010_11010101 : OUT <= 0;  //114 / 213 = 0
    16'b01110010_11010110 : OUT <= 0;  //114 / 214 = 0
    16'b01110010_11010111 : OUT <= 0;  //114 / 215 = 0
    16'b01110010_11011000 : OUT <= 0;  //114 / 216 = 0
    16'b01110010_11011001 : OUT <= 0;  //114 / 217 = 0
    16'b01110010_11011010 : OUT <= 0;  //114 / 218 = 0
    16'b01110010_11011011 : OUT <= 0;  //114 / 219 = 0
    16'b01110010_11011100 : OUT <= 0;  //114 / 220 = 0
    16'b01110010_11011101 : OUT <= 0;  //114 / 221 = 0
    16'b01110010_11011110 : OUT <= 0;  //114 / 222 = 0
    16'b01110010_11011111 : OUT <= 0;  //114 / 223 = 0
    16'b01110010_11100000 : OUT <= 0;  //114 / 224 = 0
    16'b01110010_11100001 : OUT <= 0;  //114 / 225 = 0
    16'b01110010_11100010 : OUT <= 0;  //114 / 226 = 0
    16'b01110010_11100011 : OUT <= 0;  //114 / 227 = 0
    16'b01110010_11100100 : OUT <= 0;  //114 / 228 = 0
    16'b01110010_11100101 : OUT <= 0;  //114 / 229 = 0
    16'b01110010_11100110 : OUT <= 0;  //114 / 230 = 0
    16'b01110010_11100111 : OUT <= 0;  //114 / 231 = 0
    16'b01110010_11101000 : OUT <= 0;  //114 / 232 = 0
    16'b01110010_11101001 : OUT <= 0;  //114 / 233 = 0
    16'b01110010_11101010 : OUT <= 0;  //114 / 234 = 0
    16'b01110010_11101011 : OUT <= 0;  //114 / 235 = 0
    16'b01110010_11101100 : OUT <= 0;  //114 / 236 = 0
    16'b01110010_11101101 : OUT <= 0;  //114 / 237 = 0
    16'b01110010_11101110 : OUT <= 0;  //114 / 238 = 0
    16'b01110010_11101111 : OUT <= 0;  //114 / 239 = 0
    16'b01110010_11110000 : OUT <= 0;  //114 / 240 = 0
    16'b01110010_11110001 : OUT <= 0;  //114 / 241 = 0
    16'b01110010_11110010 : OUT <= 0;  //114 / 242 = 0
    16'b01110010_11110011 : OUT <= 0;  //114 / 243 = 0
    16'b01110010_11110100 : OUT <= 0;  //114 / 244 = 0
    16'b01110010_11110101 : OUT <= 0;  //114 / 245 = 0
    16'b01110010_11110110 : OUT <= 0;  //114 / 246 = 0
    16'b01110010_11110111 : OUT <= 0;  //114 / 247 = 0
    16'b01110010_11111000 : OUT <= 0;  //114 / 248 = 0
    16'b01110010_11111001 : OUT <= 0;  //114 / 249 = 0
    16'b01110010_11111010 : OUT <= 0;  //114 / 250 = 0
    16'b01110010_11111011 : OUT <= 0;  //114 / 251 = 0
    16'b01110010_11111100 : OUT <= 0;  //114 / 252 = 0
    16'b01110010_11111101 : OUT <= 0;  //114 / 253 = 0
    16'b01110010_11111110 : OUT <= 0;  //114 / 254 = 0
    16'b01110010_11111111 : OUT <= 0;  //114 / 255 = 0
    16'b01110011_00000000 : OUT <= 0;  //115 / 0 = 0
    16'b01110011_00000001 : OUT <= 115;  //115 / 1 = 115
    16'b01110011_00000010 : OUT <= 57;  //115 / 2 = 57
    16'b01110011_00000011 : OUT <= 38;  //115 / 3 = 38
    16'b01110011_00000100 : OUT <= 28;  //115 / 4 = 28
    16'b01110011_00000101 : OUT <= 23;  //115 / 5 = 23
    16'b01110011_00000110 : OUT <= 19;  //115 / 6 = 19
    16'b01110011_00000111 : OUT <= 16;  //115 / 7 = 16
    16'b01110011_00001000 : OUT <= 14;  //115 / 8 = 14
    16'b01110011_00001001 : OUT <= 12;  //115 / 9 = 12
    16'b01110011_00001010 : OUT <= 11;  //115 / 10 = 11
    16'b01110011_00001011 : OUT <= 10;  //115 / 11 = 10
    16'b01110011_00001100 : OUT <= 9;  //115 / 12 = 9
    16'b01110011_00001101 : OUT <= 8;  //115 / 13 = 8
    16'b01110011_00001110 : OUT <= 8;  //115 / 14 = 8
    16'b01110011_00001111 : OUT <= 7;  //115 / 15 = 7
    16'b01110011_00010000 : OUT <= 7;  //115 / 16 = 7
    16'b01110011_00010001 : OUT <= 6;  //115 / 17 = 6
    16'b01110011_00010010 : OUT <= 6;  //115 / 18 = 6
    16'b01110011_00010011 : OUT <= 6;  //115 / 19 = 6
    16'b01110011_00010100 : OUT <= 5;  //115 / 20 = 5
    16'b01110011_00010101 : OUT <= 5;  //115 / 21 = 5
    16'b01110011_00010110 : OUT <= 5;  //115 / 22 = 5
    16'b01110011_00010111 : OUT <= 5;  //115 / 23 = 5
    16'b01110011_00011000 : OUT <= 4;  //115 / 24 = 4
    16'b01110011_00011001 : OUT <= 4;  //115 / 25 = 4
    16'b01110011_00011010 : OUT <= 4;  //115 / 26 = 4
    16'b01110011_00011011 : OUT <= 4;  //115 / 27 = 4
    16'b01110011_00011100 : OUT <= 4;  //115 / 28 = 4
    16'b01110011_00011101 : OUT <= 3;  //115 / 29 = 3
    16'b01110011_00011110 : OUT <= 3;  //115 / 30 = 3
    16'b01110011_00011111 : OUT <= 3;  //115 / 31 = 3
    16'b01110011_00100000 : OUT <= 3;  //115 / 32 = 3
    16'b01110011_00100001 : OUT <= 3;  //115 / 33 = 3
    16'b01110011_00100010 : OUT <= 3;  //115 / 34 = 3
    16'b01110011_00100011 : OUT <= 3;  //115 / 35 = 3
    16'b01110011_00100100 : OUT <= 3;  //115 / 36 = 3
    16'b01110011_00100101 : OUT <= 3;  //115 / 37 = 3
    16'b01110011_00100110 : OUT <= 3;  //115 / 38 = 3
    16'b01110011_00100111 : OUT <= 2;  //115 / 39 = 2
    16'b01110011_00101000 : OUT <= 2;  //115 / 40 = 2
    16'b01110011_00101001 : OUT <= 2;  //115 / 41 = 2
    16'b01110011_00101010 : OUT <= 2;  //115 / 42 = 2
    16'b01110011_00101011 : OUT <= 2;  //115 / 43 = 2
    16'b01110011_00101100 : OUT <= 2;  //115 / 44 = 2
    16'b01110011_00101101 : OUT <= 2;  //115 / 45 = 2
    16'b01110011_00101110 : OUT <= 2;  //115 / 46 = 2
    16'b01110011_00101111 : OUT <= 2;  //115 / 47 = 2
    16'b01110011_00110000 : OUT <= 2;  //115 / 48 = 2
    16'b01110011_00110001 : OUT <= 2;  //115 / 49 = 2
    16'b01110011_00110010 : OUT <= 2;  //115 / 50 = 2
    16'b01110011_00110011 : OUT <= 2;  //115 / 51 = 2
    16'b01110011_00110100 : OUT <= 2;  //115 / 52 = 2
    16'b01110011_00110101 : OUT <= 2;  //115 / 53 = 2
    16'b01110011_00110110 : OUT <= 2;  //115 / 54 = 2
    16'b01110011_00110111 : OUT <= 2;  //115 / 55 = 2
    16'b01110011_00111000 : OUT <= 2;  //115 / 56 = 2
    16'b01110011_00111001 : OUT <= 2;  //115 / 57 = 2
    16'b01110011_00111010 : OUT <= 1;  //115 / 58 = 1
    16'b01110011_00111011 : OUT <= 1;  //115 / 59 = 1
    16'b01110011_00111100 : OUT <= 1;  //115 / 60 = 1
    16'b01110011_00111101 : OUT <= 1;  //115 / 61 = 1
    16'b01110011_00111110 : OUT <= 1;  //115 / 62 = 1
    16'b01110011_00111111 : OUT <= 1;  //115 / 63 = 1
    16'b01110011_01000000 : OUT <= 1;  //115 / 64 = 1
    16'b01110011_01000001 : OUT <= 1;  //115 / 65 = 1
    16'b01110011_01000010 : OUT <= 1;  //115 / 66 = 1
    16'b01110011_01000011 : OUT <= 1;  //115 / 67 = 1
    16'b01110011_01000100 : OUT <= 1;  //115 / 68 = 1
    16'b01110011_01000101 : OUT <= 1;  //115 / 69 = 1
    16'b01110011_01000110 : OUT <= 1;  //115 / 70 = 1
    16'b01110011_01000111 : OUT <= 1;  //115 / 71 = 1
    16'b01110011_01001000 : OUT <= 1;  //115 / 72 = 1
    16'b01110011_01001001 : OUT <= 1;  //115 / 73 = 1
    16'b01110011_01001010 : OUT <= 1;  //115 / 74 = 1
    16'b01110011_01001011 : OUT <= 1;  //115 / 75 = 1
    16'b01110011_01001100 : OUT <= 1;  //115 / 76 = 1
    16'b01110011_01001101 : OUT <= 1;  //115 / 77 = 1
    16'b01110011_01001110 : OUT <= 1;  //115 / 78 = 1
    16'b01110011_01001111 : OUT <= 1;  //115 / 79 = 1
    16'b01110011_01010000 : OUT <= 1;  //115 / 80 = 1
    16'b01110011_01010001 : OUT <= 1;  //115 / 81 = 1
    16'b01110011_01010010 : OUT <= 1;  //115 / 82 = 1
    16'b01110011_01010011 : OUT <= 1;  //115 / 83 = 1
    16'b01110011_01010100 : OUT <= 1;  //115 / 84 = 1
    16'b01110011_01010101 : OUT <= 1;  //115 / 85 = 1
    16'b01110011_01010110 : OUT <= 1;  //115 / 86 = 1
    16'b01110011_01010111 : OUT <= 1;  //115 / 87 = 1
    16'b01110011_01011000 : OUT <= 1;  //115 / 88 = 1
    16'b01110011_01011001 : OUT <= 1;  //115 / 89 = 1
    16'b01110011_01011010 : OUT <= 1;  //115 / 90 = 1
    16'b01110011_01011011 : OUT <= 1;  //115 / 91 = 1
    16'b01110011_01011100 : OUT <= 1;  //115 / 92 = 1
    16'b01110011_01011101 : OUT <= 1;  //115 / 93 = 1
    16'b01110011_01011110 : OUT <= 1;  //115 / 94 = 1
    16'b01110011_01011111 : OUT <= 1;  //115 / 95 = 1
    16'b01110011_01100000 : OUT <= 1;  //115 / 96 = 1
    16'b01110011_01100001 : OUT <= 1;  //115 / 97 = 1
    16'b01110011_01100010 : OUT <= 1;  //115 / 98 = 1
    16'b01110011_01100011 : OUT <= 1;  //115 / 99 = 1
    16'b01110011_01100100 : OUT <= 1;  //115 / 100 = 1
    16'b01110011_01100101 : OUT <= 1;  //115 / 101 = 1
    16'b01110011_01100110 : OUT <= 1;  //115 / 102 = 1
    16'b01110011_01100111 : OUT <= 1;  //115 / 103 = 1
    16'b01110011_01101000 : OUT <= 1;  //115 / 104 = 1
    16'b01110011_01101001 : OUT <= 1;  //115 / 105 = 1
    16'b01110011_01101010 : OUT <= 1;  //115 / 106 = 1
    16'b01110011_01101011 : OUT <= 1;  //115 / 107 = 1
    16'b01110011_01101100 : OUT <= 1;  //115 / 108 = 1
    16'b01110011_01101101 : OUT <= 1;  //115 / 109 = 1
    16'b01110011_01101110 : OUT <= 1;  //115 / 110 = 1
    16'b01110011_01101111 : OUT <= 1;  //115 / 111 = 1
    16'b01110011_01110000 : OUT <= 1;  //115 / 112 = 1
    16'b01110011_01110001 : OUT <= 1;  //115 / 113 = 1
    16'b01110011_01110010 : OUT <= 1;  //115 / 114 = 1
    16'b01110011_01110011 : OUT <= 1;  //115 / 115 = 1
    16'b01110011_01110100 : OUT <= 0;  //115 / 116 = 0
    16'b01110011_01110101 : OUT <= 0;  //115 / 117 = 0
    16'b01110011_01110110 : OUT <= 0;  //115 / 118 = 0
    16'b01110011_01110111 : OUT <= 0;  //115 / 119 = 0
    16'b01110011_01111000 : OUT <= 0;  //115 / 120 = 0
    16'b01110011_01111001 : OUT <= 0;  //115 / 121 = 0
    16'b01110011_01111010 : OUT <= 0;  //115 / 122 = 0
    16'b01110011_01111011 : OUT <= 0;  //115 / 123 = 0
    16'b01110011_01111100 : OUT <= 0;  //115 / 124 = 0
    16'b01110011_01111101 : OUT <= 0;  //115 / 125 = 0
    16'b01110011_01111110 : OUT <= 0;  //115 / 126 = 0
    16'b01110011_01111111 : OUT <= 0;  //115 / 127 = 0
    16'b01110011_10000000 : OUT <= 0;  //115 / 128 = 0
    16'b01110011_10000001 : OUT <= 0;  //115 / 129 = 0
    16'b01110011_10000010 : OUT <= 0;  //115 / 130 = 0
    16'b01110011_10000011 : OUT <= 0;  //115 / 131 = 0
    16'b01110011_10000100 : OUT <= 0;  //115 / 132 = 0
    16'b01110011_10000101 : OUT <= 0;  //115 / 133 = 0
    16'b01110011_10000110 : OUT <= 0;  //115 / 134 = 0
    16'b01110011_10000111 : OUT <= 0;  //115 / 135 = 0
    16'b01110011_10001000 : OUT <= 0;  //115 / 136 = 0
    16'b01110011_10001001 : OUT <= 0;  //115 / 137 = 0
    16'b01110011_10001010 : OUT <= 0;  //115 / 138 = 0
    16'b01110011_10001011 : OUT <= 0;  //115 / 139 = 0
    16'b01110011_10001100 : OUT <= 0;  //115 / 140 = 0
    16'b01110011_10001101 : OUT <= 0;  //115 / 141 = 0
    16'b01110011_10001110 : OUT <= 0;  //115 / 142 = 0
    16'b01110011_10001111 : OUT <= 0;  //115 / 143 = 0
    16'b01110011_10010000 : OUT <= 0;  //115 / 144 = 0
    16'b01110011_10010001 : OUT <= 0;  //115 / 145 = 0
    16'b01110011_10010010 : OUT <= 0;  //115 / 146 = 0
    16'b01110011_10010011 : OUT <= 0;  //115 / 147 = 0
    16'b01110011_10010100 : OUT <= 0;  //115 / 148 = 0
    16'b01110011_10010101 : OUT <= 0;  //115 / 149 = 0
    16'b01110011_10010110 : OUT <= 0;  //115 / 150 = 0
    16'b01110011_10010111 : OUT <= 0;  //115 / 151 = 0
    16'b01110011_10011000 : OUT <= 0;  //115 / 152 = 0
    16'b01110011_10011001 : OUT <= 0;  //115 / 153 = 0
    16'b01110011_10011010 : OUT <= 0;  //115 / 154 = 0
    16'b01110011_10011011 : OUT <= 0;  //115 / 155 = 0
    16'b01110011_10011100 : OUT <= 0;  //115 / 156 = 0
    16'b01110011_10011101 : OUT <= 0;  //115 / 157 = 0
    16'b01110011_10011110 : OUT <= 0;  //115 / 158 = 0
    16'b01110011_10011111 : OUT <= 0;  //115 / 159 = 0
    16'b01110011_10100000 : OUT <= 0;  //115 / 160 = 0
    16'b01110011_10100001 : OUT <= 0;  //115 / 161 = 0
    16'b01110011_10100010 : OUT <= 0;  //115 / 162 = 0
    16'b01110011_10100011 : OUT <= 0;  //115 / 163 = 0
    16'b01110011_10100100 : OUT <= 0;  //115 / 164 = 0
    16'b01110011_10100101 : OUT <= 0;  //115 / 165 = 0
    16'b01110011_10100110 : OUT <= 0;  //115 / 166 = 0
    16'b01110011_10100111 : OUT <= 0;  //115 / 167 = 0
    16'b01110011_10101000 : OUT <= 0;  //115 / 168 = 0
    16'b01110011_10101001 : OUT <= 0;  //115 / 169 = 0
    16'b01110011_10101010 : OUT <= 0;  //115 / 170 = 0
    16'b01110011_10101011 : OUT <= 0;  //115 / 171 = 0
    16'b01110011_10101100 : OUT <= 0;  //115 / 172 = 0
    16'b01110011_10101101 : OUT <= 0;  //115 / 173 = 0
    16'b01110011_10101110 : OUT <= 0;  //115 / 174 = 0
    16'b01110011_10101111 : OUT <= 0;  //115 / 175 = 0
    16'b01110011_10110000 : OUT <= 0;  //115 / 176 = 0
    16'b01110011_10110001 : OUT <= 0;  //115 / 177 = 0
    16'b01110011_10110010 : OUT <= 0;  //115 / 178 = 0
    16'b01110011_10110011 : OUT <= 0;  //115 / 179 = 0
    16'b01110011_10110100 : OUT <= 0;  //115 / 180 = 0
    16'b01110011_10110101 : OUT <= 0;  //115 / 181 = 0
    16'b01110011_10110110 : OUT <= 0;  //115 / 182 = 0
    16'b01110011_10110111 : OUT <= 0;  //115 / 183 = 0
    16'b01110011_10111000 : OUT <= 0;  //115 / 184 = 0
    16'b01110011_10111001 : OUT <= 0;  //115 / 185 = 0
    16'b01110011_10111010 : OUT <= 0;  //115 / 186 = 0
    16'b01110011_10111011 : OUT <= 0;  //115 / 187 = 0
    16'b01110011_10111100 : OUT <= 0;  //115 / 188 = 0
    16'b01110011_10111101 : OUT <= 0;  //115 / 189 = 0
    16'b01110011_10111110 : OUT <= 0;  //115 / 190 = 0
    16'b01110011_10111111 : OUT <= 0;  //115 / 191 = 0
    16'b01110011_11000000 : OUT <= 0;  //115 / 192 = 0
    16'b01110011_11000001 : OUT <= 0;  //115 / 193 = 0
    16'b01110011_11000010 : OUT <= 0;  //115 / 194 = 0
    16'b01110011_11000011 : OUT <= 0;  //115 / 195 = 0
    16'b01110011_11000100 : OUT <= 0;  //115 / 196 = 0
    16'b01110011_11000101 : OUT <= 0;  //115 / 197 = 0
    16'b01110011_11000110 : OUT <= 0;  //115 / 198 = 0
    16'b01110011_11000111 : OUT <= 0;  //115 / 199 = 0
    16'b01110011_11001000 : OUT <= 0;  //115 / 200 = 0
    16'b01110011_11001001 : OUT <= 0;  //115 / 201 = 0
    16'b01110011_11001010 : OUT <= 0;  //115 / 202 = 0
    16'b01110011_11001011 : OUT <= 0;  //115 / 203 = 0
    16'b01110011_11001100 : OUT <= 0;  //115 / 204 = 0
    16'b01110011_11001101 : OUT <= 0;  //115 / 205 = 0
    16'b01110011_11001110 : OUT <= 0;  //115 / 206 = 0
    16'b01110011_11001111 : OUT <= 0;  //115 / 207 = 0
    16'b01110011_11010000 : OUT <= 0;  //115 / 208 = 0
    16'b01110011_11010001 : OUT <= 0;  //115 / 209 = 0
    16'b01110011_11010010 : OUT <= 0;  //115 / 210 = 0
    16'b01110011_11010011 : OUT <= 0;  //115 / 211 = 0
    16'b01110011_11010100 : OUT <= 0;  //115 / 212 = 0
    16'b01110011_11010101 : OUT <= 0;  //115 / 213 = 0
    16'b01110011_11010110 : OUT <= 0;  //115 / 214 = 0
    16'b01110011_11010111 : OUT <= 0;  //115 / 215 = 0
    16'b01110011_11011000 : OUT <= 0;  //115 / 216 = 0
    16'b01110011_11011001 : OUT <= 0;  //115 / 217 = 0
    16'b01110011_11011010 : OUT <= 0;  //115 / 218 = 0
    16'b01110011_11011011 : OUT <= 0;  //115 / 219 = 0
    16'b01110011_11011100 : OUT <= 0;  //115 / 220 = 0
    16'b01110011_11011101 : OUT <= 0;  //115 / 221 = 0
    16'b01110011_11011110 : OUT <= 0;  //115 / 222 = 0
    16'b01110011_11011111 : OUT <= 0;  //115 / 223 = 0
    16'b01110011_11100000 : OUT <= 0;  //115 / 224 = 0
    16'b01110011_11100001 : OUT <= 0;  //115 / 225 = 0
    16'b01110011_11100010 : OUT <= 0;  //115 / 226 = 0
    16'b01110011_11100011 : OUT <= 0;  //115 / 227 = 0
    16'b01110011_11100100 : OUT <= 0;  //115 / 228 = 0
    16'b01110011_11100101 : OUT <= 0;  //115 / 229 = 0
    16'b01110011_11100110 : OUT <= 0;  //115 / 230 = 0
    16'b01110011_11100111 : OUT <= 0;  //115 / 231 = 0
    16'b01110011_11101000 : OUT <= 0;  //115 / 232 = 0
    16'b01110011_11101001 : OUT <= 0;  //115 / 233 = 0
    16'b01110011_11101010 : OUT <= 0;  //115 / 234 = 0
    16'b01110011_11101011 : OUT <= 0;  //115 / 235 = 0
    16'b01110011_11101100 : OUT <= 0;  //115 / 236 = 0
    16'b01110011_11101101 : OUT <= 0;  //115 / 237 = 0
    16'b01110011_11101110 : OUT <= 0;  //115 / 238 = 0
    16'b01110011_11101111 : OUT <= 0;  //115 / 239 = 0
    16'b01110011_11110000 : OUT <= 0;  //115 / 240 = 0
    16'b01110011_11110001 : OUT <= 0;  //115 / 241 = 0
    16'b01110011_11110010 : OUT <= 0;  //115 / 242 = 0
    16'b01110011_11110011 : OUT <= 0;  //115 / 243 = 0
    16'b01110011_11110100 : OUT <= 0;  //115 / 244 = 0
    16'b01110011_11110101 : OUT <= 0;  //115 / 245 = 0
    16'b01110011_11110110 : OUT <= 0;  //115 / 246 = 0
    16'b01110011_11110111 : OUT <= 0;  //115 / 247 = 0
    16'b01110011_11111000 : OUT <= 0;  //115 / 248 = 0
    16'b01110011_11111001 : OUT <= 0;  //115 / 249 = 0
    16'b01110011_11111010 : OUT <= 0;  //115 / 250 = 0
    16'b01110011_11111011 : OUT <= 0;  //115 / 251 = 0
    16'b01110011_11111100 : OUT <= 0;  //115 / 252 = 0
    16'b01110011_11111101 : OUT <= 0;  //115 / 253 = 0
    16'b01110011_11111110 : OUT <= 0;  //115 / 254 = 0
    16'b01110011_11111111 : OUT <= 0;  //115 / 255 = 0
    16'b01110100_00000000 : OUT <= 0;  //116 / 0 = 0
    16'b01110100_00000001 : OUT <= 116;  //116 / 1 = 116
    16'b01110100_00000010 : OUT <= 58;  //116 / 2 = 58
    16'b01110100_00000011 : OUT <= 38;  //116 / 3 = 38
    16'b01110100_00000100 : OUT <= 29;  //116 / 4 = 29
    16'b01110100_00000101 : OUT <= 23;  //116 / 5 = 23
    16'b01110100_00000110 : OUT <= 19;  //116 / 6 = 19
    16'b01110100_00000111 : OUT <= 16;  //116 / 7 = 16
    16'b01110100_00001000 : OUT <= 14;  //116 / 8 = 14
    16'b01110100_00001001 : OUT <= 12;  //116 / 9 = 12
    16'b01110100_00001010 : OUT <= 11;  //116 / 10 = 11
    16'b01110100_00001011 : OUT <= 10;  //116 / 11 = 10
    16'b01110100_00001100 : OUT <= 9;  //116 / 12 = 9
    16'b01110100_00001101 : OUT <= 8;  //116 / 13 = 8
    16'b01110100_00001110 : OUT <= 8;  //116 / 14 = 8
    16'b01110100_00001111 : OUT <= 7;  //116 / 15 = 7
    16'b01110100_00010000 : OUT <= 7;  //116 / 16 = 7
    16'b01110100_00010001 : OUT <= 6;  //116 / 17 = 6
    16'b01110100_00010010 : OUT <= 6;  //116 / 18 = 6
    16'b01110100_00010011 : OUT <= 6;  //116 / 19 = 6
    16'b01110100_00010100 : OUT <= 5;  //116 / 20 = 5
    16'b01110100_00010101 : OUT <= 5;  //116 / 21 = 5
    16'b01110100_00010110 : OUT <= 5;  //116 / 22 = 5
    16'b01110100_00010111 : OUT <= 5;  //116 / 23 = 5
    16'b01110100_00011000 : OUT <= 4;  //116 / 24 = 4
    16'b01110100_00011001 : OUT <= 4;  //116 / 25 = 4
    16'b01110100_00011010 : OUT <= 4;  //116 / 26 = 4
    16'b01110100_00011011 : OUT <= 4;  //116 / 27 = 4
    16'b01110100_00011100 : OUT <= 4;  //116 / 28 = 4
    16'b01110100_00011101 : OUT <= 4;  //116 / 29 = 4
    16'b01110100_00011110 : OUT <= 3;  //116 / 30 = 3
    16'b01110100_00011111 : OUT <= 3;  //116 / 31 = 3
    16'b01110100_00100000 : OUT <= 3;  //116 / 32 = 3
    16'b01110100_00100001 : OUT <= 3;  //116 / 33 = 3
    16'b01110100_00100010 : OUT <= 3;  //116 / 34 = 3
    16'b01110100_00100011 : OUT <= 3;  //116 / 35 = 3
    16'b01110100_00100100 : OUT <= 3;  //116 / 36 = 3
    16'b01110100_00100101 : OUT <= 3;  //116 / 37 = 3
    16'b01110100_00100110 : OUT <= 3;  //116 / 38 = 3
    16'b01110100_00100111 : OUT <= 2;  //116 / 39 = 2
    16'b01110100_00101000 : OUT <= 2;  //116 / 40 = 2
    16'b01110100_00101001 : OUT <= 2;  //116 / 41 = 2
    16'b01110100_00101010 : OUT <= 2;  //116 / 42 = 2
    16'b01110100_00101011 : OUT <= 2;  //116 / 43 = 2
    16'b01110100_00101100 : OUT <= 2;  //116 / 44 = 2
    16'b01110100_00101101 : OUT <= 2;  //116 / 45 = 2
    16'b01110100_00101110 : OUT <= 2;  //116 / 46 = 2
    16'b01110100_00101111 : OUT <= 2;  //116 / 47 = 2
    16'b01110100_00110000 : OUT <= 2;  //116 / 48 = 2
    16'b01110100_00110001 : OUT <= 2;  //116 / 49 = 2
    16'b01110100_00110010 : OUT <= 2;  //116 / 50 = 2
    16'b01110100_00110011 : OUT <= 2;  //116 / 51 = 2
    16'b01110100_00110100 : OUT <= 2;  //116 / 52 = 2
    16'b01110100_00110101 : OUT <= 2;  //116 / 53 = 2
    16'b01110100_00110110 : OUT <= 2;  //116 / 54 = 2
    16'b01110100_00110111 : OUT <= 2;  //116 / 55 = 2
    16'b01110100_00111000 : OUT <= 2;  //116 / 56 = 2
    16'b01110100_00111001 : OUT <= 2;  //116 / 57 = 2
    16'b01110100_00111010 : OUT <= 2;  //116 / 58 = 2
    16'b01110100_00111011 : OUT <= 1;  //116 / 59 = 1
    16'b01110100_00111100 : OUT <= 1;  //116 / 60 = 1
    16'b01110100_00111101 : OUT <= 1;  //116 / 61 = 1
    16'b01110100_00111110 : OUT <= 1;  //116 / 62 = 1
    16'b01110100_00111111 : OUT <= 1;  //116 / 63 = 1
    16'b01110100_01000000 : OUT <= 1;  //116 / 64 = 1
    16'b01110100_01000001 : OUT <= 1;  //116 / 65 = 1
    16'b01110100_01000010 : OUT <= 1;  //116 / 66 = 1
    16'b01110100_01000011 : OUT <= 1;  //116 / 67 = 1
    16'b01110100_01000100 : OUT <= 1;  //116 / 68 = 1
    16'b01110100_01000101 : OUT <= 1;  //116 / 69 = 1
    16'b01110100_01000110 : OUT <= 1;  //116 / 70 = 1
    16'b01110100_01000111 : OUT <= 1;  //116 / 71 = 1
    16'b01110100_01001000 : OUT <= 1;  //116 / 72 = 1
    16'b01110100_01001001 : OUT <= 1;  //116 / 73 = 1
    16'b01110100_01001010 : OUT <= 1;  //116 / 74 = 1
    16'b01110100_01001011 : OUT <= 1;  //116 / 75 = 1
    16'b01110100_01001100 : OUT <= 1;  //116 / 76 = 1
    16'b01110100_01001101 : OUT <= 1;  //116 / 77 = 1
    16'b01110100_01001110 : OUT <= 1;  //116 / 78 = 1
    16'b01110100_01001111 : OUT <= 1;  //116 / 79 = 1
    16'b01110100_01010000 : OUT <= 1;  //116 / 80 = 1
    16'b01110100_01010001 : OUT <= 1;  //116 / 81 = 1
    16'b01110100_01010010 : OUT <= 1;  //116 / 82 = 1
    16'b01110100_01010011 : OUT <= 1;  //116 / 83 = 1
    16'b01110100_01010100 : OUT <= 1;  //116 / 84 = 1
    16'b01110100_01010101 : OUT <= 1;  //116 / 85 = 1
    16'b01110100_01010110 : OUT <= 1;  //116 / 86 = 1
    16'b01110100_01010111 : OUT <= 1;  //116 / 87 = 1
    16'b01110100_01011000 : OUT <= 1;  //116 / 88 = 1
    16'b01110100_01011001 : OUT <= 1;  //116 / 89 = 1
    16'b01110100_01011010 : OUT <= 1;  //116 / 90 = 1
    16'b01110100_01011011 : OUT <= 1;  //116 / 91 = 1
    16'b01110100_01011100 : OUT <= 1;  //116 / 92 = 1
    16'b01110100_01011101 : OUT <= 1;  //116 / 93 = 1
    16'b01110100_01011110 : OUT <= 1;  //116 / 94 = 1
    16'b01110100_01011111 : OUT <= 1;  //116 / 95 = 1
    16'b01110100_01100000 : OUT <= 1;  //116 / 96 = 1
    16'b01110100_01100001 : OUT <= 1;  //116 / 97 = 1
    16'b01110100_01100010 : OUT <= 1;  //116 / 98 = 1
    16'b01110100_01100011 : OUT <= 1;  //116 / 99 = 1
    16'b01110100_01100100 : OUT <= 1;  //116 / 100 = 1
    16'b01110100_01100101 : OUT <= 1;  //116 / 101 = 1
    16'b01110100_01100110 : OUT <= 1;  //116 / 102 = 1
    16'b01110100_01100111 : OUT <= 1;  //116 / 103 = 1
    16'b01110100_01101000 : OUT <= 1;  //116 / 104 = 1
    16'b01110100_01101001 : OUT <= 1;  //116 / 105 = 1
    16'b01110100_01101010 : OUT <= 1;  //116 / 106 = 1
    16'b01110100_01101011 : OUT <= 1;  //116 / 107 = 1
    16'b01110100_01101100 : OUT <= 1;  //116 / 108 = 1
    16'b01110100_01101101 : OUT <= 1;  //116 / 109 = 1
    16'b01110100_01101110 : OUT <= 1;  //116 / 110 = 1
    16'b01110100_01101111 : OUT <= 1;  //116 / 111 = 1
    16'b01110100_01110000 : OUT <= 1;  //116 / 112 = 1
    16'b01110100_01110001 : OUT <= 1;  //116 / 113 = 1
    16'b01110100_01110010 : OUT <= 1;  //116 / 114 = 1
    16'b01110100_01110011 : OUT <= 1;  //116 / 115 = 1
    16'b01110100_01110100 : OUT <= 1;  //116 / 116 = 1
    16'b01110100_01110101 : OUT <= 0;  //116 / 117 = 0
    16'b01110100_01110110 : OUT <= 0;  //116 / 118 = 0
    16'b01110100_01110111 : OUT <= 0;  //116 / 119 = 0
    16'b01110100_01111000 : OUT <= 0;  //116 / 120 = 0
    16'b01110100_01111001 : OUT <= 0;  //116 / 121 = 0
    16'b01110100_01111010 : OUT <= 0;  //116 / 122 = 0
    16'b01110100_01111011 : OUT <= 0;  //116 / 123 = 0
    16'b01110100_01111100 : OUT <= 0;  //116 / 124 = 0
    16'b01110100_01111101 : OUT <= 0;  //116 / 125 = 0
    16'b01110100_01111110 : OUT <= 0;  //116 / 126 = 0
    16'b01110100_01111111 : OUT <= 0;  //116 / 127 = 0
    16'b01110100_10000000 : OUT <= 0;  //116 / 128 = 0
    16'b01110100_10000001 : OUT <= 0;  //116 / 129 = 0
    16'b01110100_10000010 : OUT <= 0;  //116 / 130 = 0
    16'b01110100_10000011 : OUT <= 0;  //116 / 131 = 0
    16'b01110100_10000100 : OUT <= 0;  //116 / 132 = 0
    16'b01110100_10000101 : OUT <= 0;  //116 / 133 = 0
    16'b01110100_10000110 : OUT <= 0;  //116 / 134 = 0
    16'b01110100_10000111 : OUT <= 0;  //116 / 135 = 0
    16'b01110100_10001000 : OUT <= 0;  //116 / 136 = 0
    16'b01110100_10001001 : OUT <= 0;  //116 / 137 = 0
    16'b01110100_10001010 : OUT <= 0;  //116 / 138 = 0
    16'b01110100_10001011 : OUT <= 0;  //116 / 139 = 0
    16'b01110100_10001100 : OUT <= 0;  //116 / 140 = 0
    16'b01110100_10001101 : OUT <= 0;  //116 / 141 = 0
    16'b01110100_10001110 : OUT <= 0;  //116 / 142 = 0
    16'b01110100_10001111 : OUT <= 0;  //116 / 143 = 0
    16'b01110100_10010000 : OUT <= 0;  //116 / 144 = 0
    16'b01110100_10010001 : OUT <= 0;  //116 / 145 = 0
    16'b01110100_10010010 : OUT <= 0;  //116 / 146 = 0
    16'b01110100_10010011 : OUT <= 0;  //116 / 147 = 0
    16'b01110100_10010100 : OUT <= 0;  //116 / 148 = 0
    16'b01110100_10010101 : OUT <= 0;  //116 / 149 = 0
    16'b01110100_10010110 : OUT <= 0;  //116 / 150 = 0
    16'b01110100_10010111 : OUT <= 0;  //116 / 151 = 0
    16'b01110100_10011000 : OUT <= 0;  //116 / 152 = 0
    16'b01110100_10011001 : OUT <= 0;  //116 / 153 = 0
    16'b01110100_10011010 : OUT <= 0;  //116 / 154 = 0
    16'b01110100_10011011 : OUT <= 0;  //116 / 155 = 0
    16'b01110100_10011100 : OUT <= 0;  //116 / 156 = 0
    16'b01110100_10011101 : OUT <= 0;  //116 / 157 = 0
    16'b01110100_10011110 : OUT <= 0;  //116 / 158 = 0
    16'b01110100_10011111 : OUT <= 0;  //116 / 159 = 0
    16'b01110100_10100000 : OUT <= 0;  //116 / 160 = 0
    16'b01110100_10100001 : OUT <= 0;  //116 / 161 = 0
    16'b01110100_10100010 : OUT <= 0;  //116 / 162 = 0
    16'b01110100_10100011 : OUT <= 0;  //116 / 163 = 0
    16'b01110100_10100100 : OUT <= 0;  //116 / 164 = 0
    16'b01110100_10100101 : OUT <= 0;  //116 / 165 = 0
    16'b01110100_10100110 : OUT <= 0;  //116 / 166 = 0
    16'b01110100_10100111 : OUT <= 0;  //116 / 167 = 0
    16'b01110100_10101000 : OUT <= 0;  //116 / 168 = 0
    16'b01110100_10101001 : OUT <= 0;  //116 / 169 = 0
    16'b01110100_10101010 : OUT <= 0;  //116 / 170 = 0
    16'b01110100_10101011 : OUT <= 0;  //116 / 171 = 0
    16'b01110100_10101100 : OUT <= 0;  //116 / 172 = 0
    16'b01110100_10101101 : OUT <= 0;  //116 / 173 = 0
    16'b01110100_10101110 : OUT <= 0;  //116 / 174 = 0
    16'b01110100_10101111 : OUT <= 0;  //116 / 175 = 0
    16'b01110100_10110000 : OUT <= 0;  //116 / 176 = 0
    16'b01110100_10110001 : OUT <= 0;  //116 / 177 = 0
    16'b01110100_10110010 : OUT <= 0;  //116 / 178 = 0
    16'b01110100_10110011 : OUT <= 0;  //116 / 179 = 0
    16'b01110100_10110100 : OUT <= 0;  //116 / 180 = 0
    16'b01110100_10110101 : OUT <= 0;  //116 / 181 = 0
    16'b01110100_10110110 : OUT <= 0;  //116 / 182 = 0
    16'b01110100_10110111 : OUT <= 0;  //116 / 183 = 0
    16'b01110100_10111000 : OUT <= 0;  //116 / 184 = 0
    16'b01110100_10111001 : OUT <= 0;  //116 / 185 = 0
    16'b01110100_10111010 : OUT <= 0;  //116 / 186 = 0
    16'b01110100_10111011 : OUT <= 0;  //116 / 187 = 0
    16'b01110100_10111100 : OUT <= 0;  //116 / 188 = 0
    16'b01110100_10111101 : OUT <= 0;  //116 / 189 = 0
    16'b01110100_10111110 : OUT <= 0;  //116 / 190 = 0
    16'b01110100_10111111 : OUT <= 0;  //116 / 191 = 0
    16'b01110100_11000000 : OUT <= 0;  //116 / 192 = 0
    16'b01110100_11000001 : OUT <= 0;  //116 / 193 = 0
    16'b01110100_11000010 : OUT <= 0;  //116 / 194 = 0
    16'b01110100_11000011 : OUT <= 0;  //116 / 195 = 0
    16'b01110100_11000100 : OUT <= 0;  //116 / 196 = 0
    16'b01110100_11000101 : OUT <= 0;  //116 / 197 = 0
    16'b01110100_11000110 : OUT <= 0;  //116 / 198 = 0
    16'b01110100_11000111 : OUT <= 0;  //116 / 199 = 0
    16'b01110100_11001000 : OUT <= 0;  //116 / 200 = 0
    16'b01110100_11001001 : OUT <= 0;  //116 / 201 = 0
    16'b01110100_11001010 : OUT <= 0;  //116 / 202 = 0
    16'b01110100_11001011 : OUT <= 0;  //116 / 203 = 0
    16'b01110100_11001100 : OUT <= 0;  //116 / 204 = 0
    16'b01110100_11001101 : OUT <= 0;  //116 / 205 = 0
    16'b01110100_11001110 : OUT <= 0;  //116 / 206 = 0
    16'b01110100_11001111 : OUT <= 0;  //116 / 207 = 0
    16'b01110100_11010000 : OUT <= 0;  //116 / 208 = 0
    16'b01110100_11010001 : OUT <= 0;  //116 / 209 = 0
    16'b01110100_11010010 : OUT <= 0;  //116 / 210 = 0
    16'b01110100_11010011 : OUT <= 0;  //116 / 211 = 0
    16'b01110100_11010100 : OUT <= 0;  //116 / 212 = 0
    16'b01110100_11010101 : OUT <= 0;  //116 / 213 = 0
    16'b01110100_11010110 : OUT <= 0;  //116 / 214 = 0
    16'b01110100_11010111 : OUT <= 0;  //116 / 215 = 0
    16'b01110100_11011000 : OUT <= 0;  //116 / 216 = 0
    16'b01110100_11011001 : OUT <= 0;  //116 / 217 = 0
    16'b01110100_11011010 : OUT <= 0;  //116 / 218 = 0
    16'b01110100_11011011 : OUT <= 0;  //116 / 219 = 0
    16'b01110100_11011100 : OUT <= 0;  //116 / 220 = 0
    16'b01110100_11011101 : OUT <= 0;  //116 / 221 = 0
    16'b01110100_11011110 : OUT <= 0;  //116 / 222 = 0
    16'b01110100_11011111 : OUT <= 0;  //116 / 223 = 0
    16'b01110100_11100000 : OUT <= 0;  //116 / 224 = 0
    16'b01110100_11100001 : OUT <= 0;  //116 / 225 = 0
    16'b01110100_11100010 : OUT <= 0;  //116 / 226 = 0
    16'b01110100_11100011 : OUT <= 0;  //116 / 227 = 0
    16'b01110100_11100100 : OUT <= 0;  //116 / 228 = 0
    16'b01110100_11100101 : OUT <= 0;  //116 / 229 = 0
    16'b01110100_11100110 : OUT <= 0;  //116 / 230 = 0
    16'b01110100_11100111 : OUT <= 0;  //116 / 231 = 0
    16'b01110100_11101000 : OUT <= 0;  //116 / 232 = 0
    16'b01110100_11101001 : OUT <= 0;  //116 / 233 = 0
    16'b01110100_11101010 : OUT <= 0;  //116 / 234 = 0
    16'b01110100_11101011 : OUT <= 0;  //116 / 235 = 0
    16'b01110100_11101100 : OUT <= 0;  //116 / 236 = 0
    16'b01110100_11101101 : OUT <= 0;  //116 / 237 = 0
    16'b01110100_11101110 : OUT <= 0;  //116 / 238 = 0
    16'b01110100_11101111 : OUT <= 0;  //116 / 239 = 0
    16'b01110100_11110000 : OUT <= 0;  //116 / 240 = 0
    16'b01110100_11110001 : OUT <= 0;  //116 / 241 = 0
    16'b01110100_11110010 : OUT <= 0;  //116 / 242 = 0
    16'b01110100_11110011 : OUT <= 0;  //116 / 243 = 0
    16'b01110100_11110100 : OUT <= 0;  //116 / 244 = 0
    16'b01110100_11110101 : OUT <= 0;  //116 / 245 = 0
    16'b01110100_11110110 : OUT <= 0;  //116 / 246 = 0
    16'b01110100_11110111 : OUT <= 0;  //116 / 247 = 0
    16'b01110100_11111000 : OUT <= 0;  //116 / 248 = 0
    16'b01110100_11111001 : OUT <= 0;  //116 / 249 = 0
    16'b01110100_11111010 : OUT <= 0;  //116 / 250 = 0
    16'b01110100_11111011 : OUT <= 0;  //116 / 251 = 0
    16'b01110100_11111100 : OUT <= 0;  //116 / 252 = 0
    16'b01110100_11111101 : OUT <= 0;  //116 / 253 = 0
    16'b01110100_11111110 : OUT <= 0;  //116 / 254 = 0
    16'b01110100_11111111 : OUT <= 0;  //116 / 255 = 0
    16'b01110101_00000000 : OUT <= 0;  //117 / 0 = 0
    16'b01110101_00000001 : OUT <= 117;  //117 / 1 = 117
    16'b01110101_00000010 : OUT <= 58;  //117 / 2 = 58
    16'b01110101_00000011 : OUT <= 39;  //117 / 3 = 39
    16'b01110101_00000100 : OUT <= 29;  //117 / 4 = 29
    16'b01110101_00000101 : OUT <= 23;  //117 / 5 = 23
    16'b01110101_00000110 : OUT <= 19;  //117 / 6 = 19
    16'b01110101_00000111 : OUT <= 16;  //117 / 7 = 16
    16'b01110101_00001000 : OUT <= 14;  //117 / 8 = 14
    16'b01110101_00001001 : OUT <= 13;  //117 / 9 = 13
    16'b01110101_00001010 : OUT <= 11;  //117 / 10 = 11
    16'b01110101_00001011 : OUT <= 10;  //117 / 11 = 10
    16'b01110101_00001100 : OUT <= 9;  //117 / 12 = 9
    16'b01110101_00001101 : OUT <= 9;  //117 / 13 = 9
    16'b01110101_00001110 : OUT <= 8;  //117 / 14 = 8
    16'b01110101_00001111 : OUT <= 7;  //117 / 15 = 7
    16'b01110101_00010000 : OUT <= 7;  //117 / 16 = 7
    16'b01110101_00010001 : OUT <= 6;  //117 / 17 = 6
    16'b01110101_00010010 : OUT <= 6;  //117 / 18 = 6
    16'b01110101_00010011 : OUT <= 6;  //117 / 19 = 6
    16'b01110101_00010100 : OUT <= 5;  //117 / 20 = 5
    16'b01110101_00010101 : OUT <= 5;  //117 / 21 = 5
    16'b01110101_00010110 : OUT <= 5;  //117 / 22 = 5
    16'b01110101_00010111 : OUT <= 5;  //117 / 23 = 5
    16'b01110101_00011000 : OUT <= 4;  //117 / 24 = 4
    16'b01110101_00011001 : OUT <= 4;  //117 / 25 = 4
    16'b01110101_00011010 : OUT <= 4;  //117 / 26 = 4
    16'b01110101_00011011 : OUT <= 4;  //117 / 27 = 4
    16'b01110101_00011100 : OUT <= 4;  //117 / 28 = 4
    16'b01110101_00011101 : OUT <= 4;  //117 / 29 = 4
    16'b01110101_00011110 : OUT <= 3;  //117 / 30 = 3
    16'b01110101_00011111 : OUT <= 3;  //117 / 31 = 3
    16'b01110101_00100000 : OUT <= 3;  //117 / 32 = 3
    16'b01110101_00100001 : OUT <= 3;  //117 / 33 = 3
    16'b01110101_00100010 : OUT <= 3;  //117 / 34 = 3
    16'b01110101_00100011 : OUT <= 3;  //117 / 35 = 3
    16'b01110101_00100100 : OUT <= 3;  //117 / 36 = 3
    16'b01110101_00100101 : OUT <= 3;  //117 / 37 = 3
    16'b01110101_00100110 : OUT <= 3;  //117 / 38 = 3
    16'b01110101_00100111 : OUT <= 3;  //117 / 39 = 3
    16'b01110101_00101000 : OUT <= 2;  //117 / 40 = 2
    16'b01110101_00101001 : OUT <= 2;  //117 / 41 = 2
    16'b01110101_00101010 : OUT <= 2;  //117 / 42 = 2
    16'b01110101_00101011 : OUT <= 2;  //117 / 43 = 2
    16'b01110101_00101100 : OUT <= 2;  //117 / 44 = 2
    16'b01110101_00101101 : OUT <= 2;  //117 / 45 = 2
    16'b01110101_00101110 : OUT <= 2;  //117 / 46 = 2
    16'b01110101_00101111 : OUT <= 2;  //117 / 47 = 2
    16'b01110101_00110000 : OUT <= 2;  //117 / 48 = 2
    16'b01110101_00110001 : OUT <= 2;  //117 / 49 = 2
    16'b01110101_00110010 : OUT <= 2;  //117 / 50 = 2
    16'b01110101_00110011 : OUT <= 2;  //117 / 51 = 2
    16'b01110101_00110100 : OUT <= 2;  //117 / 52 = 2
    16'b01110101_00110101 : OUT <= 2;  //117 / 53 = 2
    16'b01110101_00110110 : OUT <= 2;  //117 / 54 = 2
    16'b01110101_00110111 : OUT <= 2;  //117 / 55 = 2
    16'b01110101_00111000 : OUT <= 2;  //117 / 56 = 2
    16'b01110101_00111001 : OUT <= 2;  //117 / 57 = 2
    16'b01110101_00111010 : OUT <= 2;  //117 / 58 = 2
    16'b01110101_00111011 : OUT <= 1;  //117 / 59 = 1
    16'b01110101_00111100 : OUT <= 1;  //117 / 60 = 1
    16'b01110101_00111101 : OUT <= 1;  //117 / 61 = 1
    16'b01110101_00111110 : OUT <= 1;  //117 / 62 = 1
    16'b01110101_00111111 : OUT <= 1;  //117 / 63 = 1
    16'b01110101_01000000 : OUT <= 1;  //117 / 64 = 1
    16'b01110101_01000001 : OUT <= 1;  //117 / 65 = 1
    16'b01110101_01000010 : OUT <= 1;  //117 / 66 = 1
    16'b01110101_01000011 : OUT <= 1;  //117 / 67 = 1
    16'b01110101_01000100 : OUT <= 1;  //117 / 68 = 1
    16'b01110101_01000101 : OUT <= 1;  //117 / 69 = 1
    16'b01110101_01000110 : OUT <= 1;  //117 / 70 = 1
    16'b01110101_01000111 : OUT <= 1;  //117 / 71 = 1
    16'b01110101_01001000 : OUT <= 1;  //117 / 72 = 1
    16'b01110101_01001001 : OUT <= 1;  //117 / 73 = 1
    16'b01110101_01001010 : OUT <= 1;  //117 / 74 = 1
    16'b01110101_01001011 : OUT <= 1;  //117 / 75 = 1
    16'b01110101_01001100 : OUT <= 1;  //117 / 76 = 1
    16'b01110101_01001101 : OUT <= 1;  //117 / 77 = 1
    16'b01110101_01001110 : OUT <= 1;  //117 / 78 = 1
    16'b01110101_01001111 : OUT <= 1;  //117 / 79 = 1
    16'b01110101_01010000 : OUT <= 1;  //117 / 80 = 1
    16'b01110101_01010001 : OUT <= 1;  //117 / 81 = 1
    16'b01110101_01010010 : OUT <= 1;  //117 / 82 = 1
    16'b01110101_01010011 : OUT <= 1;  //117 / 83 = 1
    16'b01110101_01010100 : OUT <= 1;  //117 / 84 = 1
    16'b01110101_01010101 : OUT <= 1;  //117 / 85 = 1
    16'b01110101_01010110 : OUT <= 1;  //117 / 86 = 1
    16'b01110101_01010111 : OUT <= 1;  //117 / 87 = 1
    16'b01110101_01011000 : OUT <= 1;  //117 / 88 = 1
    16'b01110101_01011001 : OUT <= 1;  //117 / 89 = 1
    16'b01110101_01011010 : OUT <= 1;  //117 / 90 = 1
    16'b01110101_01011011 : OUT <= 1;  //117 / 91 = 1
    16'b01110101_01011100 : OUT <= 1;  //117 / 92 = 1
    16'b01110101_01011101 : OUT <= 1;  //117 / 93 = 1
    16'b01110101_01011110 : OUT <= 1;  //117 / 94 = 1
    16'b01110101_01011111 : OUT <= 1;  //117 / 95 = 1
    16'b01110101_01100000 : OUT <= 1;  //117 / 96 = 1
    16'b01110101_01100001 : OUT <= 1;  //117 / 97 = 1
    16'b01110101_01100010 : OUT <= 1;  //117 / 98 = 1
    16'b01110101_01100011 : OUT <= 1;  //117 / 99 = 1
    16'b01110101_01100100 : OUT <= 1;  //117 / 100 = 1
    16'b01110101_01100101 : OUT <= 1;  //117 / 101 = 1
    16'b01110101_01100110 : OUT <= 1;  //117 / 102 = 1
    16'b01110101_01100111 : OUT <= 1;  //117 / 103 = 1
    16'b01110101_01101000 : OUT <= 1;  //117 / 104 = 1
    16'b01110101_01101001 : OUT <= 1;  //117 / 105 = 1
    16'b01110101_01101010 : OUT <= 1;  //117 / 106 = 1
    16'b01110101_01101011 : OUT <= 1;  //117 / 107 = 1
    16'b01110101_01101100 : OUT <= 1;  //117 / 108 = 1
    16'b01110101_01101101 : OUT <= 1;  //117 / 109 = 1
    16'b01110101_01101110 : OUT <= 1;  //117 / 110 = 1
    16'b01110101_01101111 : OUT <= 1;  //117 / 111 = 1
    16'b01110101_01110000 : OUT <= 1;  //117 / 112 = 1
    16'b01110101_01110001 : OUT <= 1;  //117 / 113 = 1
    16'b01110101_01110010 : OUT <= 1;  //117 / 114 = 1
    16'b01110101_01110011 : OUT <= 1;  //117 / 115 = 1
    16'b01110101_01110100 : OUT <= 1;  //117 / 116 = 1
    16'b01110101_01110101 : OUT <= 1;  //117 / 117 = 1
    16'b01110101_01110110 : OUT <= 0;  //117 / 118 = 0
    16'b01110101_01110111 : OUT <= 0;  //117 / 119 = 0
    16'b01110101_01111000 : OUT <= 0;  //117 / 120 = 0
    16'b01110101_01111001 : OUT <= 0;  //117 / 121 = 0
    16'b01110101_01111010 : OUT <= 0;  //117 / 122 = 0
    16'b01110101_01111011 : OUT <= 0;  //117 / 123 = 0
    16'b01110101_01111100 : OUT <= 0;  //117 / 124 = 0
    16'b01110101_01111101 : OUT <= 0;  //117 / 125 = 0
    16'b01110101_01111110 : OUT <= 0;  //117 / 126 = 0
    16'b01110101_01111111 : OUT <= 0;  //117 / 127 = 0
    16'b01110101_10000000 : OUT <= 0;  //117 / 128 = 0
    16'b01110101_10000001 : OUT <= 0;  //117 / 129 = 0
    16'b01110101_10000010 : OUT <= 0;  //117 / 130 = 0
    16'b01110101_10000011 : OUT <= 0;  //117 / 131 = 0
    16'b01110101_10000100 : OUT <= 0;  //117 / 132 = 0
    16'b01110101_10000101 : OUT <= 0;  //117 / 133 = 0
    16'b01110101_10000110 : OUT <= 0;  //117 / 134 = 0
    16'b01110101_10000111 : OUT <= 0;  //117 / 135 = 0
    16'b01110101_10001000 : OUT <= 0;  //117 / 136 = 0
    16'b01110101_10001001 : OUT <= 0;  //117 / 137 = 0
    16'b01110101_10001010 : OUT <= 0;  //117 / 138 = 0
    16'b01110101_10001011 : OUT <= 0;  //117 / 139 = 0
    16'b01110101_10001100 : OUT <= 0;  //117 / 140 = 0
    16'b01110101_10001101 : OUT <= 0;  //117 / 141 = 0
    16'b01110101_10001110 : OUT <= 0;  //117 / 142 = 0
    16'b01110101_10001111 : OUT <= 0;  //117 / 143 = 0
    16'b01110101_10010000 : OUT <= 0;  //117 / 144 = 0
    16'b01110101_10010001 : OUT <= 0;  //117 / 145 = 0
    16'b01110101_10010010 : OUT <= 0;  //117 / 146 = 0
    16'b01110101_10010011 : OUT <= 0;  //117 / 147 = 0
    16'b01110101_10010100 : OUT <= 0;  //117 / 148 = 0
    16'b01110101_10010101 : OUT <= 0;  //117 / 149 = 0
    16'b01110101_10010110 : OUT <= 0;  //117 / 150 = 0
    16'b01110101_10010111 : OUT <= 0;  //117 / 151 = 0
    16'b01110101_10011000 : OUT <= 0;  //117 / 152 = 0
    16'b01110101_10011001 : OUT <= 0;  //117 / 153 = 0
    16'b01110101_10011010 : OUT <= 0;  //117 / 154 = 0
    16'b01110101_10011011 : OUT <= 0;  //117 / 155 = 0
    16'b01110101_10011100 : OUT <= 0;  //117 / 156 = 0
    16'b01110101_10011101 : OUT <= 0;  //117 / 157 = 0
    16'b01110101_10011110 : OUT <= 0;  //117 / 158 = 0
    16'b01110101_10011111 : OUT <= 0;  //117 / 159 = 0
    16'b01110101_10100000 : OUT <= 0;  //117 / 160 = 0
    16'b01110101_10100001 : OUT <= 0;  //117 / 161 = 0
    16'b01110101_10100010 : OUT <= 0;  //117 / 162 = 0
    16'b01110101_10100011 : OUT <= 0;  //117 / 163 = 0
    16'b01110101_10100100 : OUT <= 0;  //117 / 164 = 0
    16'b01110101_10100101 : OUT <= 0;  //117 / 165 = 0
    16'b01110101_10100110 : OUT <= 0;  //117 / 166 = 0
    16'b01110101_10100111 : OUT <= 0;  //117 / 167 = 0
    16'b01110101_10101000 : OUT <= 0;  //117 / 168 = 0
    16'b01110101_10101001 : OUT <= 0;  //117 / 169 = 0
    16'b01110101_10101010 : OUT <= 0;  //117 / 170 = 0
    16'b01110101_10101011 : OUT <= 0;  //117 / 171 = 0
    16'b01110101_10101100 : OUT <= 0;  //117 / 172 = 0
    16'b01110101_10101101 : OUT <= 0;  //117 / 173 = 0
    16'b01110101_10101110 : OUT <= 0;  //117 / 174 = 0
    16'b01110101_10101111 : OUT <= 0;  //117 / 175 = 0
    16'b01110101_10110000 : OUT <= 0;  //117 / 176 = 0
    16'b01110101_10110001 : OUT <= 0;  //117 / 177 = 0
    16'b01110101_10110010 : OUT <= 0;  //117 / 178 = 0
    16'b01110101_10110011 : OUT <= 0;  //117 / 179 = 0
    16'b01110101_10110100 : OUT <= 0;  //117 / 180 = 0
    16'b01110101_10110101 : OUT <= 0;  //117 / 181 = 0
    16'b01110101_10110110 : OUT <= 0;  //117 / 182 = 0
    16'b01110101_10110111 : OUT <= 0;  //117 / 183 = 0
    16'b01110101_10111000 : OUT <= 0;  //117 / 184 = 0
    16'b01110101_10111001 : OUT <= 0;  //117 / 185 = 0
    16'b01110101_10111010 : OUT <= 0;  //117 / 186 = 0
    16'b01110101_10111011 : OUT <= 0;  //117 / 187 = 0
    16'b01110101_10111100 : OUT <= 0;  //117 / 188 = 0
    16'b01110101_10111101 : OUT <= 0;  //117 / 189 = 0
    16'b01110101_10111110 : OUT <= 0;  //117 / 190 = 0
    16'b01110101_10111111 : OUT <= 0;  //117 / 191 = 0
    16'b01110101_11000000 : OUT <= 0;  //117 / 192 = 0
    16'b01110101_11000001 : OUT <= 0;  //117 / 193 = 0
    16'b01110101_11000010 : OUT <= 0;  //117 / 194 = 0
    16'b01110101_11000011 : OUT <= 0;  //117 / 195 = 0
    16'b01110101_11000100 : OUT <= 0;  //117 / 196 = 0
    16'b01110101_11000101 : OUT <= 0;  //117 / 197 = 0
    16'b01110101_11000110 : OUT <= 0;  //117 / 198 = 0
    16'b01110101_11000111 : OUT <= 0;  //117 / 199 = 0
    16'b01110101_11001000 : OUT <= 0;  //117 / 200 = 0
    16'b01110101_11001001 : OUT <= 0;  //117 / 201 = 0
    16'b01110101_11001010 : OUT <= 0;  //117 / 202 = 0
    16'b01110101_11001011 : OUT <= 0;  //117 / 203 = 0
    16'b01110101_11001100 : OUT <= 0;  //117 / 204 = 0
    16'b01110101_11001101 : OUT <= 0;  //117 / 205 = 0
    16'b01110101_11001110 : OUT <= 0;  //117 / 206 = 0
    16'b01110101_11001111 : OUT <= 0;  //117 / 207 = 0
    16'b01110101_11010000 : OUT <= 0;  //117 / 208 = 0
    16'b01110101_11010001 : OUT <= 0;  //117 / 209 = 0
    16'b01110101_11010010 : OUT <= 0;  //117 / 210 = 0
    16'b01110101_11010011 : OUT <= 0;  //117 / 211 = 0
    16'b01110101_11010100 : OUT <= 0;  //117 / 212 = 0
    16'b01110101_11010101 : OUT <= 0;  //117 / 213 = 0
    16'b01110101_11010110 : OUT <= 0;  //117 / 214 = 0
    16'b01110101_11010111 : OUT <= 0;  //117 / 215 = 0
    16'b01110101_11011000 : OUT <= 0;  //117 / 216 = 0
    16'b01110101_11011001 : OUT <= 0;  //117 / 217 = 0
    16'b01110101_11011010 : OUT <= 0;  //117 / 218 = 0
    16'b01110101_11011011 : OUT <= 0;  //117 / 219 = 0
    16'b01110101_11011100 : OUT <= 0;  //117 / 220 = 0
    16'b01110101_11011101 : OUT <= 0;  //117 / 221 = 0
    16'b01110101_11011110 : OUT <= 0;  //117 / 222 = 0
    16'b01110101_11011111 : OUT <= 0;  //117 / 223 = 0
    16'b01110101_11100000 : OUT <= 0;  //117 / 224 = 0
    16'b01110101_11100001 : OUT <= 0;  //117 / 225 = 0
    16'b01110101_11100010 : OUT <= 0;  //117 / 226 = 0
    16'b01110101_11100011 : OUT <= 0;  //117 / 227 = 0
    16'b01110101_11100100 : OUT <= 0;  //117 / 228 = 0
    16'b01110101_11100101 : OUT <= 0;  //117 / 229 = 0
    16'b01110101_11100110 : OUT <= 0;  //117 / 230 = 0
    16'b01110101_11100111 : OUT <= 0;  //117 / 231 = 0
    16'b01110101_11101000 : OUT <= 0;  //117 / 232 = 0
    16'b01110101_11101001 : OUT <= 0;  //117 / 233 = 0
    16'b01110101_11101010 : OUT <= 0;  //117 / 234 = 0
    16'b01110101_11101011 : OUT <= 0;  //117 / 235 = 0
    16'b01110101_11101100 : OUT <= 0;  //117 / 236 = 0
    16'b01110101_11101101 : OUT <= 0;  //117 / 237 = 0
    16'b01110101_11101110 : OUT <= 0;  //117 / 238 = 0
    16'b01110101_11101111 : OUT <= 0;  //117 / 239 = 0
    16'b01110101_11110000 : OUT <= 0;  //117 / 240 = 0
    16'b01110101_11110001 : OUT <= 0;  //117 / 241 = 0
    16'b01110101_11110010 : OUT <= 0;  //117 / 242 = 0
    16'b01110101_11110011 : OUT <= 0;  //117 / 243 = 0
    16'b01110101_11110100 : OUT <= 0;  //117 / 244 = 0
    16'b01110101_11110101 : OUT <= 0;  //117 / 245 = 0
    16'b01110101_11110110 : OUT <= 0;  //117 / 246 = 0
    16'b01110101_11110111 : OUT <= 0;  //117 / 247 = 0
    16'b01110101_11111000 : OUT <= 0;  //117 / 248 = 0
    16'b01110101_11111001 : OUT <= 0;  //117 / 249 = 0
    16'b01110101_11111010 : OUT <= 0;  //117 / 250 = 0
    16'b01110101_11111011 : OUT <= 0;  //117 / 251 = 0
    16'b01110101_11111100 : OUT <= 0;  //117 / 252 = 0
    16'b01110101_11111101 : OUT <= 0;  //117 / 253 = 0
    16'b01110101_11111110 : OUT <= 0;  //117 / 254 = 0
    16'b01110101_11111111 : OUT <= 0;  //117 / 255 = 0
    16'b01110110_00000000 : OUT <= 0;  //118 / 0 = 0
    16'b01110110_00000001 : OUT <= 118;  //118 / 1 = 118
    16'b01110110_00000010 : OUT <= 59;  //118 / 2 = 59
    16'b01110110_00000011 : OUT <= 39;  //118 / 3 = 39
    16'b01110110_00000100 : OUT <= 29;  //118 / 4 = 29
    16'b01110110_00000101 : OUT <= 23;  //118 / 5 = 23
    16'b01110110_00000110 : OUT <= 19;  //118 / 6 = 19
    16'b01110110_00000111 : OUT <= 16;  //118 / 7 = 16
    16'b01110110_00001000 : OUT <= 14;  //118 / 8 = 14
    16'b01110110_00001001 : OUT <= 13;  //118 / 9 = 13
    16'b01110110_00001010 : OUT <= 11;  //118 / 10 = 11
    16'b01110110_00001011 : OUT <= 10;  //118 / 11 = 10
    16'b01110110_00001100 : OUT <= 9;  //118 / 12 = 9
    16'b01110110_00001101 : OUT <= 9;  //118 / 13 = 9
    16'b01110110_00001110 : OUT <= 8;  //118 / 14 = 8
    16'b01110110_00001111 : OUT <= 7;  //118 / 15 = 7
    16'b01110110_00010000 : OUT <= 7;  //118 / 16 = 7
    16'b01110110_00010001 : OUT <= 6;  //118 / 17 = 6
    16'b01110110_00010010 : OUT <= 6;  //118 / 18 = 6
    16'b01110110_00010011 : OUT <= 6;  //118 / 19 = 6
    16'b01110110_00010100 : OUT <= 5;  //118 / 20 = 5
    16'b01110110_00010101 : OUT <= 5;  //118 / 21 = 5
    16'b01110110_00010110 : OUT <= 5;  //118 / 22 = 5
    16'b01110110_00010111 : OUT <= 5;  //118 / 23 = 5
    16'b01110110_00011000 : OUT <= 4;  //118 / 24 = 4
    16'b01110110_00011001 : OUT <= 4;  //118 / 25 = 4
    16'b01110110_00011010 : OUT <= 4;  //118 / 26 = 4
    16'b01110110_00011011 : OUT <= 4;  //118 / 27 = 4
    16'b01110110_00011100 : OUT <= 4;  //118 / 28 = 4
    16'b01110110_00011101 : OUT <= 4;  //118 / 29 = 4
    16'b01110110_00011110 : OUT <= 3;  //118 / 30 = 3
    16'b01110110_00011111 : OUT <= 3;  //118 / 31 = 3
    16'b01110110_00100000 : OUT <= 3;  //118 / 32 = 3
    16'b01110110_00100001 : OUT <= 3;  //118 / 33 = 3
    16'b01110110_00100010 : OUT <= 3;  //118 / 34 = 3
    16'b01110110_00100011 : OUT <= 3;  //118 / 35 = 3
    16'b01110110_00100100 : OUT <= 3;  //118 / 36 = 3
    16'b01110110_00100101 : OUT <= 3;  //118 / 37 = 3
    16'b01110110_00100110 : OUT <= 3;  //118 / 38 = 3
    16'b01110110_00100111 : OUT <= 3;  //118 / 39 = 3
    16'b01110110_00101000 : OUT <= 2;  //118 / 40 = 2
    16'b01110110_00101001 : OUT <= 2;  //118 / 41 = 2
    16'b01110110_00101010 : OUT <= 2;  //118 / 42 = 2
    16'b01110110_00101011 : OUT <= 2;  //118 / 43 = 2
    16'b01110110_00101100 : OUT <= 2;  //118 / 44 = 2
    16'b01110110_00101101 : OUT <= 2;  //118 / 45 = 2
    16'b01110110_00101110 : OUT <= 2;  //118 / 46 = 2
    16'b01110110_00101111 : OUT <= 2;  //118 / 47 = 2
    16'b01110110_00110000 : OUT <= 2;  //118 / 48 = 2
    16'b01110110_00110001 : OUT <= 2;  //118 / 49 = 2
    16'b01110110_00110010 : OUT <= 2;  //118 / 50 = 2
    16'b01110110_00110011 : OUT <= 2;  //118 / 51 = 2
    16'b01110110_00110100 : OUT <= 2;  //118 / 52 = 2
    16'b01110110_00110101 : OUT <= 2;  //118 / 53 = 2
    16'b01110110_00110110 : OUT <= 2;  //118 / 54 = 2
    16'b01110110_00110111 : OUT <= 2;  //118 / 55 = 2
    16'b01110110_00111000 : OUT <= 2;  //118 / 56 = 2
    16'b01110110_00111001 : OUT <= 2;  //118 / 57 = 2
    16'b01110110_00111010 : OUT <= 2;  //118 / 58 = 2
    16'b01110110_00111011 : OUT <= 2;  //118 / 59 = 2
    16'b01110110_00111100 : OUT <= 1;  //118 / 60 = 1
    16'b01110110_00111101 : OUT <= 1;  //118 / 61 = 1
    16'b01110110_00111110 : OUT <= 1;  //118 / 62 = 1
    16'b01110110_00111111 : OUT <= 1;  //118 / 63 = 1
    16'b01110110_01000000 : OUT <= 1;  //118 / 64 = 1
    16'b01110110_01000001 : OUT <= 1;  //118 / 65 = 1
    16'b01110110_01000010 : OUT <= 1;  //118 / 66 = 1
    16'b01110110_01000011 : OUT <= 1;  //118 / 67 = 1
    16'b01110110_01000100 : OUT <= 1;  //118 / 68 = 1
    16'b01110110_01000101 : OUT <= 1;  //118 / 69 = 1
    16'b01110110_01000110 : OUT <= 1;  //118 / 70 = 1
    16'b01110110_01000111 : OUT <= 1;  //118 / 71 = 1
    16'b01110110_01001000 : OUT <= 1;  //118 / 72 = 1
    16'b01110110_01001001 : OUT <= 1;  //118 / 73 = 1
    16'b01110110_01001010 : OUT <= 1;  //118 / 74 = 1
    16'b01110110_01001011 : OUT <= 1;  //118 / 75 = 1
    16'b01110110_01001100 : OUT <= 1;  //118 / 76 = 1
    16'b01110110_01001101 : OUT <= 1;  //118 / 77 = 1
    16'b01110110_01001110 : OUT <= 1;  //118 / 78 = 1
    16'b01110110_01001111 : OUT <= 1;  //118 / 79 = 1
    16'b01110110_01010000 : OUT <= 1;  //118 / 80 = 1
    16'b01110110_01010001 : OUT <= 1;  //118 / 81 = 1
    16'b01110110_01010010 : OUT <= 1;  //118 / 82 = 1
    16'b01110110_01010011 : OUT <= 1;  //118 / 83 = 1
    16'b01110110_01010100 : OUT <= 1;  //118 / 84 = 1
    16'b01110110_01010101 : OUT <= 1;  //118 / 85 = 1
    16'b01110110_01010110 : OUT <= 1;  //118 / 86 = 1
    16'b01110110_01010111 : OUT <= 1;  //118 / 87 = 1
    16'b01110110_01011000 : OUT <= 1;  //118 / 88 = 1
    16'b01110110_01011001 : OUT <= 1;  //118 / 89 = 1
    16'b01110110_01011010 : OUT <= 1;  //118 / 90 = 1
    16'b01110110_01011011 : OUT <= 1;  //118 / 91 = 1
    16'b01110110_01011100 : OUT <= 1;  //118 / 92 = 1
    16'b01110110_01011101 : OUT <= 1;  //118 / 93 = 1
    16'b01110110_01011110 : OUT <= 1;  //118 / 94 = 1
    16'b01110110_01011111 : OUT <= 1;  //118 / 95 = 1
    16'b01110110_01100000 : OUT <= 1;  //118 / 96 = 1
    16'b01110110_01100001 : OUT <= 1;  //118 / 97 = 1
    16'b01110110_01100010 : OUT <= 1;  //118 / 98 = 1
    16'b01110110_01100011 : OUT <= 1;  //118 / 99 = 1
    16'b01110110_01100100 : OUT <= 1;  //118 / 100 = 1
    16'b01110110_01100101 : OUT <= 1;  //118 / 101 = 1
    16'b01110110_01100110 : OUT <= 1;  //118 / 102 = 1
    16'b01110110_01100111 : OUT <= 1;  //118 / 103 = 1
    16'b01110110_01101000 : OUT <= 1;  //118 / 104 = 1
    16'b01110110_01101001 : OUT <= 1;  //118 / 105 = 1
    16'b01110110_01101010 : OUT <= 1;  //118 / 106 = 1
    16'b01110110_01101011 : OUT <= 1;  //118 / 107 = 1
    16'b01110110_01101100 : OUT <= 1;  //118 / 108 = 1
    16'b01110110_01101101 : OUT <= 1;  //118 / 109 = 1
    16'b01110110_01101110 : OUT <= 1;  //118 / 110 = 1
    16'b01110110_01101111 : OUT <= 1;  //118 / 111 = 1
    16'b01110110_01110000 : OUT <= 1;  //118 / 112 = 1
    16'b01110110_01110001 : OUT <= 1;  //118 / 113 = 1
    16'b01110110_01110010 : OUT <= 1;  //118 / 114 = 1
    16'b01110110_01110011 : OUT <= 1;  //118 / 115 = 1
    16'b01110110_01110100 : OUT <= 1;  //118 / 116 = 1
    16'b01110110_01110101 : OUT <= 1;  //118 / 117 = 1
    16'b01110110_01110110 : OUT <= 1;  //118 / 118 = 1
    16'b01110110_01110111 : OUT <= 0;  //118 / 119 = 0
    16'b01110110_01111000 : OUT <= 0;  //118 / 120 = 0
    16'b01110110_01111001 : OUT <= 0;  //118 / 121 = 0
    16'b01110110_01111010 : OUT <= 0;  //118 / 122 = 0
    16'b01110110_01111011 : OUT <= 0;  //118 / 123 = 0
    16'b01110110_01111100 : OUT <= 0;  //118 / 124 = 0
    16'b01110110_01111101 : OUT <= 0;  //118 / 125 = 0
    16'b01110110_01111110 : OUT <= 0;  //118 / 126 = 0
    16'b01110110_01111111 : OUT <= 0;  //118 / 127 = 0
    16'b01110110_10000000 : OUT <= 0;  //118 / 128 = 0
    16'b01110110_10000001 : OUT <= 0;  //118 / 129 = 0
    16'b01110110_10000010 : OUT <= 0;  //118 / 130 = 0
    16'b01110110_10000011 : OUT <= 0;  //118 / 131 = 0
    16'b01110110_10000100 : OUT <= 0;  //118 / 132 = 0
    16'b01110110_10000101 : OUT <= 0;  //118 / 133 = 0
    16'b01110110_10000110 : OUT <= 0;  //118 / 134 = 0
    16'b01110110_10000111 : OUT <= 0;  //118 / 135 = 0
    16'b01110110_10001000 : OUT <= 0;  //118 / 136 = 0
    16'b01110110_10001001 : OUT <= 0;  //118 / 137 = 0
    16'b01110110_10001010 : OUT <= 0;  //118 / 138 = 0
    16'b01110110_10001011 : OUT <= 0;  //118 / 139 = 0
    16'b01110110_10001100 : OUT <= 0;  //118 / 140 = 0
    16'b01110110_10001101 : OUT <= 0;  //118 / 141 = 0
    16'b01110110_10001110 : OUT <= 0;  //118 / 142 = 0
    16'b01110110_10001111 : OUT <= 0;  //118 / 143 = 0
    16'b01110110_10010000 : OUT <= 0;  //118 / 144 = 0
    16'b01110110_10010001 : OUT <= 0;  //118 / 145 = 0
    16'b01110110_10010010 : OUT <= 0;  //118 / 146 = 0
    16'b01110110_10010011 : OUT <= 0;  //118 / 147 = 0
    16'b01110110_10010100 : OUT <= 0;  //118 / 148 = 0
    16'b01110110_10010101 : OUT <= 0;  //118 / 149 = 0
    16'b01110110_10010110 : OUT <= 0;  //118 / 150 = 0
    16'b01110110_10010111 : OUT <= 0;  //118 / 151 = 0
    16'b01110110_10011000 : OUT <= 0;  //118 / 152 = 0
    16'b01110110_10011001 : OUT <= 0;  //118 / 153 = 0
    16'b01110110_10011010 : OUT <= 0;  //118 / 154 = 0
    16'b01110110_10011011 : OUT <= 0;  //118 / 155 = 0
    16'b01110110_10011100 : OUT <= 0;  //118 / 156 = 0
    16'b01110110_10011101 : OUT <= 0;  //118 / 157 = 0
    16'b01110110_10011110 : OUT <= 0;  //118 / 158 = 0
    16'b01110110_10011111 : OUT <= 0;  //118 / 159 = 0
    16'b01110110_10100000 : OUT <= 0;  //118 / 160 = 0
    16'b01110110_10100001 : OUT <= 0;  //118 / 161 = 0
    16'b01110110_10100010 : OUT <= 0;  //118 / 162 = 0
    16'b01110110_10100011 : OUT <= 0;  //118 / 163 = 0
    16'b01110110_10100100 : OUT <= 0;  //118 / 164 = 0
    16'b01110110_10100101 : OUT <= 0;  //118 / 165 = 0
    16'b01110110_10100110 : OUT <= 0;  //118 / 166 = 0
    16'b01110110_10100111 : OUT <= 0;  //118 / 167 = 0
    16'b01110110_10101000 : OUT <= 0;  //118 / 168 = 0
    16'b01110110_10101001 : OUT <= 0;  //118 / 169 = 0
    16'b01110110_10101010 : OUT <= 0;  //118 / 170 = 0
    16'b01110110_10101011 : OUT <= 0;  //118 / 171 = 0
    16'b01110110_10101100 : OUT <= 0;  //118 / 172 = 0
    16'b01110110_10101101 : OUT <= 0;  //118 / 173 = 0
    16'b01110110_10101110 : OUT <= 0;  //118 / 174 = 0
    16'b01110110_10101111 : OUT <= 0;  //118 / 175 = 0
    16'b01110110_10110000 : OUT <= 0;  //118 / 176 = 0
    16'b01110110_10110001 : OUT <= 0;  //118 / 177 = 0
    16'b01110110_10110010 : OUT <= 0;  //118 / 178 = 0
    16'b01110110_10110011 : OUT <= 0;  //118 / 179 = 0
    16'b01110110_10110100 : OUT <= 0;  //118 / 180 = 0
    16'b01110110_10110101 : OUT <= 0;  //118 / 181 = 0
    16'b01110110_10110110 : OUT <= 0;  //118 / 182 = 0
    16'b01110110_10110111 : OUT <= 0;  //118 / 183 = 0
    16'b01110110_10111000 : OUT <= 0;  //118 / 184 = 0
    16'b01110110_10111001 : OUT <= 0;  //118 / 185 = 0
    16'b01110110_10111010 : OUT <= 0;  //118 / 186 = 0
    16'b01110110_10111011 : OUT <= 0;  //118 / 187 = 0
    16'b01110110_10111100 : OUT <= 0;  //118 / 188 = 0
    16'b01110110_10111101 : OUT <= 0;  //118 / 189 = 0
    16'b01110110_10111110 : OUT <= 0;  //118 / 190 = 0
    16'b01110110_10111111 : OUT <= 0;  //118 / 191 = 0
    16'b01110110_11000000 : OUT <= 0;  //118 / 192 = 0
    16'b01110110_11000001 : OUT <= 0;  //118 / 193 = 0
    16'b01110110_11000010 : OUT <= 0;  //118 / 194 = 0
    16'b01110110_11000011 : OUT <= 0;  //118 / 195 = 0
    16'b01110110_11000100 : OUT <= 0;  //118 / 196 = 0
    16'b01110110_11000101 : OUT <= 0;  //118 / 197 = 0
    16'b01110110_11000110 : OUT <= 0;  //118 / 198 = 0
    16'b01110110_11000111 : OUT <= 0;  //118 / 199 = 0
    16'b01110110_11001000 : OUT <= 0;  //118 / 200 = 0
    16'b01110110_11001001 : OUT <= 0;  //118 / 201 = 0
    16'b01110110_11001010 : OUT <= 0;  //118 / 202 = 0
    16'b01110110_11001011 : OUT <= 0;  //118 / 203 = 0
    16'b01110110_11001100 : OUT <= 0;  //118 / 204 = 0
    16'b01110110_11001101 : OUT <= 0;  //118 / 205 = 0
    16'b01110110_11001110 : OUT <= 0;  //118 / 206 = 0
    16'b01110110_11001111 : OUT <= 0;  //118 / 207 = 0
    16'b01110110_11010000 : OUT <= 0;  //118 / 208 = 0
    16'b01110110_11010001 : OUT <= 0;  //118 / 209 = 0
    16'b01110110_11010010 : OUT <= 0;  //118 / 210 = 0
    16'b01110110_11010011 : OUT <= 0;  //118 / 211 = 0
    16'b01110110_11010100 : OUT <= 0;  //118 / 212 = 0
    16'b01110110_11010101 : OUT <= 0;  //118 / 213 = 0
    16'b01110110_11010110 : OUT <= 0;  //118 / 214 = 0
    16'b01110110_11010111 : OUT <= 0;  //118 / 215 = 0
    16'b01110110_11011000 : OUT <= 0;  //118 / 216 = 0
    16'b01110110_11011001 : OUT <= 0;  //118 / 217 = 0
    16'b01110110_11011010 : OUT <= 0;  //118 / 218 = 0
    16'b01110110_11011011 : OUT <= 0;  //118 / 219 = 0
    16'b01110110_11011100 : OUT <= 0;  //118 / 220 = 0
    16'b01110110_11011101 : OUT <= 0;  //118 / 221 = 0
    16'b01110110_11011110 : OUT <= 0;  //118 / 222 = 0
    16'b01110110_11011111 : OUT <= 0;  //118 / 223 = 0
    16'b01110110_11100000 : OUT <= 0;  //118 / 224 = 0
    16'b01110110_11100001 : OUT <= 0;  //118 / 225 = 0
    16'b01110110_11100010 : OUT <= 0;  //118 / 226 = 0
    16'b01110110_11100011 : OUT <= 0;  //118 / 227 = 0
    16'b01110110_11100100 : OUT <= 0;  //118 / 228 = 0
    16'b01110110_11100101 : OUT <= 0;  //118 / 229 = 0
    16'b01110110_11100110 : OUT <= 0;  //118 / 230 = 0
    16'b01110110_11100111 : OUT <= 0;  //118 / 231 = 0
    16'b01110110_11101000 : OUT <= 0;  //118 / 232 = 0
    16'b01110110_11101001 : OUT <= 0;  //118 / 233 = 0
    16'b01110110_11101010 : OUT <= 0;  //118 / 234 = 0
    16'b01110110_11101011 : OUT <= 0;  //118 / 235 = 0
    16'b01110110_11101100 : OUT <= 0;  //118 / 236 = 0
    16'b01110110_11101101 : OUT <= 0;  //118 / 237 = 0
    16'b01110110_11101110 : OUT <= 0;  //118 / 238 = 0
    16'b01110110_11101111 : OUT <= 0;  //118 / 239 = 0
    16'b01110110_11110000 : OUT <= 0;  //118 / 240 = 0
    16'b01110110_11110001 : OUT <= 0;  //118 / 241 = 0
    16'b01110110_11110010 : OUT <= 0;  //118 / 242 = 0
    16'b01110110_11110011 : OUT <= 0;  //118 / 243 = 0
    16'b01110110_11110100 : OUT <= 0;  //118 / 244 = 0
    16'b01110110_11110101 : OUT <= 0;  //118 / 245 = 0
    16'b01110110_11110110 : OUT <= 0;  //118 / 246 = 0
    16'b01110110_11110111 : OUT <= 0;  //118 / 247 = 0
    16'b01110110_11111000 : OUT <= 0;  //118 / 248 = 0
    16'b01110110_11111001 : OUT <= 0;  //118 / 249 = 0
    16'b01110110_11111010 : OUT <= 0;  //118 / 250 = 0
    16'b01110110_11111011 : OUT <= 0;  //118 / 251 = 0
    16'b01110110_11111100 : OUT <= 0;  //118 / 252 = 0
    16'b01110110_11111101 : OUT <= 0;  //118 / 253 = 0
    16'b01110110_11111110 : OUT <= 0;  //118 / 254 = 0
    16'b01110110_11111111 : OUT <= 0;  //118 / 255 = 0
    16'b01110111_00000000 : OUT <= 0;  //119 / 0 = 0
    16'b01110111_00000001 : OUT <= 119;  //119 / 1 = 119
    16'b01110111_00000010 : OUT <= 59;  //119 / 2 = 59
    16'b01110111_00000011 : OUT <= 39;  //119 / 3 = 39
    16'b01110111_00000100 : OUT <= 29;  //119 / 4 = 29
    16'b01110111_00000101 : OUT <= 23;  //119 / 5 = 23
    16'b01110111_00000110 : OUT <= 19;  //119 / 6 = 19
    16'b01110111_00000111 : OUT <= 17;  //119 / 7 = 17
    16'b01110111_00001000 : OUT <= 14;  //119 / 8 = 14
    16'b01110111_00001001 : OUT <= 13;  //119 / 9 = 13
    16'b01110111_00001010 : OUT <= 11;  //119 / 10 = 11
    16'b01110111_00001011 : OUT <= 10;  //119 / 11 = 10
    16'b01110111_00001100 : OUT <= 9;  //119 / 12 = 9
    16'b01110111_00001101 : OUT <= 9;  //119 / 13 = 9
    16'b01110111_00001110 : OUT <= 8;  //119 / 14 = 8
    16'b01110111_00001111 : OUT <= 7;  //119 / 15 = 7
    16'b01110111_00010000 : OUT <= 7;  //119 / 16 = 7
    16'b01110111_00010001 : OUT <= 7;  //119 / 17 = 7
    16'b01110111_00010010 : OUT <= 6;  //119 / 18 = 6
    16'b01110111_00010011 : OUT <= 6;  //119 / 19 = 6
    16'b01110111_00010100 : OUT <= 5;  //119 / 20 = 5
    16'b01110111_00010101 : OUT <= 5;  //119 / 21 = 5
    16'b01110111_00010110 : OUT <= 5;  //119 / 22 = 5
    16'b01110111_00010111 : OUT <= 5;  //119 / 23 = 5
    16'b01110111_00011000 : OUT <= 4;  //119 / 24 = 4
    16'b01110111_00011001 : OUT <= 4;  //119 / 25 = 4
    16'b01110111_00011010 : OUT <= 4;  //119 / 26 = 4
    16'b01110111_00011011 : OUT <= 4;  //119 / 27 = 4
    16'b01110111_00011100 : OUT <= 4;  //119 / 28 = 4
    16'b01110111_00011101 : OUT <= 4;  //119 / 29 = 4
    16'b01110111_00011110 : OUT <= 3;  //119 / 30 = 3
    16'b01110111_00011111 : OUT <= 3;  //119 / 31 = 3
    16'b01110111_00100000 : OUT <= 3;  //119 / 32 = 3
    16'b01110111_00100001 : OUT <= 3;  //119 / 33 = 3
    16'b01110111_00100010 : OUT <= 3;  //119 / 34 = 3
    16'b01110111_00100011 : OUT <= 3;  //119 / 35 = 3
    16'b01110111_00100100 : OUT <= 3;  //119 / 36 = 3
    16'b01110111_00100101 : OUT <= 3;  //119 / 37 = 3
    16'b01110111_00100110 : OUT <= 3;  //119 / 38 = 3
    16'b01110111_00100111 : OUT <= 3;  //119 / 39 = 3
    16'b01110111_00101000 : OUT <= 2;  //119 / 40 = 2
    16'b01110111_00101001 : OUT <= 2;  //119 / 41 = 2
    16'b01110111_00101010 : OUT <= 2;  //119 / 42 = 2
    16'b01110111_00101011 : OUT <= 2;  //119 / 43 = 2
    16'b01110111_00101100 : OUT <= 2;  //119 / 44 = 2
    16'b01110111_00101101 : OUT <= 2;  //119 / 45 = 2
    16'b01110111_00101110 : OUT <= 2;  //119 / 46 = 2
    16'b01110111_00101111 : OUT <= 2;  //119 / 47 = 2
    16'b01110111_00110000 : OUT <= 2;  //119 / 48 = 2
    16'b01110111_00110001 : OUT <= 2;  //119 / 49 = 2
    16'b01110111_00110010 : OUT <= 2;  //119 / 50 = 2
    16'b01110111_00110011 : OUT <= 2;  //119 / 51 = 2
    16'b01110111_00110100 : OUT <= 2;  //119 / 52 = 2
    16'b01110111_00110101 : OUT <= 2;  //119 / 53 = 2
    16'b01110111_00110110 : OUT <= 2;  //119 / 54 = 2
    16'b01110111_00110111 : OUT <= 2;  //119 / 55 = 2
    16'b01110111_00111000 : OUT <= 2;  //119 / 56 = 2
    16'b01110111_00111001 : OUT <= 2;  //119 / 57 = 2
    16'b01110111_00111010 : OUT <= 2;  //119 / 58 = 2
    16'b01110111_00111011 : OUT <= 2;  //119 / 59 = 2
    16'b01110111_00111100 : OUT <= 1;  //119 / 60 = 1
    16'b01110111_00111101 : OUT <= 1;  //119 / 61 = 1
    16'b01110111_00111110 : OUT <= 1;  //119 / 62 = 1
    16'b01110111_00111111 : OUT <= 1;  //119 / 63 = 1
    16'b01110111_01000000 : OUT <= 1;  //119 / 64 = 1
    16'b01110111_01000001 : OUT <= 1;  //119 / 65 = 1
    16'b01110111_01000010 : OUT <= 1;  //119 / 66 = 1
    16'b01110111_01000011 : OUT <= 1;  //119 / 67 = 1
    16'b01110111_01000100 : OUT <= 1;  //119 / 68 = 1
    16'b01110111_01000101 : OUT <= 1;  //119 / 69 = 1
    16'b01110111_01000110 : OUT <= 1;  //119 / 70 = 1
    16'b01110111_01000111 : OUT <= 1;  //119 / 71 = 1
    16'b01110111_01001000 : OUT <= 1;  //119 / 72 = 1
    16'b01110111_01001001 : OUT <= 1;  //119 / 73 = 1
    16'b01110111_01001010 : OUT <= 1;  //119 / 74 = 1
    16'b01110111_01001011 : OUT <= 1;  //119 / 75 = 1
    16'b01110111_01001100 : OUT <= 1;  //119 / 76 = 1
    16'b01110111_01001101 : OUT <= 1;  //119 / 77 = 1
    16'b01110111_01001110 : OUT <= 1;  //119 / 78 = 1
    16'b01110111_01001111 : OUT <= 1;  //119 / 79 = 1
    16'b01110111_01010000 : OUT <= 1;  //119 / 80 = 1
    16'b01110111_01010001 : OUT <= 1;  //119 / 81 = 1
    16'b01110111_01010010 : OUT <= 1;  //119 / 82 = 1
    16'b01110111_01010011 : OUT <= 1;  //119 / 83 = 1
    16'b01110111_01010100 : OUT <= 1;  //119 / 84 = 1
    16'b01110111_01010101 : OUT <= 1;  //119 / 85 = 1
    16'b01110111_01010110 : OUT <= 1;  //119 / 86 = 1
    16'b01110111_01010111 : OUT <= 1;  //119 / 87 = 1
    16'b01110111_01011000 : OUT <= 1;  //119 / 88 = 1
    16'b01110111_01011001 : OUT <= 1;  //119 / 89 = 1
    16'b01110111_01011010 : OUT <= 1;  //119 / 90 = 1
    16'b01110111_01011011 : OUT <= 1;  //119 / 91 = 1
    16'b01110111_01011100 : OUT <= 1;  //119 / 92 = 1
    16'b01110111_01011101 : OUT <= 1;  //119 / 93 = 1
    16'b01110111_01011110 : OUT <= 1;  //119 / 94 = 1
    16'b01110111_01011111 : OUT <= 1;  //119 / 95 = 1
    16'b01110111_01100000 : OUT <= 1;  //119 / 96 = 1
    16'b01110111_01100001 : OUT <= 1;  //119 / 97 = 1
    16'b01110111_01100010 : OUT <= 1;  //119 / 98 = 1
    16'b01110111_01100011 : OUT <= 1;  //119 / 99 = 1
    16'b01110111_01100100 : OUT <= 1;  //119 / 100 = 1
    16'b01110111_01100101 : OUT <= 1;  //119 / 101 = 1
    16'b01110111_01100110 : OUT <= 1;  //119 / 102 = 1
    16'b01110111_01100111 : OUT <= 1;  //119 / 103 = 1
    16'b01110111_01101000 : OUT <= 1;  //119 / 104 = 1
    16'b01110111_01101001 : OUT <= 1;  //119 / 105 = 1
    16'b01110111_01101010 : OUT <= 1;  //119 / 106 = 1
    16'b01110111_01101011 : OUT <= 1;  //119 / 107 = 1
    16'b01110111_01101100 : OUT <= 1;  //119 / 108 = 1
    16'b01110111_01101101 : OUT <= 1;  //119 / 109 = 1
    16'b01110111_01101110 : OUT <= 1;  //119 / 110 = 1
    16'b01110111_01101111 : OUT <= 1;  //119 / 111 = 1
    16'b01110111_01110000 : OUT <= 1;  //119 / 112 = 1
    16'b01110111_01110001 : OUT <= 1;  //119 / 113 = 1
    16'b01110111_01110010 : OUT <= 1;  //119 / 114 = 1
    16'b01110111_01110011 : OUT <= 1;  //119 / 115 = 1
    16'b01110111_01110100 : OUT <= 1;  //119 / 116 = 1
    16'b01110111_01110101 : OUT <= 1;  //119 / 117 = 1
    16'b01110111_01110110 : OUT <= 1;  //119 / 118 = 1
    16'b01110111_01110111 : OUT <= 1;  //119 / 119 = 1
    16'b01110111_01111000 : OUT <= 0;  //119 / 120 = 0
    16'b01110111_01111001 : OUT <= 0;  //119 / 121 = 0
    16'b01110111_01111010 : OUT <= 0;  //119 / 122 = 0
    16'b01110111_01111011 : OUT <= 0;  //119 / 123 = 0
    16'b01110111_01111100 : OUT <= 0;  //119 / 124 = 0
    16'b01110111_01111101 : OUT <= 0;  //119 / 125 = 0
    16'b01110111_01111110 : OUT <= 0;  //119 / 126 = 0
    16'b01110111_01111111 : OUT <= 0;  //119 / 127 = 0
    16'b01110111_10000000 : OUT <= 0;  //119 / 128 = 0
    16'b01110111_10000001 : OUT <= 0;  //119 / 129 = 0
    16'b01110111_10000010 : OUT <= 0;  //119 / 130 = 0
    16'b01110111_10000011 : OUT <= 0;  //119 / 131 = 0
    16'b01110111_10000100 : OUT <= 0;  //119 / 132 = 0
    16'b01110111_10000101 : OUT <= 0;  //119 / 133 = 0
    16'b01110111_10000110 : OUT <= 0;  //119 / 134 = 0
    16'b01110111_10000111 : OUT <= 0;  //119 / 135 = 0
    16'b01110111_10001000 : OUT <= 0;  //119 / 136 = 0
    16'b01110111_10001001 : OUT <= 0;  //119 / 137 = 0
    16'b01110111_10001010 : OUT <= 0;  //119 / 138 = 0
    16'b01110111_10001011 : OUT <= 0;  //119 / 139 = 0
    16'b01110111_10001100 : OUT <= 0;  //119 / 140 = 0
    16'b01110111_10001101 : OUT <= 0;  //119 / 141 = 0
    16'b01110111_10001110 : OUT <= 0;  //119 / 142 = 0
    16'b01110111_10001111 : OUT <= 0;  //119 / 143 = 0
    16'b01110111_10010000 : OUT <= 0;  //119 / 144 = 0
    16'b01110111_10010001 : OUT <= 0;  //119 / 145 = 0
    16'b01110111_10010010 : OUT <= 0;  //119 / 146 = 0
    16'b01110111_10010011 : OUT <= 0;  //119 / 147 = 0
    16'b01110111_10010100 : OUT <= 0;  //119 / 148 = 0
    16'b01110111_10010101 : OUT <= 0;  //119 / 149 = 0
    16'b01110111_10010110 : OUT <= 0;  //119 / 150 = 0
    16'b01110111_10010111 : OUT <= 0;  //119 / 151 = 0
    16'b01110111_10011000 : OUT <= 0;  //119 / 152 = 0
    16'b01110111_10011001 : OUT <= 0;  //119 / 153 = 0
    16'b01110111_10011010 : OUT <= 0;  //119 / 154 = 0
    16'b01110111_10011011 : OUT <= 0;  //119 / 155 = 0
    16'b01110111_10011100 : OUT <= 0;  //119 / 156 = 0
    16'b01110111_10011101 : OUT <= 0;  //119 / 157 = 0
    16'b01110111_10011110 : OUT <= 0;  //119 / 158 = 0
    16'b01110111_10011111 : OUT <= 0;  //119 / 159 = 0
    16'b01110111_10100000 : OUT <= 0;  //119 / 160 = 0
    16'b01110111_10100001 : OUT <= 0;  //119 / 161 = 0
    16'b01110111_10100010 : OUT <= 0;  //119 / 162 = 0
    16'b01110111_10100011 : OUT <= 0;  //119 / 163 = 0
    16'b01110111_10100100 : OUT <= 0;  //119 / 164 = 0
    16'b01110111_10100101 : OUT <= 0;  //119 / 165 = 0
    16'b01110111_10100110 : OUT <= 0;  //119 / 166 = 0
    16'b01110111_10100111 : OUT <= 0;  //119 / 167 = 0
    16'b01110111_10101000 : OUT <= 0;  //119 / 168 = 0
    16'b01110111_10101001 : OUT <= 0;  //119 / 169 = 0
    16'b01110111_10101010 : OUT <= 0;  //119 / 170 = 0
    16'b01110111_10101011 : OUT <= 0;  //119 / 171 = 0
    16'b01110111_10101100 : OUT <= 0;  //119 / 172 = 0
    16'b01110111_10101101 : OUT <= 0;  //119 / 173 = 0
    16'b01110111_10101110 : OUT <= 0;  //119 / 174 = 0
    16'b01110111_10101111 : OUT <= 0;  //119 / 175 = 0
    16'b01110111_10110000 : OUT <= 0;  //119 / 176 = 0
    16'b01110111_10110001 : OUT <= 0;  //119 / 177 = 0
    16'b01110111_10110010 : OUT <= 0;  //119 / 178 = 0
    16'b01110111_10110011 : OUT <= 0;  //119 / 179 = 0
    16'b01110111_10110100 : OUT <= 0;  //119 / 180 = 0
    16'b01110111_10110101 : OUT <= 0;  //119 / 181 = 0
    16'b01110111_10110110 : OUT <= 0;  //119 / 182 = 0
    16'b01110111_10110111 : OUT <= 0;  //119 / 183 = 0
    16'b01110111_10111000 : OUT <= 0;  //119 / 184 = 0
    16'b01110111_10111001 : OUT <= 0;  //119 / 185 = 0
    16'b01110111_10111010 : OUT <= 0;  //119 / 186 = 0
    16'b01110111_10111011 : OUT <= 0;  //119 / 187 = 0
    16'b01110111_10111100 : OUT <= 0;  //119 / 188 = 0
    16'b01110111_10111101 : OUT <= 0;  //119 / 189 = 0
    16'b01110111_10111110 : OUT <= 0;  //119 / 190 = 0
    16'b01110111_10111111 : OUT <= 0;  //119 / 191 = 0
    16'b01110111_11000000 : OUT <= 0;  //119 / 192 = 0
    16'b01110111_11000001 : OUT <= 0;  //119 / 193 = 0
    16'b01110111_11000010 : OUT <= 0;  //119 / 194 = 0
    16'b01110111_11000011 : OUT <= 0;  //119 / 195 = 0
    16'b01110111_11000100 : OUT <= 0;  //119 / 196 = 0
    16'b01110111_11000101 : OUT <= 0;  //119 / 197 = 0
    16'b01110111_11000110 : OUT <= 0;  //119 / 198 = 0
    16'b01110111_11000111 : OUT <= 0;  //119 / 199 = 0
    16'b01110111_11001000 : OUT <= 0;  //119 / 200 = 0
    16'b01110111_11001001 : OUT <= 0;  //119 / 201 = 0
    16'b01110111_11001010 : OUT <= 0;  //119 / 202 = 0
    16'b01110111_11001011 : OUT <= 0;  //119 / 203 = 0
    16'b01110111_11001100 : OUT <= 0;  //119 / 204 = 0
    16'b01110111_11001101 : OUT <= 0;  //119 / 205 = 0
    16'b01110111_11001110 : OUT <= 0;  //119 / 206 = 0
    16'b01110111_11001111 : OUT <= 0;  //119 / 207 = 0
    16'b01110111_11010000 : OUT <= 0;  //119 / 208 = 0
    16'b01110111_11010001 : OUT <= 0;  //119 / 209 = 0
    16'b01110111_11010010 : OUT <= 0;  //119 / 210 = 0
    16'b01110111_11010011 : OUT <= 0;  //119 / 211 = 0
    16'b01110111_11010100 : OUT <= 0;  //119 / 212 = 0
    16'b01110111_11010101 : OUT <= 0;  //119 / 213 = 0
    16'b01110111_11010110 : OUT <= 0;  //119 / 214 = 0
    16'b01110111_11010111 : OUT <= 0;  //119 / 215 = 0
    16'b01110111_11011000 : OUT <= 0;  //119 / 216 = 0
    16'b01110111_11011001 : OUT <= 0;  //119 / 217 = 0
    16'b01110111_11011010 : OUT <= 0;  //119 / 218 = 0
    16'b01110111_11011011 : OUT <= 0;  //119 / 219 = 0
    16'b01110111_11011100 : OUT <= 0;  //119 / 220 = 0
    16'b01110111_11011101 : OUT <= 0;  //119 / 221 = 0
    16'b01110111_11011110 : OUT <= 0;  //119 / 222 = 0
    16'b01110111_11011111 : OUT <= 0;  //119 / 223 = 0
    16'b01110111_11100000 : OUT <= 0;  //119 / 224 = 0
    16'b01110111_11100001 : OUT <= 0;  //119 / 225 = 0
    16'b01110111_11100010 : OUT <= 0;  //119 / 226 = 0
    16'b01110111_11100011 : OUT <= 0;  //119 / 227 = 0
    16'b01110111_11100100 : OUT <= 0;  //119 / 228 = 0
    16'b01110111_11100101 : OUT <= 0;  //119 / 229 = 0
    16'b01110111_11100110 : OUT <= 0;  //119 / 230 = 0
    16'b01110111_11100111 : OUT <= 0;  //119 / 231 = 0
    16'b01110111_11101000 : OUT <= 0;  //119 / 232 = 0
    16'b01110111_11101001 : OUT <= 0;  //119 / 233 = 0
    16'b01110111_11101010 : OUT <= 0;  //119 / 234 = 0
    16'b01110111_11101011 : OUT <= 0;  //119 / 235 = 0
    16'b01110111_11101100 : OUT <= 0;  //119 / 236 = 0
    16'b01110111_11101101 : OUT <= 0;  //119 / 237 = 0
    16'b01110111_11101110 : OUT <= 0;  //119 / 238 = 0
    16'b01110111_11101111 : OUT <= 0;  //119 / 239 = 0
    16'b01110111_11110000 : OUT <= 0;  //119 / 240 = 0
    16'b01110111_11110001 : OUT <= 0;  //119 / 241 = 0
    16'b01110111_11110010 : OUT <= 0;  //119 / 242 = 0
    16'b01110111_11110011 : OUT <= 0;  //119 / 243 = 0
    16'b01110111_11110100 : OUT <= 0;  //119 / 244 = 0
    16'b01110111_11110101 : OUT <= 0;  //119 / 245 = 0
    16'b01110111_11110110 : OUT <= 0;  //119 / 246 = 0
    16'b01110111_11110111 : OUT <= 0;  //119 / 247 = 0
    16'b01110111_11111000 : OUT <= 0;  //119 / 248 = 0
    16'b01110111_11111001 : OUT <= 0;  //119 / 249 = 0
    16'b01110111_11111010 : OUT <= 0;  //119 / 250 = 0
    16'b01110111_11111011 : OUT <= 0;  //119 / 251 = 0
    16'b01110111_11111100 : OUT <= 0;  //119 / 252 = 0
    16'b01110111_11111101 : OUT <= 0;  //119 / 253 = 0
    16'b01110111_11111110 : OUT <= 0;  //119 / 254 = 0
    16'b01110111_11111111 : OUT <= 0;  //119 / 255 = 0
    16'b01111000_00000000 : OUT <= 0;  //120 / 0 = 0
    16'b01111000_00000001 : OUT <= 120;  //120 / 1 = 120
    16'b01111000_00000010 : OUT <= 60;  //120 / 2 = 60
    16'b01111000_00000011 : OUT <= 40;  //120 / 3 = 40
    16'b01111000_00000100 : OUT <= 30;  //120 / 4 = 30
    16'b01111000_00000101 : OUT <= 24;  //120 / 5 = 24
    16'b01111000_00000110 : OUT <= 20;  //120 / 6 = 20
    16'b01111000_00000111 : OUT <= 17;  //120 / 7 = 17
    16'b01111000_00001000 : OUT <= 15;  //120 / 8 = 15
    16'b01111000_00001001 : OUT <= 13;  //120 / 9 = 13
    16'b01111000_00001010 : OUT <= 12;  //120 / 10 = 12
    16'b01111000_00001011 : OUT <= 10;  //120 / 11 = 10
    16'b01111000_00001100 : OUT <= 10;  //120 / 12 = 10
    16'b01111000_00001101 : OUT <= 9;  //120 / 13 = 9
    16'b01111000_00001110 : OUT <= 8;  //120 / 14 = 8
    16'b01111000_00001111 : OUT <= 8;  //120 / 15 = 8
    16'b01111000_00010000 : OUT <= 7;  //120 / 16 = 7
    16'b01111000_00010001 : OUT <= 7;  //120 / 17 = 7
    16'b01111000_00010010 : OUT <= 6;  //120 / 18 = 6
    16'b01111000_00010011 : OUT <= 6;  //120 / 19 = 6
    16'b01111000_00010100 : OUT <= 6;  //120 / 20 = 6
    16'b01111000_00010101 : OUT <= 5;  //120 / 21 = 5
    16'b01111000_00010110 : OUT <= 5;  //120 / 22 = 5
    16'b01111000_00010111 : OUT <= 5;  //120 / 23 = 5
    16'b01111000_00011000 : OUT <= 5;  //120 / 24 = 5
    16'b01111000_00011001 : OUT <= 4;  //120 / 25 = 4
    16'b01111000_00011010 : OUT <= 4;  //120 / 26 = 4
    16'b01111000_00011011 : OUT <= 4;  //120 / 27 = 4
    16'b01111000_00011100 : OUT <= 4;  //120 / 28 = 4
    16'b01111000_00011101 : OUT <= 4;  //120 / 29 = 4
    16'b01111000_00011110 : OUT <= 4;  //120 / 30 = 4
    16'b01111000_00011111 : OUT <= 3;  //120 / 31 = 3
    16'b01111000_00100000 : OUT <= 3;  //120 / 32 = 3
    16'b01111000_00100001 : OUT <= 3;  //120 / 33 = 3
    16'b01111000_00100010 : OUT <= 3;  //120 / 34 = 3
    16'b01111000_00100011 : OUT <= 3;  //120 / 35 = 3
    16'b01111000_00100100 : OUT <= 3;  //120 / 36 = 3
    16'b01111000_00100101 : OUT <= 3;  //120 / 37 = 3
    16'b01111000_00100110 : OUT <= 3;  //120 / 38 = 3
    16'b01111000_00100111 : OUT <= 3;  //120 / 39 = 3
    16'b01111000_00101000 : OUT <= 3;  //120 / 40 = 3
    16'b01111000_00101001 : OUT <= 2;  //120 / 41 = 2
    16'b01111000_00101010 : OUT <= 2;  //120 / 42 = 2
    16'b01111000_00101011 : OUT <= 2;  //120 / 43 = 2
    16'b01111000_00101100 : OUT <= 2;  //120 / 44 = 2
    16'b01111000_00101101 : OUT <= 2;  //120 / 45 = 2
    16'b01111000_00101110 : OUT <= 2;  //120 / 46 = 2
    16'b01111000_00101111 : OUT <= 2;  //120 / 47 = 2
    16'b01111000_00110000 : OUT <= 2;  //120 / 48 = 2
    16'b01111000_00110001 : OUT <= 2;  //120 / 49 = 2
    16'b01111000_00110010 : OUT <= 2;  //120 / 50 = 2
    16'b01111000_00110011 : OUT <= 2;  //120 / 51 = 2
    16'b01111000_00110100 : OUT <= 2;  //120 / 52 = 2
    16'b01111000_00110101 : OUT <= 2;  //120 / 53 = 2
    16'b01111000_00110110 : OUT <= 2;  //120 / 54 = 2
    16'b01111000_00110111 : OUT <= 2;  //120 / 55 = 2
    16'b01111000_00111000 : OUT <= 2;  //120 / 56 = 2
    16'b01111000_00111001 : OUT <= 2;  //120 / 57 = 2
    16'b01111000_00111010 : OUT <= 2;  //120 / 58 = 2
    16'b01111000_00111011 : OUT <= 2;  //120 / 59 = 2
    16'b01111000_00111100 : OUT <= 2;  //120 / 60 = 2
    16'b01111000_00111101 : OUT <= 1;  //120 / 61 = 1
    16'b01111000_00111110 : OUT <= 1;  //120 / 62 = 1
    16'b01111000_00111111 : OUT <= 1;  //120 / 63 = 1
    16'b01111000_01000000 : OUT <= 1;  //120 / 64 = 1
    16'b01111000_01000001 : OUT <= 1;  //120 / 65 = 1
    16'b01111000_01000010 : OUT <= 1;  //120 / 66 = 1
    16'b01111000_01000011 : OUT <= 1;  //120 / 67 = 1
    16'b01111000_01000100 : OUT <= 1;  //120 / 68 = 1
    16'b01111000_01000101 : OUT <= 1;  //120 / 69 = 1
    16'b01111000_01000110 : OUT <= 1;  //120 / 70 = 1
    16'b01111000_01000111 : OUT <= 1;  //120 / 71 = 1
    16'b01111000_01001000 : OUT <= 1;  //120 / 72 = 1
    16'b01111000_01001001 : OUT <= 1;  //120 / 73 = 1
    16'b01111000_01001010 : OUT <= 1;  //120 / 74 = 1
    16'b01111000_01001011 : OUT <= 1;  //120 / 75 = 1
    16'b01111000_01001100 : OUT <= 1;  //120 / 76 = 1
    16'b01111000_01001101 : OUT <= 1;  //120 / 77 = 1
    16'b01111000_01001110 : OUT <= 1;  //120 / 78 = 1
    16'b01111000_01001111 : OUT <= 1;  //120 / 79 = 1
    16'b01111000_01010000 : OUT <= 1;  //120 / 80 = 1
    16'b01111000_01010001 : OUT <= 1;  //120 / 81 = 1
    16'b01111000_01010010 : OUT <= 1;  //120 / 82 = 1
    16'b01111000_01010011 : OUT <= 1;  //120 / 83 = 1
    16'b01111000_01010100 : OUT <= 1;  //120 / 84 = 1
    16'b01111000_01010101 : OUT <= 1;  //120 / 85 = 1
    16'b01111000_01010110 : OUT <= 1;  //120 / 86 = 1
    16'b01111000_01010111 : OUT <= 1;  //120 / 87 = 1
    16'b01111000_01011000 : OUT <= 1;  //120 / 88 = 1
    16'b01111000_01011001 : OUT <= 1;  //120 / 89 = 1
    16'b01111000_01011010 : OUT <= 1;  //120 / 90 = 1
    16'b01111000_01011011 : OUT <= 1;  //120 / 91 = 1
    16'b01111000_01011100 : OUT <= 1;  //120 / 92 = 1
    16'b01111000_01011101 : OUT <= 1;  //120 / 93 = 1
    16'b01111000_01011110 : OUT <= 1;  //120 / 94 = 1
    16'b01111000_01011111 : OUT <= 1;  //120 / 95 = 1
    16'b01111000_01100000 : OUT <= 1;  //120 / 96 = 1
    16'b01111000_01100001 : OUT <= 1;  //120 / 97 = 1
    16'b01111000_01100010 : OUT <= 1;  //120 / 98 = 1
    16'b01111000_01100011 : OUT <= 1;  //120 / 99 = 1
    16'b01111000_01100100 : OUT <= 1;  //120 / 100 = 1
    16'b01111000_01100101 : OUT <= 1;  //120 / 101 = 1
    16'b01111000_01100110 : OUT <= 1;  //120 / 102 = 1
    16'b01111000_01100111 : OUT <= 1;  //120 / 103 = 1
    16'b01111000_01101000 : OUT <= 1;  //120 / 104 = 1
    16'b01111000_01101001 : OUT <= 1;  //120 / 105 = 1
    16'b01111000_01101010 : OUT <= 1;  //120 / 106 = 1
    16'b01111000_01101011 : OUT <= 1;  //120 / 107 = 1
    16'b01111000_01101100 : OUT <= 1;  //120 / 108 = 1
    16'b01111000_01101101 : OUT <= 1;  //120 / 109 = 1
    16'b01111000_01101110 : OUT <= 1;  //120 / 110 = 1
    16'b01111000_01101111 : OUT <= 1;  //120 / 111 = 1
    16'b01111000_01110000 : OUT <= 1;  //120 / 112 = 1
    16'b01111000_01110001 : OUT <= 1;  //120 / 113 = 1
    16'b01111000_01110010 : OUT <= 1;  //120 / 114 = 1
    16'b01111000_01110011 : OUT <= 1;  //120 / 115 = 1
    16'b01111000_01110100 : OUT <= 1;  //120 / 116 = 1
    16'b01111000_01110101 : OUT <= 1;  //120 / 117 = 1
    16'b01111000_01110110 : OUT <= 1;  //120 / 118 = 1
    16'b01111000_01110111 : OUT <= 1;  //120 / 119 = 1
    16'b01111000_01111000 : OUT <= 1;  //120 / 120 = 1
    16'b01111000_01111001 : OUT <= 0;  //120 / 121 = 0
    16'b01111000_01111010 : OUT <= 0;  //120 / 122 = 0
    16'b01111000_01111011 : OUT <= 0;  //120 / 123 = 0
    16'b01111000_01111100 : OUT <= 0;  //120 / 124 = 0
    16'b01111000_01111101 : OUT <= 0;  //120 / 125 = 0
    16'b01111000_01111110 : OUT <= 0;  //120 / 126 = 0
    16'b01111000_01111111 : OUT <= 0;  //120 / 127 = 0
    16'b01111000_10000000 : OUT <= 0;  //120 / 128 = 0
    16'b01111000_10000001 : OUT <= 0;  //120 / 129 = 0
    16'b01111000_10000010 : OUT <= 0;  //120 / 130 = 0
    16'b01111000_10000011 : OUT <= 0;  //120 / 131 = 0
    16'b01111000_10000100 : OUT <= 0;  //120 / 132 = 0
    16'b01111000_10000101 : OUT <= 0;  //120 / 133 = 0
    16'b01111000_10000110 : OUT <= 0;  //120 / 134 = 0
    16'b01111000_10000111 : OUT <= 0;  //120 / 135 = 0
    16'b01111000_10001000 : OUT <= 0;  //120 / 136 = 0
    16'b01111000_10001001 : OUT <= 0;  //120 / 137 = 0
    16'b01111000_10001010 : OUT <= 0;  //120 / 138 = 0
    16'b01111000_10001011 : OUT <= 0;  //120 / 139 = 0
    16'b01111000_10001100 : OUT <= 0;  //120 / 140 = 0
    16'b01111000_10001101 : OUT <= 0;  //120 / 141 = 0
    16'b01111000_10001110 : OUT <= 0;  //120 / 142 = 0
    16'b01111000_10001111 : OUT <= 0;  //120 / 143 = 0
    16'b01111000_10010000 : OUT <= 0;  //120 / 144 = 0
    16'b01111000_10010001 : OUT <= 0;  //120 / 145 = 0
    16'b01111000_10010010 : OUT <= 0;  //120 / 146 = 0
    16'b01111000_10010011 : OUT <= 0;  //120 / 147 = 0
    16'b01111000_10010100 : OUT <= 0;  //120 / 148 = 0
    16'b01111000_10010101 : OUT <= 0;  //120 / 149 = 0
    16'b01111000_10010110 : OUT <= 0;  //120 / 150 = 0
    16'b01111000_10010111 : OUT <= 0;  //120 / 151 = 0
    16'b01111000_10011000 : OUT <= 0;  //120 / 152 = 0
    16'b01111000_10011001 : OUT <= 0;  //120 / 153 = 0
    16'b01111000_10011010 : OUT <= 0;  //120 / 154 = 0
    16'b01111000_10011011 : OUT <= 0;  //120 / 155 = 0
    16'b01111000_10011100 : OUT <= 0;  //120 / 156 = 0
    16'b01111000_10011101 : OUT <= 0;  //120 / 157 = 0
    16'b01111000_10011110 : OUT <= 0;  //120 / 158 = 0
    16'b01111000_10011111 : OUT <= 0;  //120 / 159 = 0
    16'b01111000_10100000 : OUT <= 0;  //120 / 160 = 0
    16'b01111000_10100001 : OUT <= 0;  //120 / 161 = 0
    16'b01111000_10100010 : OUT <= 0;  //120 / 162 = 0
    16'b01111000_10100011 : OUT <= 0;  //120 / 163 = 0
    16'b01111000_10100100 : OUT <= 0;  //120 / 164 = 0
    16'b01111000_10100101 : OUT <= 0;  //120 / 165 = 0
    16'b01111000_10100110 : OUT <= 0;  //120 / 166 = 0
    16'b01111000_10100111 : OUT <= 0;  //120 / 167 = 0
    16'b01111000_10101000 : OUT <= 0;  //120 / 168 = 0
    16'b01111000_10101001 : OUT <= 0;  //120 / 169 = 0
    16'b01111000_10101010 : OUT <= 0;  //120 / 170 = 0
    16'b01111000_10101011 : OUT <= 0;  //120 / 171 = 0
    16'b01111000_10101100 : OUT <= 0;  //120 / 172 = 0
    16'b01111000_10101101 : OUT <= 0;  //120 / 173 = 0
    16'b01111000_10101110 : OUT <= 0;  //120 / 174 = 0
    16'b01111000_10101111 : OUT <= 0;  //120 / 175 = 0
    16'b01111000_10110000 : OUT <= 0;  //120 / 176 = 0
    16'b01111000_10110001 : OUT <= 0;  //120 / 177 = 0
    16'b01111000_10110010 : OUT <= 0;  //120 / 178 = 0
    16'b01111000_10110011 : OUT <= 0;  //120 / 179 = 0
    16'b01111000_10110100 : OUT <= 0;  //120 / 180 = 0
    16'b01111000_10110101 : OUT <= 0;  //120 / 181 = 0
    16'b01111000_10110110 : OUT <= 0;  //120 / 182 = 0
    16'b01111000_10110111 : OUT <= 0;  //120 / 183 = 0
    16'b01111000_10111000 : OUT <= 0;  //120 / 184 = 0
    16'b01111000_10111001 : OUT <= 0;  //120 / 185 = 0
    16'b01111000_10111010 : OUT <= 0;  //120 / 186 = 0
    16'b01111000_10111011 : OUT <= 0;  //120 / 187 = 0
    16'b01111000_10111100 : OUT <= 0;  //120 / 188 = 0
    16'b01111000_10111101 : OUT <= 0;  //120 / 189 = 0
    16'b01111000_10111110 : OUT <= 0;  //120 / 190 = 0
    16'b01111000_10111111 : OUT <= 0;  //120 / 191 = 0
    16'b01111000_11000000 : OUT <= 0;  //120 / 192 = 0
    16'b01111000_11000001 : OUT <= 0;  //120 / 193 = 0
    16'b01111000_11000010 : OUT <= 0;  //120 / 194 = 0
    16'b01111000_11000011 : OUT <= 0;  //120 / 195 = 0
    16'b01111000_11000100 : OUT <= 0;  //120 / 196 = 0
    16'b01111000_11000101 : OUT <= 0;  //120 / 197 = 0
    16'b01111000_11000110 : OUT <= 0;  //120 / 198 = 0
    16'b01111000_11000111 : OUT <= 0;  //120 / 199 = 0
    16'b01111000_11001000 : OUT <= 0;  //120 / 200 = 0
    16'b01111000_11001001 : OUT <= 0;  //120 / 201 = 0
    16'b01111000_11001010 : OUT <= 0;  //120 / 202 = 0
    16'b01111000_11001011 : OUT <= 0;  //120 / 203 = 0
    16'b01111000_11001100 : OUT <= 0;  //120 / 204 = 0
    16'b01111000_11001101 : OUT <= 0;  //120 / 205 = 0
    16'b01111000_11001110 : OUT <= 0;  //120 / 206 = 0
    16'b01111000_11001111 : OUT <= 0;  //120 / 207 = 0
    16'b01111000_11010000 : OUT <= 0;  //120 / 208 = 0
    16'b01111000_11010001 : OUT <= 0;  //120 / 209 = 0
    16'b01111000_11010010 : OUT <= 0;  //120 / 210 = 0
    16'b01111000_11010011 : OUT <= 0;  //120 / 211 = 0
    16'b01111000_11010100 : OUT <= 0;  //120 / 212 = 0
    16'b01111000_11010101 : OUT <= 0;  //120 / 213 = 0
    16'b01111000_11010110 : OUT <= 0;  //120 / 214 = 0
    16'b01111000_11010111 : OUT <= 0;  //120 / 215 = 0
    16'b01111000_11011000 : OUT <= 0;  //120 / 216 = 0
    16'b01111000_11011001 : OUT <= 0;  //120 / 217 = 0
    16'b01111000_11011010 : OUT <= 0;  //120 / 218 = 0
    16'b01111000_11011011 : OUT <= 0;  //120 / 219 = 0
    16'b01111000_11011100 : OUT <= 0;  //120 / 220 = 0
    16'b01111000_11011101 : OUT <= 0;  //120 / 221 = 0
    16'b01111000_11011110 : OUT <= 0;  //120 / 222 = 0
    16'b01111000_11011111 : OUT <= 0;  //120 / 223 = 0
    16'b01111000_11100000 : OUT <= 0;  //120 / 224 = 0
    16'b01111000_11100001 : OUT <= 0;  //120 / 225 = 0
    16'b01111000_11100010 : OUT <= 0;  //120 / 226 = 0
    16'b01111000_11100011 : OUT <= 0;  //120 / 227 = 0
    16'b01111000_11100100 : OUT <= 0;  //120 / 228 = 0
    16'b01111000_11100101 : OUT <= 0;  //120 / 229 = 0
    16'b01111000_11100110 : OUT <= 0;  //120 / 230 = 0
    16'b01111000_11100111 : OUT <= 0;  //120 / 231 = 0
    16'b01111000_11101000 : OUT <= 0;  //120 / 232 = 0
    16'b01111000_11101001 : OUT <= 0;  //120 / 233 = 0
    16'b01111000_11101010 : OUT <= 0;  //120 / 234 = 0
    16'b01111000_11101011 : OUT <= 0;  //120 / 235 = 0
    16'b01111000_11101100 : OUT <= 0;  //120 / 236 = 0
    16'b01111000_11101101 : OUT <= 0;  //120 / 237 = 0
    16'b01111000_11101110 : OUT <= 0;  //120 / 238 = 0
    16'b01111000_11101111 : OUT <= 0;  //120 / 239 = 0
    16'b01111000_11110000 : OUT <= 0;  //120 / 240 = 0
    16'b01111000_11110001 : OUT <= 0;  //120 / 241 = 0
    16'b01111000_11110010 : OUT <= 0;  //120 / 242 = 0
    16'b01111000_11110011 : OUT <= 0;  //120 / 243 = 0
    16'b01111000_11110100 : OUT <= 0;  //120 / 244 = 0
    16'b01111000_11110101 : OUT <= 0;  //120 / 245 = 0
    16'b01111000_11110110 : OUT <= 0;  //120 / 246 = 0
    16'b01111000_11110111 : OUT <= 0;  //120 / 247 = 0
    16'b01111000_11111000 : OUT <= 0;  //120 / 248 = 0
    16'b01111000_11111001 : OUT <= 0;  //120 / 249 = 0
    16'b01111000_11111010 : OUT <= 0;  //120 / 250 = 0
    16'b01111000_11111011 : OUT <= 0;  //120 / 251 = 0
    16'b01111000_11111100 : OUT <= 0;  //120 / 252 = 0
    16'b01111000_11111101 : OUT <= 0;  //120 / 253 = 0
    16'b01111000_11111110 : OUT <= 0;  //120 / 254 = 0
    16'b01111000_11111111 : OUT <= 0;  //120 / 255 = 0
    16'b01111001_00000000 : OUT <= 0;  //121 / 0 = 0
    16'b01111001_00000001 : OUT <= 121;  //121 / 1 = 121
    16'b01111001_00000010 : OUT <= 60;  //121 / 2 = 60
    16'b01111001_00000011 : OUT <= 40;  //121 / 3 = 40
    16'b01111001_00000100 : OUT <= 30;  //121 / 4 = 30
    16'b01111001_00000101 : OUT <= 24;  //121 / 5 = 24
    16'b01111001_00000110 : OUT <= 20;  //121 / 6 = 20
    16'b01111001_00000111 : OUT <= 17;  //121 / 7 = 17
    16'b01111001_00001000 : OUT <= 15;  //121 / 8 = 15
    16'b01111001_00001001 : OUT <= 13;  //121 / 9 = 13
    16'b01111001_00001010 : OUT <= 12;  //121 / 10 = 12
    16'b01111001_00001011 : OUT <= 11;  //121 / 11 = 11
    16'b01111001_00001100 : OUT <= 10;  //121 / 12 = 10
    16'b01111001_00001101 : OUT <= 9;  //121 / 13 = 9
    16'b01111001_00001110 : OUT <= 8;  //121 / 14 = 8
    16'b01111001_00001111 : OUT <= 8;  //121 / 15 = 8
    16'b01111001_00010000 : OUT <= 7;  //121 / 16 = 7
    16'b01111001_00010001 : OUT <= 7;  //121 / 17 = 7
    16'b01111001_00010010 : OUT <= 6;  //121 / 18 = 6
    16'b01111001_00010011 : OUT <= 6;  //121 / 19 = 6
    16'b01111001_00010100 : OUT <= 6;  //121 / 20 = 6
    16'b01111001_00010101 : OUT <= 5;  //121 / 21 = 5
    16'b01111001_00010110 : OUT <= 5;  //121 / 22 = 5
    16'b01111001_00010111 : OUT <= 5;  //121 / 23 = 5
    16'b01111001_00011000 : OUT <= 5;  //121 / 24 = 5
    16'b01111001_00011001 : OUT <= 4;  //121 / 25 = 4
    16'b01111001_00011010 : OUT <= 4;  //121 / 26 = 4
    16'b01111001_00011011 : OUT <= 4;  //121 / 27 = 4
    16'b01111001_00011100 : OUT <= 4;  //121 / 28 = 4
    16'b01111001_00011101 : OUT <= 4;  //121 / 29 = 4
    16'b01111001_00011110 : OUT <= 4;  //121 / 30 = 4
    16'b01111001_00011111 : OUT <= 3;  //121 / 31 = 3
    16'b01111001_00100000 : OUT <= 3;  //121 / 32 = 3
    16'b01111001_00100001 : OUT <= 3;  //121 / 33 = 3
    16'b01111001_00100010 : OUT <= 3;  //121 / 34 = 3
    16'b01111001_00100011 : OUT <= 3;  //121 / 35 = 3
    16'b01111001_00100100 : OUT <= 3;  //121 / 36 = 3
    16'b01111001_00100101 : OUT <= 3;  //121 / 37 = 3
    16'b01111001_00100110 : OUT <= 3;  //121 / 38 = 3
    16'b01111001_00100111 : OUT <= 3;  //121 / 39 = 3
    16'b01111001_00101000 : OUT <= 3;  //121 / 40 = 3
    16'b01111001_00101001 : OUT <= 2;  //121 / 41 = 2
    16'b01111001_00101010 : OUT <= 2;  //121 / 42 = 2
    16'b01111001_00101011 : OUT <= 2;  //121 / 43 = 2
    16'b01111001_00101100 : OUT <= 2;  //121 / 44 = 2
    16'b01111001_00101101 : OUT <= 2;  //121 / 45 = 2
    16'b01111001_00101110 : OUT <= 2;  //121 / 46 = 2
    16'b01111001_00101111 : OUT <= 2;  //121 / 47 = 2
    16'b01111001_00110000 : OUT <= 2;  //121 / 48 = 2
    16'b01111001_00110001 : OUT <= 2;  //121 / 49 = 2
    16'b01111001_00110010 : OUT <= 2;  //121 / 50 = 2
    16'b01111001_00110011 : OUT <= 2;  //121 / 51 = 2
    16'b01111001_00110100 : OUT <= 2;  //121 / 52 = 2
    16'b01111001_00110101 : OUT <= 2;  //121 / 53 = 2
    16'b01111001_00110110 : OUT <= 2;  //121 / 54 = 2
    16'b01111001_00110111 : OUT <= 2;  //121 / 55 = 2
    16'b01111001_00111000 : OUT <= 2;  //121 / 56 = 2
    16'b01111001_00111001 : OUT <= 2;  //121 / 57 = 2
    16'b01111001_00111010 : OUT <= 2;  //121 / 58 = 2
    16'b01111001_00111011 : OUT <= 2;  //121 / 59 = 2
    16'b01111001_00111100 : OUT <= 2;  //121 / 60 = 2
    16'b01111001_00111101 : OUT <= 1;  //121 / 61 = 1
    16'b01111001_00111110 : OUT <= 1;  //121 / 62 = 1
    16'b01111001_00111111 : OUT <= 1;  //121 / 63 = 1
    16'b01111001_01000000 : OUT <= 1;  //121 / 64 = 1
    16'b01111001_01000001 : OUT <= 1;  //121 / 65 = 1
    16'b01111001_01000010 : OUT <= 1;  //121 / 66 = 1
    16'b01111001_01000011 : OUT <= 1;  //121 / 67 = 1
    16'b01111001_01000100 : OUT <= 1;  //121 / 68 = 1
    16'b01111001_01000101 : OUT <= 1;  //121 / 69 = 1
    16'b01111001_01000110 : OUT <= 1;  //121 / 70 = 1
    16'b01111001_01000111 : OUT <= 1;  //121 / 71 = 1
    16'b01111001_01001000 : OUT <= 1;  //121 / 72 = 1
    16'b01111001_01001001 : OUT <= 1;  //121 / 73 = 1
    16'b01111001_01001010 : OUT <= 1;  //121 / 74 = 1
    16'b01111001_01001011 : OUT <= 1;  //121 / 75 = 1
    16'b01111001_01001100 : OUT <= 1;  //121 / 76 = 1
    16'b01111001_01001101 : OUT <= 1;  //121 / 77 = 1
    16'b01111001_01001110 : OUT <= 1;  //121 / 78 = 1
    16'b01111001_01001111 : OUT <= 1;  //121 / 79 = 1
    16'b01111001_01010000 : OUT <= 1;  //121 / 80 = 1
    16'b01111001_01010001 : OUT <= 1;  //121 / 81 = 1
    16'b01111001_01010010 : OUT <= 1;  //121 / 82 = 1
    16'b01111001_01010011 : OUT <= 1;  //121 / 83 = 1
    16'b01111001_01010100 : OUT <= 1;  //121 / 84 = 1
    16'b01111001_01010101 : OUT <= 1;  //121 / 85 = 1
    16'b01111001_01010110 : OUT <= 1;  //121 / 86 = 1
    16'b01111001_01010111 : OUT <= 1;  //121 / 87 = 1
    16'b01111001_01011000 : OUT <= 1;  //121 / 88 = 1
    16'b01111001_01011001 : OUT <= 1;  //121 / 89 = 1
    16'b01111001_01011010 : OUT <= 1;  //121 / 90 = 1
    16'b01111001_01011011 : OUT <= 1;  //121 / 91 = 1
    16'b01111001_01011100 : OUT <= 1;  //121 / 92 = 1
    16'b01111001_01011101 : OUT <= 1;  //121 / 93 = 1
    16'b01111001_01011110 : OUT <= 1;  //121 / 94 = 1
    16'b01111001_01011111 : OUT <= 1;  //121 / 95 = 1
    16'b01111001_01100000 : OUT <= 1;  //121 / 96 = 1
    16'b01111001_01100001 : OUT <= 1;  //121 / 97 = 1
    16'b01111001_01100010 : OUT <= 1;  //121 / 98 = 1
    16'b01111001_01100011 : OUT <= 1;  //121 / 99 = 1
    16'b01111001_01100100 : OUT <= 1;  //121 / 100 = 1
    16'b01111001_01100101 : OUT <= 1;  //121 / 101 = 1
    16'b01111001_01100110 : OUT <= 1;  //121 / 102 = 1
    16'b01111001_01100111 : OUT <= 1;  //121 / 103 = 1
    16'b01111001_01101000 : OUT <= 1;  //121 / 104 = 1
    16'b01111001_01101001 : OUT <= 1;  //121 / 105 = 1
    16'b01111001_01101010 : OUT <= 1;  //121 / 106 = 1
    16'b01111001_01101011 : OUT <= 1;  //121 / 107 = 1
    16'b01111001_01101100 : OUT <= 1;  //121 / 108 = 1
    16'b01111001_01101101 : OUT <= 1;  //121 / 109 = 1
    16'b01111001_01101110 : OUT <= 1;  //121 / 110 = 1
    16'b01111001_01101111 : OUT <= 1;  //121 / 111 = 1
    16'b01111001_01110000 : OUT <= 1;  //121 / 112 = 1
    16'b01111001_01110001 : OUT <= 1;  //121 / 113 = 1
    16'b01111001_01110010 : OUT <= 1;  //121 / 114 = 1
    16'b01111001_01110011 : OUT <= 1;  //121 / 115 = 1
    16'b01111001_01110100 : OUT <= 1;  //121 / 116 = 1
    16'b01111001_01110101 : OUT <= 1;  //121 / 117 = 1
    16'b01111001_01110110 : OUT <= 1;  //121 / 118 = 1
    16'b01111001_01110111 : OUT <= 1;  //121 / 119 = 1
    16'b01111001_01111000 : OUT <= 1;  //121 / 120 = 1
    16'b01111001_01111001 : OUT <= 1;  //121 / 121 = 1
    16'b01111001_01111010 : OUT <= 0;  //121 / 122 = 0
    16'b01111001_01111011 : OUT <= 0;  //121 / 123 = 0
    16'b01111001_01111100 : OUT <= 0;  //121 / 124 = 0
    16'b01111001_01111101 : OUT <= 0;  //121 / 125 = 0
    16'b01111001_01111110 : OUT <= 0;  //121 / 126 = 0
    16'b01111001_01111111 : OUT <= 0;  //121 / 127 = 0
    16'b01111001_10000000 : OUT <= 0;  //121 / 128 = 0
    16'b01111001_10000001 : OUT <= 0;  //121 / 129 = 0
    16'b01111001_10000010 : OUT <= 0;  //121 / 130 = 0
    16'b01111001_10000011 : OUT <= 0;  //121 / 131 = 0
    16'b01111001_10000100 : OUT <= 0;  //121 / 132 = 0
    16'b01111001_10000101 : OUT <= 0;  //121 / 133 = 0
    16'b01111001_10000110 : OUT <= 0;  //121 / 134 = 0
    16'b01111001_10000111 : OUT <= 0;  //121 / 135 = 0
    16'b01111001_10001000 : OUT <= 0;  //121 / 136 = 0
    16'b01111001_10001001 : OUT <= 0;  //121 / 137 = 0
    16'b01111001_10001010 : OUT <= 0;  //121 / 138 = 0
    16'b01111001_10001011 : OUT <= 0;  //121 / 139 = 0
    16'b01111001_10001100 : OUT <= 0;  //121 / 140 = 0
    16'b01111001_10001101 : OUT <= 0;  //121 / 141 = 0
    16'b01111001_10001110 : OUT <= 0;  //121 / 142 = 0
    16'b01111001_10001111 : OUT <= 0;  //121 / 143 = 0
    16'b01111001_10010000 : OUT <= 0;  //121 / 144 = 0
    16'b01111001_10010001 : OUT <= 0;  //121 / 145 = 0
    16'b01111001_10010010 : OUT <= 0;  //121 / 146 = 0
    16'b01111001_10010011 : OUT <= 0;  //121 / 147 = 0
    16'b01111001_10010100 : OUT <= 0;  //121 / 148 = 0
    16'b01111001_10010101 : OUT <= 0;  //121 / 149 = 0
    16'b01111001_10010110 : OUT <= 0;  //121 / 150 = 0
    16'b01111001_10010111 : OUT <= 0;  //121 / 151 = 0
    16'b01111001_10011000 : OUT <= 0;  //121 / 152 = 0
    16'b01111001_10011001 : OUT <= 0;  //121 / 153 = 0
    16'b01111001_10011010 : OUT <= 0;  //121 / 154 = 0
    16'b01111001_10011011 : OUT <= 0;  //121 / 155 = 0
    16'b01111001_10011100 : OUT <= 0;  //121 / 156 = 0
    16'b01111001_10011101 : OUT <= 0;  //121 / 157 = 0
    16'b01111001_10011110 : OUT <= 0;  //121 / 158 = 0
    16'b01111001_10011111 : OUT <= 0;  //121 / 159 = 0
    16'b01111001_10100000 : OUT <= 0;  //121 / 160 = 0
    16'b01111001_10100001 : OUT <= 0;  //121 / 161 = 0
    16'b01111001_10100010 : OUT <= 0;  //121 / 162 = 0
    16'b01111001_10100011 : OUT <= 0;  //121 / 163 = 0
    16'b01111001_10100100 : OUT <= 0;  //121 / 164 = 0
    16'b01111001_10100101 : OUT <= 0;  //121 / 165 = 0
    16'b01111001_10100110 : OUT <= 0;  //121 / 166 = 0
    16'b01111001_10100111 : OUT <= 0;  //121 / 167 = 0
    16'b01111001_10101000 : OUT <= 0;  //121 / 168 = 0
    16'b01111001_10101001 : OUT <= 0;  //121 / 169 = 0
    16'b01111001_10101010 : OUT <= 0;  //121 / 170 = 0
    16'b01111001_10101011 : OUT <= 0;  //121 / 171 = 0
    16'b01111001_10101100 : OUT <= 0;  //121 / 172 = 0
    16'b01111001_10101101 : OUT <= 0;  //121 / 173 = 0
    16'b01111001_10101110 : OUT <= 0;  //121 / 174 = 0
    16'b01111001_10101111 : OUT <= 0;  //121 / 175 = 0
    16'b01111001_10110000 : OUT <= 0;  //121 / 176 = 0
    16'b01111001_10110001 : OUT <= 0;  //121 / 177 = 0
    16'b01111001_10110010 : OUT <= 0;  //121 / 178 = 0
    16'b01111001_10110011 : OUT <= 0;  //121 / 179 = 0
    16'b01111001_10110100 : OUT <= 0;  //121 / 180 = 0
    16'b01111001_10110101 : OUT <= 0;  //121 / 181 = 0
    16'b01111001_10110110 : OUT <= 0;  //121 / 182 = 0
    16'b01111001_10110111 : OUT <= 0;  //121 / 183 = 0
    16'b01111001_10111000 : OUT <= 0;  //121 / 184 = 0
    16'b01111001_10111001 : OUT <= 0;  //121 / 185 = 0
    16'b01111001_10111010 : OUT <= 0;  //121 / 186 = 0
    16'b01111001_10111011 : OUT <= 0;  //121 / 187 = 0
    16'b01111001_10111100 : OUT <= 0;  //121 / 188 = 0
    16'b01111001_10111101 : OUT <= 0;  //121 / 189 = 0
    16'b01111001_10111110 : OUT <= 0;  //121 / 190 = 0
    16'b01111001_10111111 : OUT <= 0;  //121 / 191 = 0
    16'b01111001_11000000 : OUT <= 0;  //121 / 192 = 0
    16'b01111001_11000001 : OUT <= 0;  //121 / 193 = 0
    16'b01111001_11000010 : OUT <= 0;  //121 / 194 = 0
    16'b01111001_11000011 : OUT <= 0;  //121 / 195 = 0
    16'b01111001_11000100 : OUT <= 0;  //121 / 196 = 0
    16'b01111001_11000101 : OUT <= 0;  //121 / 197 = 0
    16'b01111001_11000110 : OUT <= 0;  //121 / 198 = 0
    16'b01111001_11000111 : OUT <= 0;  //121 / 199 = 0
    16'b01111001_11001000 : OUT <= 0;  //121 / 200 = 0
    16'b01111001_11001001 : OUT <= 0;  //121 / 201 = 0
    16'b01111001_11001010 : OUT <= 0;  //121 / 202 = 0
    16'b01111001_11001011 : OUT <= 0;  //121 / 203 = 0
    16'b01111001_11001100 : OUT <= 0;  //121 / 204 = 0
    16'b01111001_11001101 : OUT <= 0;  //121 / 205 = 0
    16'b01111001_11001110 : OUT <= 0;  //121 / 206 = 0
    16'b01111001_11001111 : OUT <= 0;  //121 / 207 = 0
    16'b01111001_11010000 : OUT <= 0;  //121 / 208 = 0
    16'b01111001_11010001 : OUT <= 0;  //121 / 209 = 0
    16'b01111001_11010010 : OUT <= 0;  //121 / 210 = 0
    16'b01111001_11010011 : OUT <= 0;  //121 / 211 = 0
    16'b01111001_11010100 : OUT <= 0;  //121 / 212 = 0
    16'b01111001_11010101 : OUT <= 0;  //121 / 213 = 0
    16'b01111001_11010110 : OUT <= 0;  //121 / 214 = 0
    16'b01111001_11010111 : OUT <= 0;  //121 / 215 = 0
    16'b01111001_11011000 : OUT <= 0;  //121 / 216 = 0
    16'b01111001_11011001 : OUT <= 0;  //121 / 217 = 0
    16'b01111001_11011010 : OUT <= 0;  //121 / 218 = 0
    16'b01111001_11011011 : OUT <= 0;  //121 / 219 = 0
    16'b01111001_11011100 : OUT <= 0;  //121 / 220 = 0
    16'b01111001_11011101 : OUT <= 0;  //121 / 221 = 0
    16'b01111001_11011110 : OUT <= 0;  //121 / 222 = 0
    16'b01111001_11011111 : OUT <= 0;  //121 / 223 = 0
    16'b01111001_11100000 : OUT <= 0;  //121 / 224 = 0
    16'b01111001_11100001 : OUT <= 0;  //121 / 225 = 0
    16'b01111001_11100010 : OUT <= 0;  //121 / 226 = 0
    16'b01111001_11100011 : OUT <= 0;  //121 / 227 = 0
    16'b01111001_11100100 : OUT <= 0;  //121 / 228 = 0
    16'b01111001_11100101 : OUT <= 0;  //121 / 229 = 0
    16'b01111001_11100110 : OUT <= 0;  //121 / 230 = 0
    16'b01111001_11100111 : OUT <= 0;  //121 / 231 = 0
    16'b01111001_11101000 : OUT <= 0;  //121 / 232 = 0
    16'b01111001_11101001 : OUT <= 0;  //121 / 233 = 0
    16'b01111001_11101010 : OUT <= 0;  //121 / 234 = 0
    16'b01111001_11101011 : OUT <= 0;  //121 / 235 = 0
    16'b01111001_11101100 : OUT <= 0;  //121 / 236 = 0
    16'b01111001_11101101 : OUT <= 0;  //121 / 237 = 0
    16'b01111001_11101110 : OUT <= 0;  //121 / 238 = 0
    16'b01111001_11101111 : OUT <= 0;  //121 / 239 = 0
    16'b01111001_11110000 : OUT <= 0;  //121 / 240 = 0
    16'b01111001_11110001 : OUT <= 0;  //121 / 241 = 0
    16'b01111001_11110010 : OUT <= 0;  //121 / 242 = 0
    16'b01111001_11110011 : OUT <= 0;  //121 / 243 = 0
    16'b01111001_11110100 : OUT <= 0;  //121 / 244 = 0
    16'b01111001_11110101 : OUT <= 0;  //121 / 245 = 0
    16'b01111001_11110110 : OUT <= 0;  //121 / 246 = 0
    16'b01111001_11110111 : OUT <= 0;  //121 / 247 = 0
    16'b01111001_11111000 : OUT <= 0;  //121 / 248 = 0
    16'b01111001_11111001 : OUT <= 0;  //121 / 249 = 0
    16'b01111001_11111010 : OUT <= 0;  //121 / 250 = 0
    16'b01111001_11111011 : OUT <= 0;  //121 / 251 = 0
    16'b01111001_11111100 : OUT <= 0;  //121 / 252 = 0
    16'b01111001_11111101 : OUT <= 0;  //121 / 253 = 0
    16'b01111001_11111110 : OUT <= 0;  //121 / 254 = 0
    16'b01111001_11111111 : OUT <= 0;  //121 / 255 = 0
    16'b01111010_00000000 : OUT <= 0;  //122 / 0 = 0
    16'b01111010_00000001 : OUT <= 122;  //122 / 1 = 122
    16'b01111010_00000010 : OUT <= 61;  //122 / 2 = 61
    16'b01111010_00000011 : OUT <= 40;  //122 / 3 = 40
    16'b01111010_00000100 : OUT <= 30;  //122 / 4 = 30
    16'b01111010_00000101 : OUT <= 24;  //122 / 5 = 24
    16'b01111010_00000110 : OUT <= 20;  //122 / 6 = 20
    16'b01111010_00000111 : OUT <= 17;  //122 / 7 = 17
    16'b01111010_00001000 : OUT <= 15;  //122 / 8 = 15
    16'b01111010_00001001 : OUT <= 13;  //122 / 9 = 13
    16'b01111010_00001010 : OUT <= 12;  //122 / 10 = 12
    16'b01111010_00001011 : OUT <= 11;  //122 / 11 = 11
    16'b01111010_00001100 : OUT <= 10;  //122 / 12 = 10
    16'b01111010_00001101 : OUT <= 9;  //122 / 13 = 9
    16'b01111010_00001110 : OUT <= 8;  //122 / 14 = 8
    16'b01111010_00001111 : OUT <= 8;  //122 / 15 = 8
    16'b01111010_00010000 : OUT <= 7;  //122 / 16 = 7
    16'b01111010_00010001 : OUT <= 7;  //122 / 17 = 7
    16'b01111010_00010010 : OUT <= 6;  //122 / 18 = 6
    16'b01111010_00010011 : OUT <= 6;  //122 / 19 = 6
    16'b01111010_00010100 : OUT <= 6;  //122 / 20 = 6
    16'b01111010_00010101 : OUT <= 5;  //122 / 21 = 5
    16'b01111010_00010110 : OUT <= 5;  //122 / 22 = 5
    16'b01111010_00010111 : OUT <= 5;  //122 / 23 = 5
    16'b01111010_00011000 : OUT <= 5;  //122 / 24 = 5
    16'b01111010_00011001 : OUT <= 4;  //122 / 25 = 4
    16'b01111010_00011010 : OUT <= 4;  //122 / 26 = 4
    16'b01111010_00011011 : OUT <= 4;  //122 / 27 = 4
    16'b01111010_00011100 : OUT <= 4;  //122 / 28 = 4
    16'b01111010_00011101 : OUT <= 4;  //122 / 29 = 4
    16'b01111010_00011110 : OUT <= 4;  //122 / 30 = 4
    16'b01111010_00011111 : OUT <= 3;  //122 / 31 = 3
    16'b01111010_00100000 : OUT <= 3;  //122 / 32 = 3
    16'b01111010_00100001 : OUT <= 3;  //122 / 33 = 3
    16'b01111010_00100010 : OUT <= 3;  //122 / 34 = 3
    16'b01111010_00100011 : OUT <= 3;  //122 / 35 = 3
    16'b01111010_00100100 : OUT <= 3;  //122 / 36 = 3
    16'b01111010_00100101 : OUT <= 3;  //122 / 37 = 3
    16'b01111010_00100110 : OUT <= 3;  //122 / 38 = 3
    16'b01111010_00100111 : OUT <= 3;  //122 / 39 = 3
    16'b01111010_00101000 : OUT <= 3;  //122 / 40 = 3
    16'b01111010_00101001 : OUT <= 2;  //122 / 41 = 2
    16'b01111010_00101010 : OUT <= 2;  //122 / 42 = 2
    16'b01111010_00101011 : OUT <= 2;  //122 / 43 = 2
    16'b01111010_00101100 : OUT <= 2;  //122 / 44 = 2
    16'b01111010_00101101 : OUT <= 2;  //122 / 45 = 2
    16'b01111010_00101110 : OUT <= 2;  //122 / 46 = 2
    16'b01111010_00101111 : OUT <= 2;  //122 / 47 = 2
    16'b01111010_00110000 : OUT <= 2;  //122 / 48 = 2
    16'b01111010_00110001 : OUT <= 2;  //122 / 49 = 2
    16'b01111010_00110010 : OUT <= 2;  //122 / 50 = 2
    16'b01111010_00110011 : OUT <= 2;  //122 / 51 = 2
    16'b01111010_00110100 : OUT <= 2;  //122 / 52 = 2
    16'b01111010_00110101 : OUT <= 2;  //122 / 53 = 2
    16'b01111010_00110110 : OUT <= 2;  //122 / 54 = 2
    16'b01111010_00110111 : OUT <= 2;  //122 / 55 = 2
    16'b01111010_00111000 : OUT <= 2;  //122 / 56 = 2
    16'b01111010_00111001 : OUT <= 2;  //122 / 57 = 2
    16'b01111010_00111010 : OUT <= 2;  //122 / 58 = 2
    16'b01111010_00111011 : OUT <= 2;  //122 / 59 = 2
    16'b01111010_00111100 : OUT <= 2;  //122 / 60 = 2
    16'b01111010_00111101 : OUT <= 2;  //122 / 61 = 2
    16'b01111010_00111110 : OUT <= 1;  //122 / 62 = 1
    16'b01111010_00111111 : OUT <= 1;  //122 / 63 = 1
    16'b01111010_01000000 : OUT <= 1;  //122 / 64 = 1
    16'b01111010_01000001 : OUT <= 1;  //122 / 65 = 1
    16'b01111010_01000010 : OUT <= 1;  //122 / 66 = 1
    16'b01111010_01000011 : OUT <= 1;  //122 / 67 = 1
    16'b01111010_01000100 : OUT <= 1;  //122 / 68 = 1
    16'b01111010_01000101 : OUT <= 1;  //122 / 69 = 1
    16'b01111010_01000110 : OUT <= 1;  //122 / 70 = 1
    16'b01111010_01000111 : OUT <= 1;  //122 / 71 = 1
    16'b01111010_01001000 : OUT <= 1;  //122 / 72 = 1
    16'b01111010_01001001 : OUT <= 1;  //122 / 73 = 1
    16'b01111010_01001010 : OUT <= 1;  //122 / 74 = 1
    16'b01111010_01001011 : OUT <= 1;  //122 / 75 = 1
    16'b01111010_01001100 : OUT <= 1;  //122 / 76 = 1
    16'b01111010_01001101 : OUT <= 1;  //122 / 77 = 1
    16'b01111010_01001110 : OUT <= 1;  //122 / 78 = 1
    16'b01111010_01001111 : OUT <= 1;  //122 / 79 = 1
    16'b01111010_01010000 : OUT <= 1;  //122 / 80 = 1
    16'b01111010_01010001 : OUT <= 1;  //122 / 81 = 1
    16'b01111010_01010010 : OUT <= 1;  //122 / 82 = 1
    16'b01111010_01010011 : OUT <= 1;  //122 / 83 = 1
    16'b01111010_01010100 : OUT <= 1;  //122 / 84 = 1
    16'b01111010_01010101 : OUT <= 1;  //122 / 85 = 1
    16'b01111010_01010110 : OUT <= 1;  //122 / 86 = 1
    16'b01111010_01010111 : OUT <= 1;  //122 / 87 = 1
    16'b01111010_01011000 : OUT <= 1;  //122 / 88 = 1
    16'b01111010_01011001 : OUT <= 1;  //122 / 89 = 1
    16'b01111010_01011010 : OUT <= 1;  //122 / 90 = 1
    16'b01111010_01011011 : OUT <= 1;  //122 / 91 = 1
    16'b01111010_01011100 : OUT <= 1;  //122 / 92 = 1
    16'b01111010_01011101 : OUT <= 1;  //122 / 93 = 1
    16'b01111010_01011110 : OUT <= 1;  //122 / 94 = 1
    16'b01111010_01011111 : OUT <= 1;  //122 / 95 = 1
    16'b01111010_01100000 : OUT <= 1;  //122 / 96 = 1
    16'b01111010_01100001 : OUT <= 1;  //122 / 97 = 1
    16'b01111010_01100010 : OUT <= 1;  //122 / 98 = 1
    16'b01111010_01100011 : OUT <= 1;  //122 / 99 = 1
    16'b01111010_01100100 : OUT <= 1;  //122 / 100 = 1
    16'b01111010_01100101 : OUT <= 1;  //122 / 101 = 1
    16'b01111010_01100110 : OUT <= 1;  //122 / 102 = 1
    16'b01111010_01100111 : OUT <= 1;  //122 / 103 = 1
    16'b01111010_01101000 : OUT <= 1;  //122 / 104 = 1
    16'b01111010_01101001 : OUT <= 1;  //122 / 105 = 1
    16'b01111010_01101010 : OUT <= 1;  //122 / 106 = 1
    16'b01111010_01101011 : OUT <= 1;  //122 / 107 = 1
    16'b01111010_01101100 : OUT <= 1;  //122 / 108 = 1
    16'b01111010_01101101 : OUT <= 1;  //122 / 109 = 1
    16'b01111010_01101110 : OUT <= 1;  //122 / 110 = 1
    16'b01111010_01101111 : OUT <= 1;  //122 / 111 = 1
    16'b01111010_01110000 : OUT <= 1;  //122 / 112 = 1
    16'b01111010_01110001 : OUT <= 1;  //122 / 113 = 1
    16'b01111010_01110010 : OUT <= 1;  //122 / 114 = 1
    16'b01111010_01110011 : OUT <= 1;  //122 / 115 = 1
    16'b01111010_01110100 : OUT <= 1;  //122 / 116 = 1
    16'b01111010_01110101 : OUT <= 1;  //122 / 117 = 1
    16'b01111010_01110110 : OUT <= 1;  //122 / 118 = 1
    16'b01111010_01110111 : OUT <= 1;  //122 / 119 = 1
    16'b01111010_01111000 : OUT <= 1;  //122 / 120 = 1
    16'b01111010_01111001 : OUT <= 1;  //122 / 121 = 1
    16'b01111010_01111010 : OUT <= 1;  //122 / 122 = 1
    16'b01111010_01111011 : OUT <= 0;  //122 / 123 = 0
    16'b01111010_01111100 : OUT <= 0;  //122 / 124 = 0
    16'b01111010_01111101 : OUT <= 0;  //122 / 125 = 0
    16'b01111010_01111110 : OUT <= 0;  //122 / 126 = 0
    16'b01111010_01111111 : OUT <= 0;  //122 / 127 = 0
    16'b01111010_10000000 : OUT <= 0;  //122 / 128 = 0
    16'b01111010_10000001 : OUT <= 0;  //122 / 129 = 0
    16'b01111010_10000010 : OUT <= 0;  //122 / 130 = 0
    16'b01111010_10000011 : OUT <= 0;  //122 / 131 = 0
    16'b01111010_10000100 : OUT <= 0;  //122 / 132 = 0
    16'b01111010_10000101 : OUT <= 0;  //122 / 133 = 0
    16'b01111010_10000110 : OUT <= 0;  //122 / 134 = 0
    16'b01111010_10000111 : OUT <= 0;  //122 / 135 = 0
    16'b01111010_10001000 : OUT <= 0;  //122 / 136 = 0
    16'b01111010_10001001 : OUT <= 0;  //122 / 137 = 0
    16'b01111010_10001010 : OUT <= 0;  //122 / 138 = 0
    16'b01111010_10001011 : OUT <= 0;  //122 / 139 = 0
    16'b01111010_10001100 : OUT <= 0;  //122 / 140 = 0
    16'b01111010_10001101 : OUT <= 0;  //122 / 141 = 0
    16'b01111010_10001110 : OUT <= 0;  //122 / 142 = 0
    16'b01111010_10001111 : OUT <= 0;  //122 / 143 = 0
    16'b01111010_10010000 : OUT <= 0;  //122 / 144 = 0
    16'b01111010_10010001 : OUT <= 0;  //122 / 145 = 0
    16'b01111010_10010010 : OUT <= 0;  //122 / 146 = 0
    16'b01111010_10010011 : OUT <= 0;  //122 / 147 = 0
    16'b01111010_10010100 : OUT <= 0;  //122 / 148 = 0
    16'b01111010_10010101 : OUT <= 0;  //122 / 149 = 0
    16'b01111010_10010110 : OUT <= 0;  //122 / 150 = 0
    16'b01111010_10010111 : OUT <= 0;  //122 / 151 = 0
    16'b01111010_10011000 : OUT <= 0;  //122 / 152 = 0
    16'b01111010_10011001 : OUT <= 0;  //122 / 153 = 0
    16'b01111010_10011010 : OUT <= 0;  //122 / 154 = 0
    16'b01111010_10011011 : OUT <= 0;  //122 / 155 = 0
    16'b01111010_10011100 : OUT <= 0;  //122 / 156 = 0
    16'b01111010_10011101 : OUT <= 0;  //122 / 157 = 0
    16'b01111010_10011110 : OUT <= 0;  //122 / 158 = 0
    16'b01111010_10011111 : OUT <= 0;  //122 / 159 = 0
    16'b01111010_10100000 : OUT <= 0;  //122 / 160 = 0
    16'b01111010_10100001 : OUT <= 0;  //122 / 161 = 0
    16'b01111010_10100010 : OUT <= 0;  //122 / 162 = 0
    16'b01111010_10100011 : OUT <= 0;  //122 / 163 = 0
    16'b01111010_10100100 : OUT <= 0;  //122 / 164 = 0
    16'b01111010_10100101 : OUT <= 0;  //122 / 165 = 0
    16'b01111010_10100110 : OUT <= 0;  //122 / 166 = 0
    16'b01111010_10100111 : OUT <= 0;  //122 / 167 = 0
    16'b01111010_10101000 : OUT <= 0;  //122 / 168 = 0
    16'b01111010_10101001 : OUT <= 0;  //122 / 169 = 0
    16'b01111010_10101010 : OUT <= 0;  //122 / 170 = 0
    16'b01111010_10101011 : OUT <= 0;  //122 / 171 = 0
    16'b01111010_10101100 : OUT <= 0;  //122 / 172 = 0
    16'b01111010_10101101 : OUT <= 0;  //122 / 173 = 0
    16'b01111010_10101110 : OUT <= 0;  //122 / 174 = 0
    16'b01111010_10101111 : OUT <= 0;  //122 / 175 = 0
    16'b01111010_10110000 : OUT <= 0;  //122 / 176 = 0
    16'b01111010_10110001 : OUT <= 0;  //122 / 177 = 0
    16'b01111010_10110010 : OUT <= 0;  //122 / 178 = 0
    16'b01111010_10110011 : OUT <= 0;  //122 / 179 = 0
    16'b01111010_10110100 : OUT <= 0;  //122 / 180 = 0
    16'b01111010_10110101 : OUT <= 0;  //122 / 181 = 0
    16'b01111010_10110110 : OUT <= 0;  //122 / 182 = 0
    16'b01111010_10110111 : OUT <= 0;  //122 / 183 = 0
    16'b01111010_10111000 : OUT <= 0;  //122 / 184 = 0
    16'b01111010_10111001 : OUT <= 0;  //122 / 185 = 0
    16'b01111010_10111010 : OUT <= 0;  //122 / 186 = 0
    16'b01111010_10111011 : OUT <= 0;  //122 / 187 = 0
    16'b01111010_10111100 : OUT <= 0;  //122 / 188 = 0
    16'b01111010_10111101 : OUT <= 0;  //122 / 189 = 0
    16'b01111010_10111110 : OUT <= 0;  //122 / 190 = 0
    16'b01111010_10111111 : OUT <= 0;  //122 / 191 = 0
    16'b01111010_11000000 : OUT <= 0;  //122 / 192 = 0
    16'b01111010_11000001 : OUT <= 0;  //122 / 193 = 0
    16'b01111010_11000010 : OUT <= 0;  //122 / 194 = 0
    16'b01111010_11000011 : OUT <= 0;  //122 / 195 = 0
    16'b01111010_11000100 : OUT <= 0;  //122 / 196 = 0
    16'b01111010_11000101 : OUT <= 0;  //122 / 197 = 0
    16'b01111010_11000110 : OUT <= 0;  //122 / 198 = 0
    16'b01111010_11000111 : OUT <= 0;  //122 / 199 = 0
    16'b01111010_11001000 : OUT <= 0;  //122 / 200 = 0
    16'b01111010_11001001 : OUT <= 0;  //122 / 201 = 0
    16'b01111010_11001010 : OUT <= 0;  //122 / 202 = 0
    16'b01111010_11001011 : OUT <= 0;  //122 / 203 = 0
    16'b01111010_11001100 : OUT <= 0;  //122 / 204 = 0
    16'b01111010_11001101 : OUT <= 0;  //122 / 205 = 0
    16'b01111010_11001110 : OUT <= 0;  //122 / 206 = 0
    16'b01111010_11001111 : OUT <= 0;  //122 / 207 = 0
    16'b01111010_11010000 : OUT <= 0;  //122 / 208 = 0
    16'b01111010_11010001 : OUT <= 0;  //122 / 209 = 0
    16'b01111010_11010010 : OUT <= 0;  //122 / 210 = 0
    16'b01111010_11010011 : OUT <= 0;  //122 / 211 = 0
    16'b01111010_11010100 : OUT <= 0;  //122 / 212 = 0
    16'b01111010_11010101 : OUT <= 0;  //122 / 213 = 0
    16'b01111010_11010110 : OUT <= 0;  //122 / 214 = 0
    16'b01111010_11010111 : OUT <= 0;  //122 / 215 = 0
    16'b01111010_11011000 : OUT <= 0;  //122 / 216 = 0
    16'b01111010_11011001 : OUT <= 0;  //122 / 217 = 0
    16'b01111010_11011010 : OUT <= 0;  //122 / 218 = 0
    16'b01111010_11011011 : OUT <= 0;  //122 / 219 = 0
    16'b01111010_11011100 : OUT <= 0;  //122 / 220 = 0
    16'b01111010_11011101 : OUT <= 0;  //122 / 221 = 0
    16'b01111010_11011110 : OUT <= 0;  //122 / 222 = 0
    16'b01111010_11011111 : OUT <= 0;  //122 / 223 = 0
    16'b01111010_11100000 : OUT <= 0;  //122 / 224 = 0
    16'b01111010_11100001 : OUT <= 0;  //122 / 225 = 0
    16'b01111010_11100010 : OUT <= 0;  //122 / 226 = 0
    16'b01111010_11100011 : OUT <= 0;  //122 / 227 = 0
    16'b01111010_11100100 : OUT <= 0;  //122 / 228 = 0
    16'b01111010_11100101 : OUT <= 0;  //122 / 229 = 0
    16'b01111010_11100110 : OUT <= 0;  //122 / 230 = 0
    16'b01111010_11100111 : OUT <= 0;  //122 / 231 = 0
    16'b01111010_11101000 : OUT <= 0;  //122 / 232 = 0
    16'b01111010_11101001 : OUT <= 0;  //122 / 233 = 0
    16'b01111010_11101010 : OUT <= 0;  //122 / 234 = 0
    16'b01111010_11101011 : OUT <= 0;  //122 / 235 = 0
    16'b01111010_11101100 : OUT <= 0;  //122 / 236 = 0
    16'b01111010_11101101 : OUT <= 0;  //122 / 237 = 0
    16'b01111010_11101110 : OUT <= 0;  //122 / 238 = 0
    16'b01111010_11101111 : OUT <= 0;  //122 / 239 = 0
    16'b01111010_11110000 : OUT <= 0;  //122 / 240 = 0
    16'b01111010_11110001 : OUT <= 0;  //122 / 241 = 0
    16'b01111010_11110010 : OUT <= 0;  //122 / 242 = 0
    16'b01111010_11110011 : OUT <= 0;  //122 / 243 = 0
    16'b01111010_11110100 : OUT <= 0;  //122 / 244 = 0
    16'b01111010_11110101 : OUT <= 0;  //122 / 245 = 0
    16'b01111010_11110110 : OUT <= 0;  //122 / 246 = 0
    16'b01111010_11110111 : OUT <= 0;  //122 / 247 = 0
    16'b01111010_11111000 : OUT <= 0;  //122 / 248 = 0
    16'b01111010_11111001 : OUT <= 0;  //122 / 249 = 0
    16'b01111010_11111010 : OUT <= 0;  //122 / 250 = 0
    16'b01111010_11111011 : OUT <= 0;  //122 / 251 = 0
    16'b01111010_11111100 : OUT <= 0;  //122 / 252 = 0
    16'b01111010_11111101 : OUT <= 0;  //122 / 253 = 0
    16'b01111010_11111110 : OUT <= 0;  //122 / 254 = 0
    16'b01111010_11111111 : OUT <= 0;  //122 / 255 = 0
    16'b01111011_00000000 : OUT <= 0;  //123 / 0 = 0
    16'b01111011_00000001 : OUT <= 123;  //123 / 1 = 123
    16'b01111011_00000010 : OUT <= 61;  //123 / 2 = 61
    16'b01111011_00000011 : OUT <= 41;  //123 / 3 = 41
    16'b01111011_00000100 : OUT <= 30;  //123 / 4 = 30
    16'b01111011_00000101 : OUT <= 24;  //123 / 5 = 24
    16'b01111011_00000110 : OUT <= 20;  //123 / 6 = 20
    16'b01111011_00000111 : OUT <= 17;  //123 / 7 = 17
    16'b01111011_00001000 : OUT <= 15;  //123 / 8 = 15
    16'b01111011_00001001 : OUT <= 13;  //123 / 9 = 13
    16'b01111011_00001010 : OUT <= 12;  //123 / 10 = 12
    16'b01111011_00001011 : OUT <= 11;  //123 / 11 = 11
    16'b01111011_00001100 : OUT <= 10;  //123 / 12 = 10
    16'b01111011_00001101 : OUT <= 9;  //123 / 13 = 9
    16'b01111011_00001110 : OUT <= 8;  //123 / 14 = 8
    16'b01111011_00001111 : OUT <= 8;  //123 / 15 = 8
    16'b01111011_00010000 : OUT <= 7;  //123 / 16 = 7
    16'b01111011_00010001 : OUT <= 7;  //123 / 17 = 7
    16'b01111011_00010010 : OUT <= 6;  //123 / 18 = 6
    16'b01111011_00010011 : OUT <= 6;  //123 / 19 = 6
    16'b01111011_00010100 : OUT <= 6;  //123 / 20 = 6
    16'b01111011_00010101 : OUT <= 5;  //123 / 21 = 5
    16'b01111011_00010110 : OUT <= 5;  //123 / 22 = 5
    16'b01111011_00010111 : OUT <= 5;  //123 / 23 = 5
    16'b01111011_00011000 : OUT <= 5;  //123 / 24 = 5
    16'b01111011_00011001 : OUT <= 4;  //123 / 25 = 4
    16'b01111011_00011010 : OUT <= 4;  //123 / 26 = 4
    16'b01111011_00011011 : OUT <= 4;  //123 / 27 = 4
    16'b01111011_00011100 : OUT <= 4;  //123 / 28 = 4
    16'b01111011_00011101 : OUT <= 4;  //123 / 29 = 4
    16'b01111011_00011110 : OUT <= 4;  //123 / 30 = 4
    16'b01111011_00011111 : OUT <= 3;  //123 / 31 = 3
    16'b01111011_00100000 : OUT <= 3;  //123 / 32 = 3
    16'b01111011_00100001 : OUT <= 3;  //123 / 33 = 3
    16'b01111011_00100010 : OUT <= 3;  //123 / 34 = 3
    16'b01111011_00100011 : OUT <= 3;  //123 / 35 = 3
    16'b01111011_00100100 : OUT <= 3;  //123 / 36 = 3
    16'b01111011_00100101 : OUT <= 3;  //123 / 37 = 3
    16'b01111011_00100110 : OUT <= 3;  //123 / 38 = 3
    16'b01111011_00100111 : OUT <= 3;  //123 / 39 = 3
    16'b01111011_00101000 : OUT <= 3;  //123 / 40 = 3
    16'b01111011_00101001 : OUT <= 3;  //123 / 41 = 3
    16'b01111011_00101010 : OUT <= 2;  //123 / 42 = 2
    16'b01111011_00101011 : OUT <= 2;  //123 / 43 = 2
    16'b01111011_00101100 : OUT <= 2;  //123 / 44 = 2
    16'b01111011_00101101 : OUT <= 2;  //123 / 45 = 2
    16'b01111011_00101110 : OUT <= 2;  //123 / 46 = 2
    16'b01111011_00101111 : OUT <= 2;  //123 / 47 = 2
    16'b01111011_00110000 : OUT <= 2;  //123 / 48 = 2
    16'b01111011_00110001 : OUT <= 2;  //123 / 49 = 2
    16'b01111011_00110010 : OUT <= 2;  //123 / 50 = 2
    16'b01111011_00110011 : OUT <= 2;  //123 / 51 = 2
    16'b01111011_00110100 : OUT <= 2;  //123 / 52 = 2
    16'b01111011_00110101 : OUT <= 2;  //123 / 53 = 2
    16'b01111011_00110110 : OUT <= 2;  //123 / 54 = 2
    16'b01111011_00110111 : OUT <= 2;  //123 / 55 = 2
    16'b01111011_00111000 : OUT <= 2;  //123 / 56 = 2
    16'b01111011_00111001 : OUT <= 2;  //123 / 57 = 2
    16'b01111011_00111010 : OUT <= 2;  //123 / 58 = 2
    16'b01111011_00111011 : OUT <= 2;  //123 / 59 = 2
    16'b01111011_00111100 : OUT <= 2;  //123 / 60 = 2
    16'b01111011_00111101 : OUT <= 2;  //123 / 61 = 2
    16'b01111011_00111110 : OUT <= 1;  //123 / 62 = 1
    16'b01111011_00111111 : OUT <= 1;  //123 / 63 = 1
    16'b01111011_01000000 : OUT <= 1;  //123 / 64 = 1
    16'b01111011_01000001 : OUT <= 1;  //123 / 65 = 1
    16'b01111011_01000010 : OUT <= 1;  //123 / 66 = 1
    16'b01111011_01000011 : OUT <= 1;  //123 / 67 = 1
    16'b01111011_01000100 : OUT <= 1;  //123 / 68 = 1
    16'b01111011_01000101 : OUT <= 1;  //123 / 69 = 1
    16'b01111011_01000110 : OUT <= 1;  //123 / 70 = 1
    16'b01111011_01000111 : OUT <= 1;  //123 / 71 = 1
    16'b01111011_01001000 : OUT <= 1;  //123 / 72 = 1
    16'b01111011_01001001 : OUT <= 1;  //123 / 73 = 1
    16'b01111011_01001010 : OUT <= 1;  //123 / 74 = 1
    16'b01111011_01001011 : OUT <= 1;  //123 / 75 = 1
    16'b01111011_01001100 : OUT <= 1;  //123 / 76 = 1
    16'b01111011_01001101 : OUT <= 1;  //123 / 77 = 1
    16'b01111011_01001110 : OUT <= 1;  //123 / 78 = 1
    16'b01111011_01001111 : OUT <= 1;  //123 / 79 = 1
    16'b01111011_01010000 : OUT <= 1;  //123 / 80 = 1
    16'b01111011_01010001 : OUT <= 1;  //123 / 81 = 1
    16'b01111011_01010010 : OUT <= 1;  //123 / 82 = 1
    16'b01111011_01010011 : OUT <= 1;  //123 / 83 = 1
    16'b01111011_01010100 : OUT <= 1;  //123 / 84 = 1
    16'b01111011_01010101 : OUT <= 1;  //123 / 85 = 1
    16'b01111011_01010110 : OUT <= 1;  //123 / 86 = 1
    16'b01111011_01010111 : OUT <= 1;  //123 / 87 = 1
    16'b01111011_01011000 : OUT <= 1;  //123 / 88 = 1
    16'b01111011_01011001 : OUT <= 1;  //123 / 89 = 1
    16'b01111011_01011010 : OUT <= 1;  //123 / 90 = 1
    16'b01111011_01011011 : OUT <= 1;  //123 / 91 = 1
    16'b01111011_01011100 : OUT <= 1;  //123 / 92 = 1
    16'b01111011_01011101 : OUT <= 1;  //123 / 93 = 1
    16'b01111011_01011110 : OUT <= 1;  //123 / 94 = 1
    16'b01111011_01011111 : OUT <= 1;  //123 / 95 = 1
    16'b01111011_01100000 : OUT <= 1;  //123 / 96 = 1
    16'b01111011_01100001 : OUT <= 1;  //123 / 97 = 1
    16'b01111011_01100010 : OUT <= 1;  //123 / 98 = 1
    16'b01111011_01100011 : OUT <= 1;  //123 / 99 = 1
    16'b01111011_01100100 : OUT <= 1;  //123 / 100 = 1
    16'b01111011_01100101 : OUT <= 1;  //123 / 101 = 1
    16'b01111011_01100110 : OUT <= 1;  //123 / 102 = 1
    16'b01111011_01100111 : OUT <= 1;  //123 / 103 = 1
    16'b01111011_01101000 : OUT <= 1;  //123 / 104 = 1
    16'b01111011_01101001 : OUT <= 1;  //123 / 105 = 1
    16'b01111011_01101010 : OUT <= 1;  //123 / 106 = 1
    16'b01111011_01101011 : OUT <= 1;  //123 / 107 = 1
    16'b01111011_01101100 : OUT <= 1;  //123 / 108 = 1
    16'b01111011_01101101 : OUT <= 1;  //123 / 109 = 1
    16'b01111011_01101110 : OUT <= 1;  //123 / 110 = 1
    16'b01111011_01101111 : OUT <= 1;  //123 / 111 = 1
    16'b01111011_01110000 : OUT <= 1;  //123 / 112 = 1
    16'b01111011_01110001 : OUT <= 1;  //123 / 113 = 1
    16'b01111011_01110010 : OUT <= 1;  //123 / 114 = 1
    16'b01111011_01110011 : OUT <= 1;  //123 / 115 = 1
    16'b01111011_01110100 : OUT <= 1;  //123 / 116 = 1
    16'b01111011_01110101 : OUT <= 1;  //123 / 117 = 1
    16'b01111011_01110110 : OUT <= 1;  //123 / 118 = 1
    16'b01111011_01110111 : OUT <= 1;  //123 / 119 = 1
    16'b01111011_01111000 : OUT <= 1;  //123 / 120 = 1
    16'b01111011_01111001 : OUT <= 1;  //123 / 121 = 1
    16'b01111011_01111010 : OUT <= 1;  //123 / 122 = 1
    16'b01111011_01111011 : OUT <= 1;  //123 / 123 = 1
    16'b01111011_01111100 : OUT <= 0;  //123 / 124 = 0
    16'b01111011_01111101 : OUT <= 0;  //123 / 125 = 0
    16'b01111011_01111110 : OUT <= 0;  //123 / 126 = 0
    16'b01111011_01111111 : OUT <= 0;  //123 / 127 = 0
    16'b01111011_10000000 : OUT <= 0;  //123 / 128 = 0
    16'b01111011_10000001 : OUT <= 0;  //123 / 129 = 0
    16'b01111011_10000010 : OUT <= 0;  //123 / 130 = 0
    16'b01111011_10000011 : OUT <= 0;  //123 / 131 = 0
    16'b01111011_10000100 : OUT <= 0;  //123 / 132 = 0
    16'b01111011_10000101 : OUT <= 0;  //123 / 133 = 0
    16'b01111011_10000110 : OUT <= 0;  //123 / 134 = 0
    16'b01111011_10000111 : OUT <= 0;  //123 / 135 = 0
    16'b01111011_10001000 : OUT <= 0;  //123 / 136 = 0
    16'b01111011_10001001 : OUT <= 0;  //123 / 137 = 0
    16'b01111011_10001010 : OUT <= 0;  //123 / 138 = 0
    16'b01111011_10001011 : OUT <= 0;  //123 / 139 = 0
    16'b01111011_10001100 : OUT <= 0;  //123 / 140 = 0
    16'b01111011_10001101 : OUT <= 0;  //123 / 141 = 0
    16'b01111011_10001110 : OUT <= 0;  //123 / 142 = 0
    16'b01111011_10001111 : OUT <= 0;  //123 / 143 = 0
    16'b01111011_10010000 : OUT <= 0;  //123 / 144 = 0
    16'b01111011_10010001 : OUT <= 0;  //123 / 145 = 0
    16'b01111011_10010010 : OUT <= 0;  //123 / 146 = 0
    16'b01111011_10010011 : OUT <= 0;  //123 / 147 = 0
    16'b01111011_10010100 : OUT <= 0;  //123 / 148 = 0
    16'b01111011_10010101 : OUT <= 0;  //123 / 149 = 0
    16'b01111011_10010110 : OUT <= 0;  //123 / 150 = 0
    16'b01111011_10010111 : OUT <= 0;  //123 / 151 = 0
    16'b01111011_10011000 : OUT <= 0;  //123 / 152 = 0
    16'b01111011_10011001 : OUT <= 0;  //123 / 153 = 0
    16'b01111011_10011010 : OUT <= 0;  //123 / 154 = 0
    16'b01111011_10011011 : OUT <= 0;  //123 / 155 = 0
    16'b01111011_10011100 : OUT <= 0;  //123 / 156 = 0
    16'b01111011_10011101 : OUT <= 0;  //123 / 157 = 0
    16'b01111011_10011110 : OUT <= 0;  //123 / 158 = 0
    16'b01111011_10011111 : OUT <= 0;  //123 / 159 = 0
    16'b01111011_10100000 : OUT <= 0;  //123 / 160 = 0
    16'b01111011_10100001 : OUT <= 0;  //123 / 161 = 0
    16'b01111011_10100010 : OUT <= 0;  //123 / 162 = 0
    16'b01111011_10100011 : OUT <= 0;  //123 / 163 = 0
    16'b01111011_10100100 : OUT <= 0;  //123 / 164 = 0
    16'b01111011_10100101 : OUT <= 0;  //123 / 165 = 0
    16'b01111011_10100110 : OUT <= 0;  //123 / 166 = 0
    16'b01111011_10100111 : OUT <= 0;  //123 / 167 = 0
    16'b01111011_10101000 : OUT <= 0;  //123 / 168 = 0
    16'b01111011_10101001 : OUT <= 0;  //123 / 169 = 0
    16'b01111011_10101010 : OUT <= 0;  //123 / 170 = 0
    16'b01111011_10101011 : OUT <= 0;  //123 / 171 = 0
    16'b01111011_10101100 : OUT <= 0;  //123 / 172 = 0
    16'b01111011_10101101 : OUT <= 0;  //123 / 173 = 0
    16'b01111011_10101110 : OUT <= 0;  //123 / 174 = 0
    16'b01111011_10101111 : OUT <= 0;  //123 / 175 = 0
    16'b01111011_10110000 : OUT <= 0;  //123 / 176 = 0
    16'b01111011_10110001 : OUT <= 0;  //123 / 177 = 0
    16'b01111011_10110010 : OUT <= 0;  //123 / 178 = 0
    16'b01111011_10110011 : OUT <= 0;  //123 / 179 = 0
    16'b01111011_10110100 : OUT <= 0;  //123 / 180 = 0
    16'b01111011_10110101 : OUT <= 0;  //123 / 181 = 0
    16'b01111011_10110110 : OUT <= 0;  //123 / 182 = 0
    16'b01111011_10110111 : OUT <= 0;  //123 / 183 = 0
    16'b01111011_10111000 : OUT <= 0;  //123 / 184 = 0
    16'b01111011_10111001 : OUT <= 0;  //123 / 185 = 0
    16'b01111011_10111010 : OUT <= 0;  //123 / 186 = 0
    16'b01111011_10111011 : OUT <= 0;  //123 / 187 = 0
    16'b01111011_10111100 : OUT <= 0;  //123 / 188 = 0
    16'b01111011_10111101 : OUT <= 0;  //123 / 189 = 0
    16'b01111011_10111110 : OUT <= 0;  //123 / 190 = 0
    16'b01111011_10111111 : OUT <= 0;  //123 / 191 = 0
    16'b01111011_11000000 : OUT <= 0;  //123 / 192 = 0
    16'b01111011_11000001 : OUT <= 0;  //123 / 193 = 0
    16'b01111011_11000010 : OUT <= 0;  //123 / 194 = 0
    16'b01111011_11000011 : OUT <= 0;  //123 / 195 = 0
    16'b01111011_11000100 : OUT <= 0;  //123 / 196 = 0
    16'b01111011_11000101 : OUT <= 0;  //123 / 197 = 0
    16'b01111011_11000110 : OUT <= 0;  //123 / 198 = 0
    16'b01111011_11000111 : OUT <= 0;  //123 / 199 = 0
    16'b01111011_11001000 : OUT <= 0;  //123 / 200 = 0
    16'b01111011_11001001 : OUT <= 0;  //123 / 201 = 0
    16'b01111011_11001010 : OUT <= 0;  //123 / 202 = 0
    16'b01111011_11001011 : OUT <= 0;  //123 / 203 = 0
    16'b01111011_11001100 : OUT <= 0;  //123 / 204 = 0
    16'b01111011_11001101 : OUT <= 0;  //123 / 205 = 0
    16'b01111011_11001110 : OUT <= 0;  //123 / 206 = 0
    16'b01111011_11001111 : OUT <= 0;  //123 / 207 = 0
    16'b01111011_11010000 : OUT <= 0;  //123 / 208 = 0
    16'b01111011_11010001 : OUT <= 0;  //123 / 209 = 0
    16'b01111011_11010010 : OUT <= 0;  //123 / 210 = 0
    16'b01111011_11010011 : OUT <= 0;  //123 / 211 = 0
    16'b01111011_11010100 : OUT <= 0;  //123 / 212 = 0
    16'b01111011_11010101 : OUT <= 0;  //123 / 213 = 0
    16'b01111011_11010110 : OUT <= 0;  //123 / 214 = 0
    16'b01111011_11010111 : OUT <= 0;  //123 / 215 = 0
    16'b01111011_11011000 : OUT <= 0;  //123 / 216 = 0
    16'b01111011_11011001 : OUT <= 0;  //123 / 217 = 0
    16'b01111011_11011010 : OUT <= 0;  //123 / 218 = 0
    16'b01111011_11011011 : OUT <= 0;  //123 / 219 = 0
    16'b01111011_11011100 : OUT <= 0;  //123 / 220 = 0
    16'b01111011_11011101 : OUT <= 0;  //123 / 221 = 0
    16'b01111011_11011110 : OUT <= 0;  //123 / 222 = 0
    16'b01111011_11011111 : OUT <= 0;  //123 / 223 = 0
    16'b01111011_11100000 : OUT <= 0;  //123 / 224 = 0
    16'b01111011_11100001 : OUT <= 0;  //123 / 225 = 0
    16'b01111011_11100010 : OUT <= 0;  //123 / 226 = 0
    16'b01111011_11100011 : OUT <= 0;  //123 / 227 = 0
    16'b01111011_11100100 : OUT <= 0;  //123 / 228 = 0
    16'b01111011_11100101 : OUT <= 0;  //123 / 229 = 0
    16'b01111011_11100110 : OUT <= 0;  //123 / 230 = 0
    16'b01111011_11100111 : OUT <= 0;  //123 / 231 = 0
    16'b01111011_11101000 : OUT <= 0;  //123 / 232 = 0
    16'b01111011_11101001 : OUT <= 0;  //123 / 233 = 0
    16'b01111011_11101010 : OUT <= 0;  //123 / 234 = 0
    16'b01111011_11101011 : OUT <= 0;  //123 / 235 = 0
    16'b01111011_11101100 : OUT <= 0;  //123 / 236 = 0
    16'b01111011_11101101 : OUT <= 0;  //123 / 237 = 0
    16'b01111011_11101110 : OUT <= 0;  //123 / 238 = 0
    16'b01111011_11101111 : OUT <= 0;  //123 / 239 = 0
    16'b01111011_11110000 : OUT <= 0;  //123 / 240 = 0
    16'b01111011_11110001 : OUT <= 0;  //123 / 241 = 0
    16'b01111011_11110010 : OUT <= 0;  //123 / 242 = 0
    16'b01111011_11110011 : OUT <= 0;  //123 / 243 = 0
    16'b01111011_11110100 : OUT <= 0;  //123 / 244 = 0
    16'b01111011_11110101 : OUT <= 0;  //123 / 245 = 0
    16'b01111011_11110110 : OUT <= 0;  //123 / 246 = 0
    16'b01111011_11110111 : OUT <= 0;  //123 / 247 = 0
    16'b01111011_11111000 : OUT <= 0;  //123 / 248 = 0
    16'b01111011_11111001 : OUT <= 0;  //123 / 249 = 0
    16'b01111011_11111010 : OUT <= 0;  //123 / 250 = 0
    16'b01111011_11111011 : OUT <= 0;  //123 / 251 = 0
    16'b01111011_11111100 : OUT <= 0;  //123 / 252 = 0
    16'b01111011_11111101 : OUT <= 0;  //123 / 253 = 0
    16'b01111011_11111110 : OUT <= 0;  //123 / 254 = 0
    16'b01111011_11111111 : OUT <= 0;  //123 / 255 = 0
    16'b01111100_00000000 : OUT <= 0;  //124 / 0 = 0
    16'b01111100_00000001 : OUT <= 124;  //124 / 1 = 124
    16'b01111100_00000010 : OUT <= 62;  //124 / 2 = 62
    16'b01111100_00000011 : OUT <= 41;  //124 / 3 = 41
    16'b01111100_00000100 : OUT <= 31;  //124 / 4 = 31
    16'b01111100_00000101 : OUT <= 24;  //124 / 5 = 24
    16'b01111100_00000110 : OUT <= 20;  //124 / 6 = 20
    16'b01111100_00000111 : OUT <= 17;  //124 / 7 = 17
    16'b01111100_00001000 : OUT <= 15;  //124 / 8 = 15
    16'b01111100_00001001 : OUT <= 13;  //124 / 9 = 13
    16'b01111100_00001010 : OUT <= 12;  //124 / 10 = 12
    16'b01111100_00001011 : OUT <= 11;  //124 / 11 = 11
    16'b01111100_00001100 : OUT <= 10;  //124 / 12 = 10
    16'b01111100_00001101 : OUT <= 9;  //124 / 13 = 9
    16'b01111100_00001110 : OUT <= 8;  //124 / 14 = 8
    16'b01111100_00001111 : OUT <= 8;  //124 / 15 = 8
    16'b01111100_00010000 : OUT <= 7;  //124 / 16 = 7
    16'b01111100_00010001 : OUT <= 7;  //124 / 17 = 7
    16'b01111100_00010010 : OUT <= 6;  //124 / 18 = 6
    16'b01111100_00010011 : OUT <= 6;  //124 / 19 = 6
    16'b01111100_00010100 : OUT <= 6;  //124 / 20 = 6
    16'b01111100_00010101 : OUT <= 5;  //124 / 21 = 5
    16'b01111100_00010110 : OUT <= 5;  //124 / 22 = 5
    16'b01111100_00010111 : OUT <= 5;  //124 / 23 = 5
    16'b01111100_00011000 : OUT <= 5;  //124 / 24 = 5
    16'b01111100_00011001 : OUT <= 4;  //124 / 25 = 4
    16'b01111100_00011010 : OUT <= 4;  //124 / 26 = 4
    16'b01111100_00011011 : OUT <= 4;  //124 / 27 = 4
    16'b01111100_00011100 : OUT <= 4;  //124 / 28 = 4
    16'b01111100_00011101 : OUT <= 4;  //124 / 29 = 4
    16'b01111100_00011110 : OUT <= 4;  //124 / 30 = 4
    16'b01111100_00011111 : OUT <= 4;  //124 / 31 = 4
    16'b01111100_00100000 : OUT <= 3;  //124 / 32 = 3
    16'b01111100_00100001 : OUT <= 3;  //124 / 33 = 3
    16'b01111100_00100010 : OUT <= 3;  //124 / 34 = 3
    16'b01111100_00100011 : OUT <= 3;  //124 / 35 = 3
    16'b01111100_00100100 : OUT <= 3;  //124 / 36 = 3
    16'b01111100_00100101 : OUT <= 3;  //124 / 37 = 3
    16'b01111100_00100110 : OUT <= 3;  //124 / 38 = 3
    16'b01111100_00100111 : OUT <= 3;  //124 / 39 = 3
    16'b01111100_00101000 : OUT <= 3;  //124 / 40 = 3
    16'b01111100_00101001 : OUT <= 3;  //124 / 41 = 3
    16'b01111100_00101010 : OUT <= 2;  //124 / 42 = 2
    16'b01111100_00101011 : OUT <= 2;  //124 / 43 = 2
    16'b01111100_00101100 : OUT <= 2;  //124 / 44 = 2
    16'b01111100_00101101 : OUT <= 2;  //124 / 45 = 2
    16'b01111100_00101110 : OUT <= 2;  //124 / 46 = 2
    16'b01111100_00101111 : OUT <= 2;  //124 / 47 = 2
    16'b01111100_00110000 : OUT <= 2;  //124 / 48 = 2
    16'b01111100_00110001 : OUT <= 2;  //124 / 49 = 2
    16'b01111100_00110010 : OUT <= 2;  //124 / 50 = 2
    16'b01111100_00110011 : OUT <= 2;  //124 / 51 = 2
    16'b01111100_00110100 : OUT <= 2;  //124 / 52 = 2
    16'b01111100_00110101 : OUT <= 2;  //124 / 53 = 2
    16'b01111100_00110110 : OUT <= 2;  //124 / 54 = 2
    16'b01111100_00110111 : OUT <= 2;  //124 / 55 = 2
    16'b01111100_00111000 : OUT <= 2;  //124 / 56 = 2
    16'b01111100_00111001 : OUT <= 2;  //124 / 57 = 2
    16'b01111100_00111010 : OUT <= 2;  //124 / 58 = 2
    16'b01111100_00111011 : OUT <= 2;  //124 / 59 = 2
    16'b01111100_00111100 : OUT <= 2;  //124 / 60 = 2
    16'b01111100_00111101 : OUT <= 2;  //124 / 61 = 2
    16'b01111100_00111110 : OUT <= 2;  //124 / 62 = 2
    16'b01111100_00111111 : OUT <= 1;  //124 / 63 = 1
    16'b01111100_01000000 : OUT <= 1;  //124 / 64 = 1
    16'b01111100_01000001 : OUT <= 1;  //124 / 65 = 1
    16'b01111100_01000010 : OUT <= 1;  //124 / 66 = 1
    16'b01111100_01000011 : OUT <= 1;  //124 / 67 = 1
    16'b01111100_01000100 : OUT <= 1;  //124 / 68 = 1
    16'b01111100_01000101 : OUT <= 1;  //124 / 69 = 1
    16'b01111100_01000110 : OUT <= 1;  //124 / 70 = 1
    16'b01111100_01000111 : OUT <= 1;  //124 / 71 = 1
    16'b01111100_01001000 : OUT <= 1;  //124 / 72 = 1
    16'b01111100_01001001 : OUT <= 1;  //124 / 73 = 1
    16'b01111100_01001010 : OUT <= 1;  //124 / 74 = 1
    16'b01111100_01001011 : OUT <= 1;  //124 / 75 = 1
    16'b01111100_01001100 : OUT <= 1;  //124 / 76 = 1
    16'b01111100_01001101 : OUT <= 1;  //124 / 77 = 1
    16'b01111100_01001110 : OUT <= 1;  //124 / 78 = 1
    16'b01111100_01001111 : OUT <= 1;  //124 / 79 = 1
    16'b01111100_01010000 : OUT <= 1;  //124 / 80 = 1
    16'b01111100_01010001 : OUT <= 1;  //124 / 81 = 1
    16'b01111100_01010010 : OUT <= 1;  //124 / 82 = 1
    16'b01111100_01010011 : OUT <= 1;  //124 / 83 = 1
    16'b01111100_01010100 : OUT <= 1;  //124 / 84 = 1
    16'b01111100_01010101 : OUT <= 1;  //124 / 85 = 1
    16'b01111100_01010110 : OUT <= 1;  //124 / 86 = 1
    16'b01111100_01010111 : OUT <= 1;  //124 / 87 = 1
    16'b01111100_01011000 : OUT <= 1;  //124 / 88 = 1
    16'b01111100_01011001 : OUT <= 1;  //124 / 89 = 1
    16'b01111100_01011010 : OUT <= 1;  //124 / 90 = 1
    16'b01111100_01011011 : OUT <= 1;  //124 / 91 = 1
    16'b01111100_01011100 : OUT <= 1;  //124 / 92 = 1
    16'b01111100_01011101 : OUT <= 1;  //124 / 93 = 1
    16'b01111100_01011110 : OUT <= 1;  //124 / 94 = 1
    16'b01111100_01011111 : OUT <= 1;  //124 / 95 = 1
    16'b01111100_01100000 : OUT <= 1;  //124 / 96 = 1
    16'b01111100_01100001 : OUT <= 1;  //124 / 97 = 1
    16'b01111100_01100010 : OUT <= 1;  //124 / 98 = 1
    16'b01111100_01100011 : OUT <= 1;  //124 / 99 = 1
    16'b01111100_01100100 : OUT <= 1;  //124 / 100 = 1
    16'b01111100_01100101 : OUT <= 1;  //124 / 101 = 1
    16'b01111100_01100110 : OUT <= 1;  //124 / 102 = 1
    16'b01111100_01100111 : OUT <= 1;  //124 / 103 = 1
    16'b01111100_01101000 : OUT <= 1;  //124 / 104 = 1
    16'b01111100_01101001 : OUT <= 1;  //124 / 105 = 1
    16'b01111100_01101010 : OUT <= 1;  //124 / 106 = 1
    16'b01111100_01101011 : OUT <= 1;  //124 / 107 = 1
    16'b01111100_01101100 : OUT <= 1;  //124 / 108 = 1
    16'b01111100_01101101 : OUT <= 1;  //124 / 109 = 1
    16'b01111100_01101110 : OUT <= 1;  //124 / 110 = 1
    16'b01111100_01101111 : OUT <= 1;  //124 / 111 = 1
    16'b01111100_01110000 : OUT <= 1;  //124 / 112 = 1
    16'b01111100_01110001 : OUT <= 1;  //124 / 113 = 1
    16'b01111100_01110010 : OUT <= 1;  //124 / 114 = 1
    16'b01111100_01110011 : OUT <= 1;  //124 / 115 = 1
    16'b01111100_01110100 : OUT <= 1;  //124 / 116 = 1
    16'b01111100_01110101 : OUT <= 1;  //124 / 117 = 1
    16'b01111100_01110110 : OUT <= 1;  //124 / 118 = 1
    16'b01111100_01110111 : OUT <= 1;  //124 / 119 = 1
    16'b01111100_01111000 : OUT <= 1;  //124 / 120 = 1
    16'b01111100_01111001 : OUT <= 1;  //124 / 121 = 1
    16'b01111100_01111010 : OUT <= 1;  //124 / 122 = 1
    16'b01111100_01111011 : OUT <= 1;  //124 / 123 = 1
    16'b01111100_01111100 : OUT <= 1;  //124 / 124 = 1
    16'b01111100_01111101 : OUT <= 0;  //124 / 125 = 0
    16'b01111100_01111110 : OUT <= 0;  //124 / 126 = 0
    16'b01111100_01111111 : OUT <= 0;  //124 / 127 = 0
    16'b01111100_10000000 : OUT <= 0;  //124 / 128 = 0
    16'b01111100_10000001 : OUT <= 0;  //124 / 129 = 0
    16'b01111100_10000010 : OUT <= 0;  //124 / 130 = 0
    16'b01111100_10000011 : OUT <= 0;  //124 / 131 = 0
    16'b01111100_10000100 : OUT <= 0;  //124 / 132 = 0
    16'b01111100_10000101 : OUT <= 0;  //124 / 133 = 0
    16'b01111100_10000110 : OUT <= 0;  //124 / 134 = 0
    16'b01111100_10000111 : OUT <= 0;  //124 / 135 = 0
    16'b01111100_10001000 : OUT <= 0;  //124 / 136 = 0
    16'b01111100_10001001 : OUT <= 0;  //124 / 137 = 0
    16'b01111100_10001010 : OUT <= 0;  //124 / 138 = 0
    16'b01111100_10001011 : OUT <= 0;  //124 / 139 = 0
    16'b01111100_10001100 : OUT <= 0;  //124 / 140 = 0
    16'b01111100_10001101 : OUT <= 0;  //124 / 141 = 0
    16'b01111100_10001110 : OUT <= 0;  //124 / 142 = 0
    16'b01111100_10001111 : OUT <= 0;  //124 / 143 = 0
    16'b01111100_10010000 : OUT <= 0;  //124 / 144 = 0
    16'b01111100_10010001 : OUT <= 0;  //124 / 145 = 0
    16'b01111100_10010010 : OUT <= 0;  //124 / 146 = 0
    16'b01111100_10010011 : OUT <= 0;  //124 / 147 = 0
    16'b01111100_10010100 : OUT <= 0;  //124 / 148 = 0
    16'b01111100_10010101 : OUT <= 0;  //124 / 149 = 0
    16'b01111100_10010110 : OUT <= 0;  //124 / 150 = 0
    16'b01111100_10010111 : OUT <= 0;  //124 / 151 = 0
    16'b01111100_10011000 : OUT <= 0;  //124 / 152 = 0
    16'b01111100_10011001 : OUT <= 0;  //124 / 153 = 0
    16'b01111100_10011010 : OUT <= 0;  //124 / 154 = 0
    16'b01111100_10011011 : OUT <= 0;  //124 / 155 = 0
    16'b01111100_10011100 : OUT <= 0;  //124 / 156 = 0
    16'b01111100_10011101 : OUT <= 0;  //124 / 157 = 0
    16'b01111100_10011110 : OUT <= 0;  //124 / 158 = 0
    16'b01111100_10011111 : OUT <= 0;  //124 / 159 = 0
    16'b01111100_10100000 : OUT <= 0;  //124 / 160 = 0
    16'b01111100_10100001 : OUT <= 0;  //124 / 161 = 0
    16'b01111100_10100010 : OUT <= 0;  //124 / 162 = 0
    16'b01111100_10100011 : OUT <= 0;  //124 / 163 = 0
    16'b01111100_10100100 : OUT <= 0;  //124 / 164 = 0
    16'b01111100_10100101 : OUT <= 0;  //124 / 165 = 0
    16'b01111100_10100110 : OUT <= 0;  //124 / 166 = 0
    16'b01111100_10100111 : OUT <= 0;  //124 / 167 = 0
    16'b01111100_10101000 : OUT <= 0;  //124 / 168 = 0
    16'b01111100_10101001 : OUT <= 0;  //124 / 169 = 0
    16'b01111100_10101010 : OUT <= 0;  //124 / 170 = 0
    16'b01111100_10101011 : OUT <= 0;  //124 / 171 = 0
    16'b01111100_10101100 : OUT <= 0;  //124 / 172 = 0
    16'b01111100_10101101 : OUT <= 0;  //124 / 173 = 0
    16'b01111100_10101110 : OUT <= 0;  //124 / 174 = 0
    16'b01111100_10101111 : OUT <= 0;  //124 / 175 = 0
    16'b01111100_10110000 : OUT <= 0;  //124 / 176 = 0
    16'b01111100_10110001 : OUT <= 0;  //124 / 177 = 0
    16'b01111100_10110010 : OUT <= 0;  //124 / 178 = 0
    16'b01111100_10110011 : OUT <= 0;  //124 / 179 = 0
    16'b01111100_10110100 : OUT <= 0;  //124 / 180 = 0
    16'b01111100_10110101 : OUT <= 0;  //124 / 181 = 0
    16'b01111100_10110110 : OUT <= 0;  //124 / 182 = 0
    16'b01111100_10110111 : OUT <= 0;  //124 / 183 = 0
    16'b01111100_10111000 : OUT <= 0;  //124 / 184 = 0
    16'b01111100_10111001 : OUT <= 0;  //124 / 185 = 0
    16'b01111100_10111010 : OUT <= 0;  //124 / 186 = 0
    16'b01111100_10111011 : OUT <= 0;  //124 / 187 = 0
    16'b01111100_10111100 : OUT <= 0;  //124 / 188 = 0
    16'b01111100_10111101 : OUT <= 0;  //124 / 189 = 0
    16'b01111100_10111110 : OUT <= 0;  //124 / 190 = 0
    16'b01111100_10111111 : OUT <= 0;  //124 / 191 = 0
    16'b01111100_11000000 : OUT <= 0;  //124 / 192 = 0
    16'b01111100_11000001 : OUT <= 0;  //124 / 193 = 0
    16'b01111100_11000010 : OUT <= 0;  //124 / 194 = 0
    16'b01111100_11000011 : OUT <= 0;  //124 / 195 = 0
    16'b01111100_11000100 : OUT <= 0;  //124 / 196 = 0
    16'b01111100_11000101 : OUT <= 0;  //124 / 197 = 0
    16'b01111100_11000110 : OUT <= 0;  //124 / 198 = 0
    16'b01111100_11000111 : OUT <= 0;  //124 / 199 = 0
    16'b01111100_11001000 : OUT <= 0;  //124 / 200 = 0
    16'b01111100_11001001 : OUT <= 0;  //124 / 201 = 0
    16'b01111100_11001010 : OUT <= 0;  //124 / 202 = 0
    16'b01111100_11001011 : OUT <= 0;  //124 / 203 = 0
    16'b01111100_11001100 : OUT <= 0;  //124 / 204 = 0
    16'b01111100_11001101 : OUT <= 0;  //124 / 205 = 0
    16'b01111100_11001110 : OUT <= 0;  //124 / 206 = 0
    16'b01111100_11001111 : OUT <= 0;  //124 / 207 = 0
    16'b01111100_11010000 : OUT <= 0;  //124 / 208 = 0
    16'b01111100_11010001 : OUT <= 0;  //124 / 209 = 0
    16'b01111100_11010010 : OUT <= 0;  //124 / 210 = 0
    16'b01111100_11010011 : OUT <= 0;  //124 / 211 = 0
    16'b01111100_11010100 : OUT <= 0;  //124 / 212 = 0
    16'b01111100_11010101 : OUT <= 0;  //124 / 213 = 0
    16'b01111100_11010110 : OUT <= 0;  //124 / 214 = 0
    16'b01111100_11010111 : OUT <= 0;  //124 / 215 = 0
    16'b01111100_11011000 : OUT <= 0;  //124 / 216 = 0
    16'b01111100_11011001 : OUT <= 0;  //124 / 217 = 0
    16'b01111100_11011010 : OUT <= 0;  //124 / 218 = 0
    16'b01111100_11011011 : OUT <= 0;  //124 / 219 = 0
    16'b01111100_11011100 : OUT <= 0;  //124 / 220 = 0
    16'b01111100_11011101 : OUT <= 0;  //124 / 221 = 0
    16'b01111100_11011110 : OUT <= 0;  //124 / 222 = 0
    16'b01111100_11011111 : OUT <= 0;  //124 / 223 = 0
    16'b01111100_11100000 : OUT <= 0;  //124 / 224 = 0
    16'b01111100_11100001 : OUT <= 0;  //124 / 225 = 0
    16'b01111100_11100010 : OUT <= 0;  //124 / 226 = 0
    16'b01111100_11100011 : OUT <= 0;  //124 / 227 = 0
    16'b01111100_11100100 : OUT <= 0;  //124 / 228 = 0
    16'b01111100_11100101 : OUT <= 0;  //124 / 229 = 0
    16'b01111100_11100110 : OUT <= 0;  //124 / 230 = 0
    16'b01111100_11100111 : OUT <= 0;  //124 / 231 = 0
    16'b01111100_11101000 : OUT <= 0;  //124 / 232 = 0
    16'b01111100_11101001 : OUT <= 0;  //124 / 233 = 0
    16'b01111100_11101010 : OUT <= 0;  //124 / 234 = 0
    16'b01111100_11101011 : OUT <= 0;  //124 / 235 = 0
    16'b01111100_11101100 : OUT <= 0;  //124 / 236 = 0
    16'b01111100_11101101 : OUT <= 0;  //124 / 237 = 0
    16'b01111100_11101110 : OUT <= 0;  //124 / 238 = 0
    16'b01111100_11101111 : OUT <= 0;  //124 / 239 = 0
    16'b01111100_11110000 : OUT <= 0;  //124 / 240 = 0
    16'b01111100_11110001 : OUT <= 0;  //124 / 241 = 0
    16'b01111100_11110010 : OUT <= 0;  //124 / 242 = 0
    16'b01111100_11110011 : OUT <= 0;  //124 / 243 = 0
    16'b01111100_11110100 : OUT <= 0;  //124 / 244 = 0
    16'b01111100_11110101 : OUT <= 0;  //124 / 245 = 0
    16'b01111100_11110110 : OUT <= 0;  //124 / 246 = 0
    16'b01111100_11110111 : OUT <= 0;  //124 / 247 = 0
    16'b01111100_11111000 : OUT <= 0;  //124 / 248 = 0
    16'b01111100_11111001 : OUT <= 0;  //124 / 249 = 0
    16'b01111100_11111010 : OUT <= 0;  //124 / 250 = 0
    16'b01111100_11111011 : OUT <= 0;  //124 / 251 = 0
    16'b01111100_11111100 : OUT <= 0;  //124 / 252 = 0
    16'b01111100_11111101 : OUT <= 0;  //124 / 253 = 0
    16'b01111100_11111110 : OUT <= 0;  //124 / 254 = 0
    16'b01111100_11111111 : OUT <= 0;  //124 / 255 = 0
    16'b01111101_00000000 : OUT <= 0;  //125 / 0 = 0
    16'b01111101_00000001 : OUT <= 125;  //125 / 1 = 125
    16'b01111101_00000010 : OUT <= 62;  //125 / 2 = 62
    16'b01111101_00000011 : OUT <= 41;  //125 / 3 = 41
    16'b01111101_00000100 : OUT <= 31;  //125 / 4 = 31
    16'b01111101_00000101 : OUT <= 25;  //125 / 5 = 25
    16'b01111101_00000110 : OUT <= 20;  //125 / 6 = 20
    16'b01111101_00000111 : OUT <= 17;  //125 / 7 = 17
    16'b01111101_00001000 : OUT <= 15;  //125 / 8 = 15
    16'b01111101_00001001 : OUT <= 13;  //125 / 9 = 13
    16'b01111101_00001010 : OUT <= 12;  //125 / 10 = 12
    16'b01111101_00001011 : OUT <= 11;  //125 / 11 = 11
    16'b01111101_00001100 : OUT <= 10;  //125 / 12 = 10
    16'b01111101_00001101 : OUT <= 9;  //125 / 13 = 9
    16'b01111101_00001110 : OUT <= 8;  //125 / 14 = 8
    16'b01111101_00001111 : OUT <= 8;  //125 / 15 = 8
    16'b01111101_00010000 : OUT <= 7;  //125 / 16 = 7
    16'b01111101_00010001 : OUT <= 7;  //125 / 17 = 7
    16'b01111101_00010010 : OUT <= 6;  //125 / 18 = 6
    16'b01111101_00010011 : OUT <= 6;  //125 / 19 = 6
    16'b01111101_00010100 : OUT <= 6;  //125 / 20 = 6
    16'b01111101_00010101 : OUT <= 5;  //125 / 21 = 5
    16'b01111101_00010110 : OUT <= 5;  //125 / 22 = 5
    16'b01111101_00010111 : OUT <= 5;  //125 / 23 = 5
    16'b01111101_00011000 : OUT <= 5;  //125 / 24 = 5
    16'b01111101_00011001 : OUT <= 5;  //125 / 25 = 5
    16'b01111101_00011010 : OUT <= 4;  //125 / 26 = 4
    16'b01111101_00011011 : OUT <= 4;  //125 / 27 = 4
    16'b01111101_00011100 : OUT <= 4;  //125 / 28 = 4
    16'b01111101_00011101 : OUT <= 4;  //125 / 29 = 4
    16'b01111101_00011110 : OUT <= 4;  //125 / 30 = 4
    16'b01111101_00011111 : OUT <= 4;  //125 / 31 = 4
    16'b01111101_00100000 : OUT <= 3;  //125 / 32 = 3
    16'b01111101_00100001 : OUT <= 3;  //125 / 33 = 3
    16'b01111101_00100010 : OUT <= 3;  //125 / 34 = 3
    16'b01111101_00100011 : OUT <= 3;  //125 / 35 = 3
    16'b01111101_00100100 : OUT <= 3;  //125 / 36 = 3
    16'b01111101_00100101 : OUT <= 3;  //125 / 37 = 3
    16'b01111101_00100110 : OUT <= 3;  //125 / 38 = 3
    16'b01111101_00100111 : OUT <= 3;  //125 / 39 = 3
    16'b01111101_00101000 : OUT <= 3;  //125 / 40 = 3
    16'b01111101_00101001 : OUT <= 3;  //125 / 41 = 3
    16'b01111101_00101010 : OUT <= 2;  //125 / 42 = 2
    16'b01111101_00101011 : OUT <= 2;  //125 / 43 = 2
    16'b01111101_00101100 : OUT <= 2;  //125 / 44 = 2
    16'b01111101_00101101 : OUT <= 2;  //125 / 45 = 2
    16'b01111101_00101110 : OUT <= 2;  //125 / 46 = 2
    16'b01111101_00101111 : OUT <= 2;  //125 / 47 = 2
    16'b01111101_00110000 : OUT <= 2;  //125 / 48 = 2
    16'b01111101_00110001 : OUT <= 2;  //125 / 49 = 2
    16'b01111101_00110010 : OUT <= 2;  //125 / 50 = 2
    16'b01111101_00110011 : OUT <= 2;  //125 / 51 = 2
    16'b01111101_00110100 : OUT <= 2;  //125 / 52 = 2
    16'b01111101_00110101 : OUT <= 2;  //125 / 53 = 2
    16'b01111101_00110110 : OUT <= 2;  //125 / 54 = 2
    16'b01111101_00110111 : OUT <= 2;  //125 / 55 = 2
    16'b01111101_00111000 : OUT <= 2;  //125 / 56 = 2
    16'b01111101_00111001 : OUT <= 2;  //125 / 57 = 2
    16'b01111101_00111010 : OUT <= 2;  //125 / 58 = 2
    16'b01111101_00111011 : OUT <= 2;  //125 / 59 = 2
    16'b01111101_00111100 : OUT <= 2;  //125 / 60 = 2
    16'b01111101_00111101 : OUT <= 2;  //125 / 61 = 2
    16'b01111101_00111110 : OUT <= 2;  //125 / 62 = 2
    16'b01111101_00111111 : OUT <= 1;  //125 / 63 = 1
    16'b01111101_01000000 : OUT <= 1;  //125 / 64 = 1
    16'b01111101_01000001 : OUT <= 1;  //125 / 65 = 1
    16'b01111101_01000010 : OUT <= 1;  //125 / 66 = 1
    16'b01111101_01000011 : OUT <= 1;  //125 / 67 = 1
    16'b01111101_01000100 : OUT <= 1;  //125 / 68 = 1
    16'b01111101_01000101 : OUT <= 1;  //125 / 69 = 1
    16'b01111101_01000110 : OUT <= 1;  //125 / 70 = 1
    16'b01111101_01000111 : OUT <= 1;  //125 / 71 = 1
    16'b01111101_01001000 : OUT <= 1;  //125 / 72 = 1
    16'b01111101_01001001 : OUT <= 1;  //125 / 73 = 1
    16'b01111101_01001010 : OUT <= 1;  //125 / 74 = 1
    16'b01111101_01001011 : OUT <= 1;  //125 / 75 = 1
    16'b01111101_01001100 : OUT <= 1;  //125 / 76 = 1
    16'b01111101_01001101 : OUT <= 1;  //125 / 77 = 1
    16'b01111101_01001110 : OUT <= 1;  //125 / 78 = 1
    16'b01111101_01001111 : OUT <= 1;  //125 / 79 = 1
    16'b01111101_01010000 : OUT <= 1;  //125 / 80 = 1
    16'b01111101_01010001 : OUT <= 1;  //125 / 81 = 1
    16'b01111101_01010010 : OUT <= 1;  //125 / 82 = 1
    16'b01111101_01010011 : OUT <= 1;  //125 / 83 = 1
    16'b01111101_01010100 : OUT <= 1;  //125 / 84 = 1
    16'b01111101_01010101 : OUT <= 1;  //125 / 85 = 1
    16'b01111101_01010110 : OUT <= 1;  //125 / 86 = 1
    16'b01111101_01010111 : OUT <= 1;  //125 / 87 = 1
    16'b01111101_01011000 : OUT <= 1;  //125 / 88 = 1
    16'b01111101_01011001 : OUT <= 1;  //125 / 89 = 1
    16'b01111101_01011010 : OUT <= 1;  //125 / 90 = 1
    16'b01111101_01011011 : OUT <= 1;  //125 / 91 = 1
    16'b01111101_01011100 : OUT <= 1;  //125 / 92 = 1
    16'b01111101_01011101 : OUT <= 1;  //125 / 93 = 1
    16'b01111101_01011110 : OUT <= 1;  //125 / 94 = 1
    16'b01111101_01011111 : OUT <= 1;  //125 / 95 = 1
    16'b01111101_01100000 : OUT <= 1;  //125 / 96 = 1
    16'b01111101_01100001 : OUT <= 1;  //125 / 97 = 1
    16'b01111101_01100010 : OUT <= 1;  //125 / 98 = 1
    16'b01111101_01100011 : OUT <= 1;  //125 / 99 = 1
    16'b01111101_01100100 : OUT <= 1;  //125 / 100 = 1
    16'b01111101_01100101 : OUT <= 1;  //125 / 101 = 1
    16'b01111101_01100110 : OUT <= 1;  //125 / 102 = 1
    16'b01111101_01100111 : OUT <= 1;  //125 / 103 = 1
    16'b01111101_01101000 : OUT <= 1;  //125 / 104 = 1
    16'b01111101_01101001 : OUT <= 1;  //125 / 105 = 1
    16'b01111101_01101010 : OUT <= 1;  //125 / 106 = 1
    16'b01111101_01101011 : OUT <= 1;  //125 / 107 = 1
    16'b01111101_01101100 : OUT <= 1;  //125 / 108 = 1
    16'b01111101_01101101 : OUT <= 1;  //125 / 109 = 1
    16'b01111101_01101110 : OUT <= 1;  //125 / 110 = 1
    16'b01111101_01101111 : OUT <= 1;  //125 / 111 = 1
    16'b01111101_01110000 : OUT <= 1;  //125 / 112 = 1
    16'b01111101_01110001 : OUT <= 1;  //125 / 113 = 1
    16'b01111101_01110010 : OUT <= 1;  //125 / 114 = 1
    16'b01111101_01110011 : OUT <= 1;  //125 / 115 = 1
    16'b01111101_01110100 : OUT <= 1;  //125 / 116 = 1
    16'b01111101_01110101 : OUT <= 1;  //125 / 117 = 1
    16'b01111101_01110110 : OUT <= 1;  //125 / 118 = 1
    16'b01111101_01110111 : OUT <= 1;  //125 / 119 = 1
    16'b01111101_01111000 : OUT <= 1;  //125 / 120 = 1
    16'b01111101_01111001 : OUT <= 1;  //125 / 121 = 1
    16'b01111101_01111010 : OUT <= 1;  //125 / 122 = 1
    16'b01111101_01111011 : OUT <= 1;  //125 / 123 = 1
    16'b01111101_01111100 : OUT <= 1;  //125 / 124 = 1
    16'b01111101_01111101 : OUT <= 1;  //125 / 125 = 1
    16'b01111101_01111110 : OUT <= 0;  //125 / 126 = 0
    16'b01111101_01111111 : OUT <= 0;  //125 / 127 = 0
    16'b01111101_10000000 : OUT <= 0;  //125 / 128 = 0
    16'b01111101_10000001 : OUT <= 0;  //125 / 129 = 0
    16'b01111101_10000010 : OUT <= 0;  //125 / 130 = 0
    16'b01111101_10000011 : OUT <= 0;  //125 / 131 = 0
    16'b01111101_10000100 : OUT <= 0;  //125 / 132 = 0
    16'b01111101_10000101 : OUT <= 0;  //125 / 133 = 0
    16'b01111101_10000110 : OUT <= 0;  //125 / 134 = 0
    16'b01111101_10000111 : OUT <= 0;  //125 / 135 = 0
    16'b01111101_10001000 : OUT <= 0;  //125 / 136 = 0
    16'b01111101_10001001 : OUT <= 0;  //125 / 137 = 0
    16'b01111101_10001010 : OUT <= 0;  //125 / 138 = 0
    16'b01111101_10001011 : OUT <= 0;  //125 / 139 = 0
    16'b01111101_10001100 : OUT <= 0;  //125 / 140 = 0
    16'b01111101_10001101 : OUT <= 0;  //125 / 141 = 0
    16'b01111101_10001110 : OUT <= 0;  //125 / 142 = 0
    16'b01111101_10001111 : OUT <= 0;  //125 / 143 = 0
    16'b01111101_10010000 : OUT <= 0;  //125 / 144 = 0
    16'b01111101_10010001 : OUT <= 0;  //125 / 145 = 0
    16'b01111101_10010010 : OUT <= 0;  //125 / 146 = 0
    16'b01111101_10010011 : OUT <= 0;  //125 / 147 = 0
    16'b01111101_10010100 : OUT <= 0;  //125 / 148 = 0
    16'b01111101_10010101 : OUT <= 0;  //125 / 149 = 0
    16'b01111101_10010110 : OUT <= 0;  //125 / 150 = 0
    16'b01111101_10010111 : OUT <= 0;  //125 / 151 = 0
    16'b01111101_10011000 : OUT <= 0;  //125 / 152 = 0
    16'b01111101_10011001 : OUT <= 0;  //125 / 153 = 0
    16'b01111101_10011010 : OUT <= 0;  //125 / 154 = 0
    16'b01111101_10011011 : OUT <= 0;  //125 / 155 = 0
    16'b01111101_10011100 : OUT <= 0;  //125 / 156 = 0
    16'b01111101_10011101 : OUT <= 0;  //125 / 157 = 0
    16'b01111101_10011110 : OUT <= 0;  //125 / 158 = 0
    16'b01111101_10011111 : OUT <= 0;  //125 / 159 = 0
    16'b01111101_10100000 : OUT <= 0;  //125 / 160 = 0
    16'b01111101_10100001 : OUT <= 0;  //125 / 161 = 0
    16'b01111101_10100010 : OUT <= 0;  //125 / 162 = 0
    16'b01111101_10100011 : OUT <= 0;  //125 / 163 = 0
    16'b01111101_10100100 : OUT <= 0;  //125 / 164 = 0
    16'b01111101_10100101 : OUT <= 0;  //125 / 165 = 0
    16'b01111101_10100110 : OUT <= 0;  //125 / 166 = 0
    16'b01111101_10100111 : OUT <= 0;  //125 / 167 = 0
    16'b01111101_10101000 : OUT <= 0;  //125 / 168 = 0
    16'b01111101_10101001 : OUT <= 0;  //125 / 169 = 0
    16'b01111101_10101010 : OUT <= 0;  //125 / 170 = 0
    16'b01111101_10101011 : OUT <= 0;  //125 / 171 = 0
    16'b01111101_10101100 : OUT <= 0;  //125 / 172 = 0
    16'b01111101_10101101 : OUT <= 0;  //125 / 173 = 0
    16'b01111101_10101110 : OUT <= 0;  //125 / 174 = 0
    16'b01111101_10101111 : OUT <= 0;  //125 / 175 = 0
    16'b01111101_10110000 : OUT <= 0;  //125 / 176 = 0
    16'b01111101_10110001 : OUT <= 0;  //125 / 177 = 0
    16'b01111101_10110010 : OUT <= 0;  //125 / 178 = 0
    16'b01111101_10110011 : OUT <= 0;  //125 / 179 = 0
    16'b01111101_10110100 : OUT <= 0;  //125 / 180 = 0
    16'b01111101_10110101 : OUT <= 0;  //125 / 181 = 0
    16'b01111101_10110110 : OUT <= 0;  //125 / 182 = 0
    16'b01111101_10110111 : OUT <= 0;  //125 / 183 = 0
    16'b01111101_10111000 : OUT <= 0;  //125 / 184 = 0
    16'b01111101_10111001 : OUT <= 0;  //125 / 185 = 0
    16'b01111101_10111010 : OUT <= 0;  //125 / 186 = 0
    16'b01111101_10111011 : OUT <= 0;  //125 / 187 = 0
    16'b01111101_10111100 : OUT <= 0;  //125 / 188 = 0
    16'b01111101_10111101 : OUT <= 0;  //125 / 189 = 0
    16'b01111101_10111110 : OUT <= 0;  //125 / 190 = 0
    16'b01111101_10111111 : OUT <= 0;  //125 / 191 = 0
    16'b01111101_11000000 : OUT <= 0;  //125 / 192 = 0
    16'b01111101_11000001 : OUT <= 0;  //125 / 193 = 0
    16'b01111101_11000010 : OUT <= 0;  //125 / 194 = 0
    16'b01111101_11000011 : OUT <= 0;  //125 / 195 = 0
    16'b01111101_11000100 : OUT <= 0;  //125 / 196 = 0
    16'b01111101_11000101 : OUT <= 0;  //125 / 197 = 0
    16'b01111101_11000110 : OUT <= 0;  //125 / 198 = 0
    16'b01111101_11000111 : OUT <= 0;  //125 / 199 = 0
    16'b01111101_11001000 : OUT <= 0;  //125 / 200 = 0
    16'b01111101_11001001 : OUT <= 0;  //125 / 201 = 0
    16'b01111101_11001010 : OUT <= 0;  //125 / 202 = 0
    16'b01111101_11001011 : OUT <= 0;  //125 / 203 = 0
    16'b01111101_11001100 : OUT <= 0;  //125 / 204 = 0
    16'b01111101_11001101 : OUT <= 0;  //125 / 205 = 0
    16'b01111101_11001110 : OUT <= 0;  //125 / 206 = 0
    16'b01111101_11001111 : OUT <= 0;  //125 / 207 = 0
    16'b01111101_11010000 : OUT <= 0;  //125 / 208 = 0
    16'b01111101_11010001 : OUT <= 0;  //125 / 209 = 0
    16'b01111101_11010010 : OUT <= 0;  //125 / 210 = 0
    16'b01111101_11010011 : OUT <= 0;  //125 / 211 = 0
    16'b01111101_11010100 : OUT <= 0;  //125 / 212 = 0
    16'b01111101_11010101 : OUT <= 0;  //125 / 213 = 0
    16'b01111101_11010110 : OUT <= 0;  //125 / 214 = 0
    16'b01111101_11010111 : OUT <= 0;  //125 / 215 = 0
    16'b01111101_11011000 : OUT <= 0;  //125 / 216 = 0
    16'b01111101_11011001 : OUT <= 0;  //125 / 217 = 0
    16'b01111101_11011010 : OUT <= 0;  //125 / 218 = 0
    16'b01111101_11011011 : OUT <= 0;  //125 / 219 = 0
    16'b01111101_11011100 : OUT <= 0;  //125 / 220 = 0
    16'b01111101_11011101 : OUT <= 0;  //125 / 221 = 0
    16'b01111101_11011110 : OUT <= 0;  //125 / 222 = 0
    16'b01111101_11011111 : OUT <= 0;  //125 / 223 = 0
    16'b01111101_11100000 : OUT <= 0;  //125 / 224 = 0
    16'b01111101_11100001 : OUT <= 0;  //125 / 225 = 0
    16'b01111101_11100010 : OUT <= 0;  //125 / 226 = 0
    16'b01111101_11100011 : OUT <= 0;  //125 / 227 = 0
    16'b01111101_11100100 : OUT <= 0;  //125 / 228 = 0
    16'b01111101_11100101 : OUT <= 0;  //125 / 229 = 0
    16'b01111101_11100110 : OUT <= 0;  //125 / 230 = 0
    16'b01111101_11100111 : OUT <= 0;  //125 / 231 = 0
    16'b01111101_11101000 : OUT <= 0;  //125 / 232 = 0
    16'b01111101_11101001 : OUT <= 0;  //125 / 233 = 0
    16'b01111101_11101010 : OUT <= 0;  //125 / 234 = 0
    16'b01111101_11101011 : OUT <= 0;  //125 / 235 = 0
    16'b01111101_11101100 : OUT <= 0;  //125 / 236 = 0
    16'b01111101_11101101 : OUT <= 0;  //125 / 237 = 0
    16'b01111101_11101110 : OUT <= 0;  //125 / 238 = 0
    16'b01111101_11101111 : OUT <= 0;  //125 / 239 = 0
    16'b01111101_11110000 : OUT <= 0;  //125 / 240 = 0
    16'b01111101_11110001 : OUT <= 0;  //125 / 241 = 0
    16'b01111101_11110010 : OUT <= 0;  //125 / 242 = 0
    16'b01111101_11110011 : OUT <= 0;  //125 / 243 = 0
    16'b01111101_11110100 : OUT <= 0;  //125 / 244 = 0
    16'b01111101_11110101 : OUT <= 0;  //125 / 245 = 0
    16'b01111101_11110110 : OUT <= 0;  //125 / 246 = 0
    16'b01111101_11110111 : OUT <= 0;  //125 / 247 = 0
    16'b01111101_11111000 : OUT <= 0;  //125 / 248 = 0
    16'b01111101_11111001 : OUT <= 0;  //125 / 249 = 0
    16'b01111101_11111010 : OUT <= 0;  //125 / 250 = 0
    16'b01111101_11111011 : OUT <= 0;  //125 / 251 = 0
    16'b01111101_11111100 : OUT <= 0;  //125 / 252 = 0
    16'b01111101_11111101 : OUT <= 0;  //125 / 253 = 0
    16'b01111101_11111110 : OUT <= 0;  //125 / 254 = 0
    16'b01111101_11111111 : OUT <= 0;  //125 / 255 = 0
    16'b01111110_00000000 : OUT <= 0;  //126 / 0 = 0
    16'b01111110_00000001 : OUT <= 126;  //126 / 1 = 126
    16'b01111110_00000010 : OUT <= 63;  //126 / 2 = 63
    16'b01111110_00000011 : OUT <= 42;  //126 / 3 = 42
    16'b01111110_00000100 : OUT <= 31;  //126 / 4 = 31
    16'b01111110_00000101 : OUT <= 25;  //126 / 5 = 25
    16'b01111110_00000110 : OUT <= 21;  //126 / 6 = 21
    16'b01111110_00000111 : OUT <= 18;  //126 / 7 = 18
    16'b01111110_00001000 : OUT <= 15;  //126 / 8 = 15
    16'b01111110_00001001 : OUT <= 14;  //126 / 9 = 14
    16'b01111110_00001010 : OUT <= 12;  //126 / 10 = 12
    16'b01111110_00001011 : OUT <= 11;  //126 / 11 = 11
    16'b01111110_00001100 : OUT <= 10;  //126 / 12 = 10
    16'b01111110_00001101 : OUT <= 9;  //126 / 13 = 9
    16'b01111110_00001110 : OUT <= 9;  //126 / 14 = 9
    16'b01111110_00001111 : OUT <= 8;  //126 / 15 = 8
    16'b01111110_00010000 : OUT <= 7;  //126 / 16 = 7
    16'b01111110_00010001 : OUT <= 7;  //126 / 17 = 7
    16'b01111110_00010010 : OUT <= 7;  //126 / 18 = 7
    16'b01111110_00010011 : OUT <= 6;  //126 / 19 = 6
    16'b01111110_00010100 : OUT <= 6;  //126 / 20 = 6
    16'b01111110_00010101 : OUT <= 6;  //126 / 21 = 6
    16'b01111110_00010110 : OUT <= 5;  //126 / 22 = 5
    16'b01111110_00010111 : OUT <= 5;  //126 / 23 = 5
    16'b01111110_00011000 : OUT <= 5;  //126 / 24 = 5
    16'b01111110_00011001 : OUT <= 5;  //126 / 25 = 5
    16'b01111110_00011010 : OUT <= 4;  //126 / 26 = 4
    16'b01111110_00011011 : OUT <= 4;  //126 / 27 = 4
    16'b01111110_00011100 : OUT <= 4;  //126 / 28 = 4
    16'b01111110_00011101 : OUT <= 4;  //126 / 29 = 4
    16'b01111110_00011110 : OUT <= 4;  //126 / 30 = 4
    16'b01111110_00011111 : OUT <= 4;  //126 / 31 = 4
    16'b01111110_00100000 : OUT <= 3;  //126 / 32 = 3
    16'b01111110_00100001 : OUT <= 3;  //126 / 33 = 3
    16'b01111110_00100010 : OUT <= 3;  //126 / 34 = 3
    16'b01111110_00100011 : OUT <= 3;  //126 / 35 = 3
    16'b01111110_00100100 : OUT <= 3;  //126 / 36 = 3
    16'b01111110_00100101 : OUT <= 3;  //126 / 37 = 3
    16'b01111110_00100110 : OUT <= 3;  //126 / 38 = 3
    16'b01111110_00100111 : OUT <= 3;  //126 / 39 = 3
    16'b01111110_00101000 : OUT <= 3;  //126 / 40 = 3
    16'b01111110_00101001 : OUT <= 3;  //126 / 41 = 3
    16'b01111110_00101010 : OUT <= 3;  //126 / 42 = 3
    16'b01111110_00101011 : OUT <= 2;  //126 / 43 = 2
    16'b01111110_00101100 : OUT <= 2;  //126 / 44 = 2
    16'b01111110_00101101 : OUT <= 2;  //126 / 45 = 2
    16'b01111110_00101110 : OUT <= 2;  //126 / 46 = 2
    16'b01111110_00101111 : OUT <= 2;  //126 / 47 = 2
    16'b01111110_00110000 : OUT <= 2;  //126 / 48 = 2
    16'b01111110_00110001 : OUT <= 2;  //126 / 49 = 2
    16'b01111110_00110010 : OUT <= 2;  //126 / 50 = 2
    16'b01111110_00110011 : OUT <= 2;  //126 / 51 = 2
    16'b01111110_00110100 : OUT <= 2;  //126 / 52 = 2
    16'b01111110_00110101 : OUT <= 2;  //126 / 53 = 2
    16'b01111110_00110110 : OUT <= 2;  //126 / 54 = 2
    16'b01111110_00110111 : OUT <= 2;  //126 / 55 = 2
    16'b01111110_00111000 : OUT <= 2;  //126 / 56 = 2
    16'b01111110_00111001 : OUT <= 2;  //126 / 57 = 2
    16'b01111110_00111010 : OUT <= 2;  //126 / 58 = 2
    16'b01111110_00111011 : OUT <= 2;  //126 / 59 = 2
    16'b01111110_00111100 : OUT <= 2;  //126 / 60 = 2
    16'b01111110_00111101 : OUT <= 2;  //126 / 61 = 2
    16'b01111110_00111110 : OUT <= 2;  //126 / 62 = 2
    16'b01111110_00111111 : OUT <= 2;  //126 / 63 = 2
    16'b01111110_01000000 : OUT <= 1;  //126 / 64 = 1
    16'b01111110_01000001 : OUT <= 1;  //126 / 65 = 1
    16'b01111110_01000010 : OUT <= 1;  //126 / 66 = 1
    16'b01111110_01000011 : OUT <= 1;  //126 / 67 = 1
    16'b01111110_01000100 : OUT <= 1;  //126 / 68 = 1
    16'b01111110_01000101 : OUT <= 1;  //126 / 69 = 1
    16'b01111110_01000110 : OUT <= 1;  //126 / 70 = 1
    16'b01111110_01000111 : OUT <= 1;  //126 / 71 = 1
    16'b01111110_01001000 : OUT <= 1;  //126 / 72 = 1
    16'b01111110_01001001 : OUT <= 1;  //126 / 73 = 1
    16'b01111110_01001010 : OUT <= 1;  //126 / 74 = 1
    16'b01111110_01001011 : OUT <= 1;  //126 / 75 = 1
    16'b01111110_01001100 : OUT <= 1;  //126 / 76 = 1
    16'b01111110_01001101 : OUT <= 1;  //126 / 77 = 1
    16'b01111110_01001110 : OUT <= 1;  //126 / 78 = 1
    16'b01111110_01001111 : OUT <= 1;  //126 / 79 = 1
    16'b01111110_01010000 : OUT <= 1;  //126 / 80 = 1
    16'b01111110_01010001 : OUT <= 1;  //126 / 81 = 1
    16'b01111110_01010010 : OUT <= 1;  //126 / 82 = 1
    16'b01111110_01010011 : OUT <= 1;  //126 / 83 = 1
    16'b01111110_01010100 : OUT <= 1;  //126 / 84 = 1
    16'b01111110_01010101 : OUT <= 1;  //126 / 85 = 1
    16'b01111110_01010110 : OUT <= 1;  //126 / 86 = 1
    16'b01111110_01010111 : OUT <= 1;  //126 / 87 = 1
    16'b01111110_01011000 : OUT <= 1;  //126 / 88 = 1
    16'b01111110_01011001 : OUT <= 1;  //126 / 89 = 1
    16'b01111110_01011010 : OUT <= 1;  //126 / 90 = 1
    16'b01111110_01011011 : OUT <= 1;  //126 / 91 = 1
    16'b01111110_01011100 : OUT <= 1;  //126 / 92 = 1
    16'b01111110_01011101 : OUT <= 1;  //126 / 93 = 1
    16'b01111110_01011110 : OUT <= 1;  //126 / 94 = 1
    16'b01111110_01011111 : OUT <= 1;  //126 / 95 = 1
    16'b01111110_01100000 : OUT <= 1;  //126 / 96 = 1
    16'b01111110_01100001 : OUT <= 1;  //126 / 97 = 1
    16'b01111110_01100010 : OUT <= 1;  //126 / 98 = 1
    16'b01111110_01100011 : OUT <= 1;  //126 / 99 = 1
    16'b01111110_01100100 : OUT <= 1;  //126 / 100 = 1
    16'b01111110_01100101 : OUT <= 1;  //126 / 101 = 1
    16'b01111110_01100110 : OUT <= 1;  //126 / 102 = 1
    16'b01111110_01100111 : OUT <= 1;  //126 / 103 = 1
    16'b01111110_01101000 : OUT <= 1;  //126 / 104 = 1
    16'b01111110_01101001 : OUT <= 1;  //126 / 105 = 1
    16'b01111110_01101010 : OUT <= 1;  //126 / 106 = 1
    16'b01111110_01101011 : OUT <= 1;  //126 / 107 = 1
    16'b01111110_01101100 : OUT <= 1;  //126 / 108 = 1
    16'b01111110_01101101 : OUT <= 1;  //126 / 109 = 1
    16'b01111110_01101110 : OUT <= 1;  //126 / 110 = 1
    16'b01111110_01101111 : OUT <= 1;  //126 / 111 = 1
    16'b01111110_01110000 : OUT <= 1;  //126 / 112 = 1
    16'b01111110_01110001 : OUT <= 1;  //126 / 113 = 1
    16'b01111110_01110010 : OUT <= 1;  //126 / 114 = 1
    16'b01111110_01110011 : OUT <= 1;  //126 / 115 = 1
    16'b01111110_01110100 : OUT <= 1;  //126 / 116 = 1
    16'b01111110_01110101 : OUT <= 1;  //126 / 117 = 1
    16'b01111110_01110110 : OUT <= 1;  //126 / 118 = 1
    16'b01111110_01110111 : OUT <= 1;  //126 / 119 = 1
    16'b01111110_01111000 : OUT <= 1;  //126 / 120 = 1
    16'b01111110_01111001 : OUT <= 1;  //126 / 121 = 1
    16'b01111110_01111010 : OUT <= 1;  //126 / 122 = 1
    16'b01111110_01111011 : OUT <= 1;  //126 / 123 = 1
    16'b01111110_01111100 : OUT <= 1;  //126 / 124 = 1
    16'b01111110_01111101 : OUT <= 1;  //126 / 125 = 1
    16'b01111110_01111110 : OUT <= 1;  //126 / 126 = 1
    16'b01111110_01111111 : OUT <= 0;  //126 / 127 = 0
    16'b01111110_10000000 : OUT <= 0;  //126 / 128 = 0
    16'b01111110_10000001 : OUT <= 0;  //126 / 129 = 0
    16'b01111110_10000010 : OUT <= 0;  //126 / 130 = 0
    16'b01111110_10000011 : OUT <= 0;  //126 / 131 = 0
    16'b01111110_10000100 : OUT <= 0;  //126 / 132 = 0
    16'b01111110_10000101 : OUT <= 0;  //126 / 133 = 0
    16'b01111110_10000110 : OUT <= 0;  //126 / 134 = 0
    16'b01111110_10000111 : OUT <= 0;  //126 / 135 = 0
    16'b01111110_10001000 : OUT <= 0;  //126 / 136 = 0
    16'b01111110_10001001 : OUT <= 0;  //126 / 137 = 0
    16'b01111110_10001010 : OUT <= 0;  //126 / 138 = 0
    16'b01111110_10001011 : OUT <= 0;  //126 / 139 = 0
    16'b01111110_10001100 : OUT <= 0;  //126 / 140 = 0
    16'b01111110_10001101 : OUT <= 0;  //126 / 141 = 0
    16'b01111110_10001110 : OUT <= 0;  //126 / 142 = 0
    16'b01111110_10001111 : OUT <= 0;  //126 / 143 = 0
    16'b01111110_10010000 : OUT <= 0;  //126 / 144 = 0
    16'b01111110_10010001 : OUT <= 0;  //126 / 145 = 0
    16'b01111110_10010010 : OUT <= 0;  //126 / 146 = 0
    16'b01111110_10010011 : OUT <= 0;  //126 / 147 = 0
    16'b01111110_10010100 : OUT <= 0;  //126 / 148 = 0
    16'b01111110_10010101 : OUT <= 0;  //126 / 149 = 0
    16'b01111110_10010110 : OUT <= 0;  //126 / 150 = 0
    16'b01111110_10010111 : OUT <= 0;  //126 / 151 = 0
    16'b01111110_10011000 : OUT <= 0;  //126 / 152 = 0
    16'b01111110_10011001 : OUT <= 0;  //126 / 153 = 0
    16'b01111110_10011010 : OUT <= 0;  //126 / 154 = 0
    16'b01111110_10011011 : OUT <= 0;  //126 / 155 = 0
    16'b01111110_10011100 : OUT <= 0;  //126 / 156 = 0
    16'b01111110_10011101 : OUT <= 0;  //126 / 157 = 0
    16'b01111110_10011110 : OUT <= 0;  //126 / 158 = 0
    16'b01111110_10011111 : OUT <= 0;  //126 / 159 = 0
    16'b01111110_10100000 : OUT <= 0;  //126 / 160 = 0
    16'b01111110_10100001 : OUT <= 0;  //126 / 161 = 0
    16'b01111110_10100010 : OUT <= 0;  //126 / 162 = 0
    16'b01111110_10100011 : OUT <= 0;  //126 / 163 = 0
    16'b01111110_10100100 : OUT <= 0;  //126 / 164 = 0
    16'b01111110_10100101 : OUT <= 0;  //126 / 165 = 0
    16'b01111110_10100110 : OUT <= 0;  //126 / 166 = 0
    16'b01111110_10100111 : OUT <= 0;  //126 / 167 = 0
    16'b01111110_10101000 : OUT <= 0;  //126 / 168 = 0
    16'b01111110_10101001 : OUT <= 0;  //126 / 169 = 0
    16'b01111110_10101010 : OUT <= 0;  //126 / 170 = 0
    16'b01111110_10101011 : OUT <= 0;  //126 / 171 = 0
    16'b01111110_10101100 : OUT <= 0;  //126 / 172 = 0
    16'b01111110_10101101 : OUT <= 0;  //126 / 173 = 0
    16'b01111110_10101110 : OUT <= 0;  //126 / 174 = 0
    16'b01111110_10101111 : OUT <= 0;  //126 / 175 = 0
    16'b01111110_10110000 : OUT <= 0;  //126 / 176 = 0
    16'b01111110_10110001 : OUT <= 0;  //126 / 177 = 0
    16'b01111110_10110010 : OUT <= 0;  //126 / 178 = 0
    16'b01111110_10110011 : OUT <= 0;  //126 / 179 = 0
    16'b01111110_10110100 : OUT <= 0;  //126 / 180 = 0
    16'b01111110_10110101 : OUT <= 0;  //126 / 181 = 0
    16'b01111110_10110110 : OUT <= 0;  //126 / 182 = 0
    16'b01111110_10110111 : OUT <= 0;  //126 / 183 = 0
    16'b01111110_10111000 : OUT <= 0;  //126 / 184 = 0
    16'b01111110_10111001 : OUT <= 0;  //126 / 185 = 0
    16'b01111110_10111010 : OUT <= 0;  //126 / 186 = 0
    16'b01111110_10111011 : OUT <= 0;  //126 / 187 = 0
    16'b01111110_10111100 : OUT <= 0;  //126 / 188 = 0
    16'b01111110_10111101 : OUT <= 0;  //126 / 189 = 0
    16'b01111110_10111110 : OUT <= 0;  //126 / 190 = 0
    16'b01111110_10111111 : OUT <= 0;  //126 / 191 = 0
    16'b01111110_11000000 : OUT <= 0;  //126 / 192 = 0
    16'b01111110_11000001 : OUT <= 0;  //126 / 193 = 0
    16'b01111110_11000010 : OUT <= 0;  //126 / 194 = 0
    16'b01111110_11000011 : OUT <= 0;  //126 / 195 = 0
    16'b01111110_11000100 : OUT <= 0;  //126 / 196 = 0
    16'b01111110_11000101 : OUT <= 0;  //126 / 197 = 0
    16'b01111110_11000110 : OUT <= 0;  //126 / 198 = 0
    16'b01111110_11000111 : OUT <= 0;  //126 / 199 = 0
    16'b01111110_11001000 : OUT <= 0;  //126 / 200 = 0
    16'b01111110_11001001 : OUT <= 0;  //126 / 201 = 0
    16'b01111110_11001010 : OUT <= 0;  //126 / 202 = 0
    16'b01111110_11001011 : OUT <= 0;  //126 / 203 = 0
    16'b01111110_11001100 : OUT <= 0;  //126 / 204 = 0
    16'b01111110_11001101 : OUT <= 0;  //126 / 205 = 0
    16'b01111110_11001110 : OUT <= 0;  //126 / 206 = 0
    16'b01111110_11001111 : OUT <= 0;  //126 / 207 = 0
    16'b01111110_11010000 : OUT <= 0;  //126 / 208 = 0
    16'b01111110_11010001 : OUT <= 0;  //126 / 209 = 0
    16'b01111110_11010010 : OUT <= 0;  //126 / 210 = 0
    16'b01111110_11010011 : OUT <= 0;  //126 / 211 = 0
    16'b01111110_11010100 : OUT <= 0;  //126 / 212 = 0
    16'b01111110_11010101 : OUT <= 0;  //126 / 213 = 0
    16'b01111110_11010110 : OUT <= 0;  //126 / 214 = 0
    16'b01111110_11010111 : OUT <= 0;  //126 / 215 = 0
    16'b01111110_11011000 : OUT <= 0;  //126 / 216 = 0
    16'b01111110_11011001 : OUT <= 0;  //126 / 217 = 0
    16'b01111110_11011010 : OUT <= 0;  //126 / 218 = 0
    16'b01111110_11011011 : OUT <= 0;  //126 / 219 = 0
    16'b01111110_11011100 : OUT <= 0;  //126 / 220 = 0
    16'b01111110_11011101 : OUT <= 0;  //126 / 221 = 0
    16'b01111110_11011110 : OUT <= 0;  //126 / 222 = 0
    16'b01111110_11011111 : OUT <= 0;  //126 / 223 = 0
    16'b01111110_11100000 : OUT <= 0;  //126 / 224 = 0
    16'b01111110_11100001 : OUT <= 0;  //126 / 225 = 0
    16'b01111110_11100010 : OUT <= 0;  //126 / 226 = 0
    16'b01111110_11100011 : OUT <= 0;  //126 / 227 = 0
    16'b01111110_11100100 : OUT <= 0;  //126 / 228 = 0
    16'b01111110_11100101 : OUT <= 0;  //126 / 229 = 0
    16'b01111110_11100110 : OUT <= 0;  //126 / 230 = 0
    16'b01111110_11100111 : OUT <= 0;  //126 / 231 = 0
    16'b01111110_11101000 : OUT <= 0;  //126 / 232 = 0
    16'b01111110_11101001 : OUT <= 0;  //126 / 233 = 0
    16'b01111110_11101010 : OUT <= 0;  //126 / 234 = 0
    16'b01111110_11101011 : OUT <= 0;  //126 / 235 = 0
    16'b01111110_11101100 : OUT <= 0;  //126 / 236 = 0
    16'b01111110_11101101 : OUT <= 0;  //126 / 237 = 0
    16'b01111110_11101110 : OUT <= 0;  //126 / 238 = 0
    16'b01111110_11101111 : OUT <= 0;  //126 / 239 = 0
    16'b01111110_11110000 : OUT <= 0;  //126 / 240 = 0
    16'b01111110_11110001 : OUT <= 0;  //126 / 241 = 0
    16'b01111110_11110010 : OUT <= 0;  //126 / 242 = 0
    16'b01111110_11110011 : OUT <= 0;  //126 / 243 = 0
    16'b01111110_11110100 : OUT <= 0;  //126 / 244 = 0
    16'b01111110_11110101 : OUT <= 0;  //126 / 245 = 0
    16'b01111110_11110110 : OUT <= 0;  //126 / 246 = 0
    16'b01111110_11110111 : OUT <= 0;  //126 / 247 = 0
    16'b01111110_11111000 : OUT <= 0;  //126 / 248 = 0
    16'b01111110_11111001 : OUT <= 0;  //126 / 249 = 0
    16'b01111110_11111010 : OUT <= 0;  //126 / 250 = 0
    16'b01111110_11111011 : OUT <= 0;  //126 / 251 = 0
    16'b01111110_11111100 : OUT <= 0;  //126 / 252 = 0
    16'b01111110_11111101 : OUT <= 0;  //126 / 253 = 0
    16'b01111110_11111110 : OUT <= 0;  //126 / 254 = 0
    16'b01111110_11111111 : OUT <= 0;  //126 / 255 = 0
    16'b01111111_00000000 : OUT <= 0;  //127 / 0 = 0
    16'b01111111_00000001 : OUT <= 127;  //127 / 1 = 127
    16'b01111111_00000010 : OUT <= 63;  //127 / 2 = 63
    16'b01111111_00000011 : OUT <= 42;  //127 / 3 = 42
    16'b01111111_00000100 : OUT <= 31;  //127 / 4 = 31
    16'b01111111_00000101 : OUT <= 25;  //127 / 5 = 25
    16'b01111111_00000110 : OUT <= 21;  //127 / 6 = 21
    16'b01111111_00000111 : OUT <= 18;  //127 / 7 = 18
    16'b01111111_00001000 : OUT <= 15;  //127 / 8 = 15
    16'b01111111_00001001 : OUT <= 14;  //127 / 9 = 14
    16'b01111111_00001010 : OUT <= 12;  //127 / 10 = 12
    16'b01111111_00001011 : OUT <= 11;  //127 / 11 = 11
    16'b01111111_00001100 : OUT <= 10;  //127 / 12 = 10
    16'b01111111_00001101 : OUT <= 9;  //127 / 13 = 9
    16'b01111111_00001110 : OUT <= 9;  //127 / 14 = 9
    16'b01111111_00001111 : OUT <= 8;  //127 / 15 = 8
    16'b01111111_00010000 : OUT <= 7;  //127 / 16 = 7
    16'b01111111_00010001 : OUT <= 7;  //127 / 17 = 7
    16'b01111111_00010010 : OUT <= 7;  //127 / 18 = 7
    16'b01111111_00010011 : OUT <= 6;  //127 / 19 = 6
    16'b01111111_00010100 : OUT <= 6;  //127 / 20 = 6
    16'b01111111_00010101 : OUT <= 6;  //127 / 21 = 6
    16'b01111111_00010110 : OUT <= 5;  //127 / 22 = 5
    16'b01111111_00010111 : OUT <= 5;  //127 / 23 = 5
    16'b01111111_00011000 : OUT <= 5;  //127 / 24 = 5
    16'b01111111_00011001 : OUT <= 5;  //127 / 25 = 5
    16'b01111111_00011010 : OUT <= 4;  //127 / 26 = 4
    16'b01111111_00011011 : OUT <= 4;  //127 / 27 = 4
    16'b01111111_00011100 : OUT <= 4;  //127 / 28 = 4
    16'b01111111_00011101 : OUT <= 4;  //127 / 29 = 4
    16'b01111111_00011110 : OUT <= 4;  //127 / 30 = 4
    16'b01111111_00011111 : OUT <= 4;  //127 / 31 = 4
    16'b01111111_00100000 : OUT <= 3;  //127 / 32 = 3
    16'b01111111_00100001 : OUT <= 3;  //127 / 33 = 3
    16'b01111111_00100010 : OUT <= 3;  //127 / 34 = 3
    16'b01111111_00100011 : OUT <= 3;  //127 / 35 = 3
    16'b01111111_00100100 : OUT <= 3;  //127 / 36 = 3
    16'b01111111_00100101 : OUT <= 3;  //127 / 37 = 3
    16'b01111111_00100110 : OUT <= 3;  //127 / 38 = 3
    16'b01111111_00100111 : OUT <= 3;  //127 / 39 = 3
    16'b01111111_00101000 : OUT <= 3;  //127 / 40 = 3
    16'b01111111_00101001 : OUT <= 3;  //127 / 41 = 3
    16'b01111111_00101010 : OUT <= 3;  //127 / 42 = 3
    16'b01111111_00101011 : OUT <= 2;  //127 / 43 = 2
    16'b01111111_00101100 : OUT <= 2;  //127 / 44 = 2
    16'b01111111_00101101 : OUT <= 2;  //127 / 45 = 2
    16'b01111111_00101110 : OUT <= 2;  //127 / 46 = 2
    16'b01111111_00101111 : OUT <= 2;  //127 / 47 = 2
    16'b01111111_00110000 : OUT <= 2;  //127 / 48 = 2
    16'b01111111_00110001 : OUT <= 2;  //127 / 49 = 2
    16'b01111111_00110010 : OUT <= 2;  //127 / 50 = 2
    16'b01111111_00110011 : OUT <= 2;  //127 / 51 = 2
    16'b01111111_00110100 : OUT <= 2;  //127 / 52 = 2
    16'b01111111_00110101 : OUT <= 2;  //127 / 53 = 2
    16'b01111111_00110110 : OUT <= 2;  //127 / 54 = 2
    16'b01111111_00110111 : OUT <= 2;  //127 / 55 = 2
    16'b01111111_00111000 : OUT <= 2;  //127 / 56 = 2
    16'b01111111_00111001 : OUT <= 2;  //127 / 57 = 2
    16'b01111111_00111010 : OUT <= 2;  //127 / 58 = 2
    16'b01111111_00111011 : OUT <= 2;  //127 / 59 = 2
    16'b01111111_00111100 : OUT <= 2;  //127 / 60 = 2
    16'b01111111_00111101 : OUT <= 2;  //127 / 61 = 2
    16'b01111111_00111110 : OUT <= 2;  //127 / 62 = 2
    16'b01111111_00111111 : OUT <= 2;  //127 / 63 = 2
    16'b01111111_01000000 : OUT <= 1;  //127 / 64 = 1
    16'b01111111_01000001 : OUT <= 1;  //127 / 65 = 1
    16'b01111111_01000010 : OUT <= 1;  //127 / 66 = 1
    16'b01111111_01000011 : OUT <= 1;  //127 / 67 = 1
    16'b01111111_01000100 : OUT <= 1;  //127 / 68 = 1
    16'b01111111_01000101 : OUT <= 1;  //127 / 69 = 1
    16'b01111111_01000110 : OUT <= 1;  //127 / 70 = 1
    16'b01111111_01000111 : OUT <= 1;  //127 / 71 = 1
    16'b01111111_01001000 : OUT <= 1;  //127 / 72 = 1
    16'b01111111_01001001 : OUT <= 1;  //127 / 73 = 1
    16'b01111111_01001010 : OUT <= 1;  //127 / 74 = 1
    16'b01111111_01001011 : OUT <= 1;  //127 / 75 = 1
    16'b01111111_01001100 : OUT <= 1;  //127 / 76 = 1
    16'b01111111_01001101 : OUT <= 1;  //127 / 77 = 1
    16'b01111111_01001110 : OUT <= 1;  //127 / 78 = 1
    16'b01111111_01001111 : OUT <= 1;  //127 / 79 = 1
    16'b01111111_01010000 : OUT <= 1;  //127 / 80 = 1
    16'b01111111_01010001 : OUT <= 1;  //127 / 81 = 1
    16'b01111111_01010010 : OUT <= 1;  //127 / 82 = 1
    16'b01111111_01010011 : OUT <= 1;  //127 / 83 = 1
    16'b01111111_01010100 : OUT <= 1;  //127 / 84 = 1
    16'b01111111_01010101 : OUT <= 1;  //127 / 85 = 1
    16'b01111111_01010110 : OUT <= 1;  //127 / 86 = 1
    16'b01111111_01010111 : OUT <= 1;  //127 / 87 = 1
    16'b01111111_01011000 : OUT <= 1;  //127 / 88 = 1
    16'b01111111_01011001 : OUT <= 1;  //127 / 89 = 1
    16'b01111111_01011010 : OUT <= 1;  //127 / 90 = 1
    16'b01111111_01011011 : OUT <= 1;  //127 / 91 = 1
    16'b01111111_01011100 : OUT <= 1;  //127 / 92 = 1
    16'b01111111_01011101 : OUT <= 1;  //127 / 93 = 1
    16'b01111111_01011110 : OUT <= 1;  //127 / 94 = 1
    16'b01111111_01011111 : OUT <= 1;  //127 / 95 = 1
    16'b01111111_01100000 : OUT <= 1;  //127 / 96 = 1
    16'b01111111_01100001 : OUT <= 1;  //127 / 97 = 1
    16'b01111111_01100010 : OUT <= 1;  //127 / 98 = 1
    16'b01111111_01100011 : OUT <= 1;  //127 / 99 = 1
    16'b01111111_01100100 : OUT <= 1;  //127 / 100 = 1
    16'b01111111_01100101 : OUT <= 1;  //127 / 101 = 1
    16'b01111111_01100110 : OUT <= 1;  //127 / 102 = 1
    16'b01111111_01100111 : OUT <= 1;  //127 / 103 = 1
    16'b01111111_01101000 : OUT <= 1;  //127 / 104 = 1
    16'b01111111_01101001 : OUT <= 1;  //127 / 105 = 1
    16'b01111111_01101010 : OUT <= 1;  //127 / 106 = 1
    16'b01111111_01101011 : OUT <= 1;  //127 / 107 = 1
    16'b01111111_01101100 : OUT <= 1;  //127 / 108 = 1
    16'b01111111_01101101 : OUT <= 1;  //127 / 109 = 1
    16'b01111111_01101110 : OUT <= 1;  //127 / 110 = 1
    16'b01111111_01101111 : OUT <= 1;  //127 / 111 = 1
    16'b01111111_01110000 : OUT <= 1;  //127 / 112 = 1
    16'b01111111_01110001 : OUT <= 1;  //127 / 113 = 1
    16'b01111111_01110010 : OUT <= 1;  //127 / 114 = 1
    16'b01111111_01110011 : OUT <= 1;  //127 / 115 = 1
    16'b01111111_01110100 : OUT <= 1;  //127 / 116 = 1
    16'b01111111_01110101 : OUT <= 1;  //127 / 117 = 1
    16'b01111111_01110110 : OUT <= 1;  //127 / 118 = 1
    16'b01111111_01110111 : OUT <= 1;  //127 / 119 = 1
    16'b01111111_01111000 : OUT <= 1;  //127 / 120 = 1
    16'b01111111_01111001 : OUT <= 1;  //127 / 121 = 1
    16'b01111111_01111010 : OUT <= 1;  //127 / 122 = 1
    16'b01111111_01111011 : OUT <= 1;  //127 / 123 = 1
    16'b01111111_01111100 : OUT <= 1;  //127 / 124 = 1
    16'b01111111_01111101 : OUT <= 1;  //127 / 125 = 1
    16'b01111111_01111110 : OUT <= 1;  //127 / 126 = 1
    16'b01111111_01111111 : OUT <= 1;  //127 / 127 = 1
    16'b01111111_10000000 : OUT <= 0;  //127 / 128 = 0
    16'b01111111_10000001 : OUT <= 0;  //127 / 129 = 0
    16'b01111111_10000010 : OUT <= 0;  //127 / 130 = 0
    16'b01111111_10000011 : OUT <= 0;  //127 / 131 = 0
    16'b01111111_10000100 : OUT <= 0;  //127 / 132 = 0
    16'b01111111_10000101 : OUT <= 0;  //127 / 133 = 0
    16'b01111111_10000110 : OUT <= 0;  //127 / 134 = 0
    16'b01111111_10000111 : OUT <= 0;  //127 / 135 = 0
    16'b01111111_10001000 : OUT <= 0;  //127 / 136 = 0
    16'b01111111_10001001 : OUT <= 0;  //127 / 137 = 0
    16'b01111111_10001010 : OUT <= 0;  //127 / 138 = 0
    16'b01111111_10001011 : OUT <= 0;  //127 / 139 = 0
    16'b01111111_10001100 : OUT <= 0;  //127 / 140 = 0
    16'b01111111_10001101 : OUT <= 0;  //127 / 141 = 0
    16'b01111111_10001110 : OUT <= 0;  //127 / 142 = 0
    16'b01111111_10001111 : OUT <= 0;  //127 / 143 = 0
    16'b01111111_10010000 : OUT <= 0;  //127 / 144 = 0
    16'b01111111_10010001 : OUT <= 0;  //127 / 145 = 0
    16'b01111111_10010010 : OUT <= 0;  //127 / 146 = 0
    16'b01111111_10010011 : OUT <= 0;  //127 / 147 = 0
    16'b01111111_10010100 : OUT <= 0;  //127 / 148 = 0
    16'b01111111_10010101 : OUT <= 0;  //127 / 149 = 0
    16'b01111111_10010110 : OUT <= 0;  //127 / 150 = 0
    16'b01111111_10010111 : OUT <= 0;  //127 / 151 = 0
    16'b01111111_10011000 : OUT <= 0;  //127 / 152 = 0
    16'b01111111_10011001 : OUT <= 0;  //127 / 153 = 0
    16'b01111111_10011010 : OUT <= 0;  //127 / 154 = 0
    16'b01111111_10011011 : OUT <= 0;  //127 / 155 = 0
    16'b01111111_10011100 : OUT <= 0;  //127 / 156 = 0
    16'b01111111_10011101 : OUT <= 0;  //127 / 157 = 0
    16'b01111111_10011110 : OUT <= 0;  //127 / 158 = 0
    16'b01111111_10011111 : OUT <= 0;  //127 / 159 = 0
    16'b01111111_10100000 : OUT <= 0;  //127 / 160 = 0
    16'b01111111_10100001 : OUT <= 0;  //127 / 161 = 0
    16'b01111111_10100010 : OUT <= 0;  //127 / 162 = 0
    16'b01111111_10100011 : OUT <= 0;  //127 / 163 = 0
    16'b01111111_10100100 : OUT <= 0;  //127 / 164 = 0
    16'b01111111_10100101 : OUT <= 0;  //127 / 165 = 0
    16'b01111111_10100110 : OUT <= 0;  //127 / 166 = 0
    16'b01111111_10100111 : OUT <= 0;  //127 / 167 = 0
    16'b01111111_10101000 : OUT <= 0;  //127 / 168 = 0
    16'b01111111_10101001 : OUT <= 0;  //127 / 169 = 0
    16'b01111111_10101010 : OUT <= 0;  //127 / 170 = 0
    16'b01111111_10101011 : OUT <= 0;  //127 / 171 = 0
    16'b01111111_10101100 : OUT <= 0;  //127 / 172 = 0
    16'b01111111_10101101 : OUT <= 0;  //127 / 173 = 0
    16'b01111111_10101110 : OUT <= 0;  //127 / 174 = 0
    16'b01111111_10101111 : OUT <= 0;  //127 / 175 = 0
    16'b01111111_10110000 : OUT <= 0;  //127 / 176 = 0
    16'b01111111_10110001 : OUT <= 0;  //127 / 177 = 0
    16'b01111111_10110010 : OUT <= 0;  //127 / 178 = 0
    16'b01111111_10110011 : OUT <= 0;  //127 / 179 = 0
    16'b01111111_10110100 : OUT <= 0;  //127 / 180 = 0
    16'b01111111_10110101 : OUT <= 0;  //127 / 181 = 0
    16'b01111111_10110110 : OUT <= 0;  //127 / 182 = 0
    16'b01111111_10110111 : OUT <= 0;  //127 / 183 = 0
    16'b01111111_10111000 : OUT <= 0;  //127 / 184 = 0
    16'b01111111_10111001 : OUT <= 0;  //127 / 185 = 0
    16'b01111111_10111010 : OUT <= 0;  //127 / 186 = 0
    16'b01111111_10111011 : OUT <= 0;  //127 / 187 = 0
    16'b01111111_10111100 : OUT <= 0;  //127 / 188 = 0
    16'b01111111_10111101 : OUT <= 0;  //127 / 189 = 0
    16'b01111111_10111110 : OUT <= 0;  //127 / 190 = 0
    16'b01111111_10111111 : OUT <= 0;  //127 / 191 = 0
    16'b01111111_11000000 : OUT <= 0;  //127 / 192 = 0
    16'b01111111_11000001 : OUT <= 0;  //127 / 193 = 0
    16'b01111111_11000010 : OUT <= 0;  //127 / 194 = 0
    16'b01111111_11000011 : OUT <= 0;  //127 / 195 = 0
    16'b01111111_11000100 : OUT <= 0;  //127 / 196 = 0
    16'b01111111_11000101 : OUT <= 0;  //127 / 197 = 0
    16'b01111111_11000110 : OUT <= 0;  //127 / 198 = 0
    16'b01111111_11000111 : OUT <= 0;  //127 / 199 = 0
    16'b01111111_11001000 : OUT <= 0;  //127 / 200 = 0
    16'b01111111_11001001 : OUT <= 0;  //127 / 201 = 0
    16'b01111111_11001010 : OUT <= 0;  //127 / 202 = 0
    16'b01111111_11001011 : OUT <= 0;  //127 / 203 = 0
    16'b01111111_11001100 : OUT <= 0;  //127 / 204 = 0
    16'b01111111_11001101 : OUT <= 0;  //127 / 205 = 0
    16'b01111111_11001110 : OUT <= 0;  //127 / 206 = 0
    16'b01111111_11001111 : OUT <= 0;  //127 / 207 = 0
    16'b01111111_11010000 : OUT <= 0;  //127 / 208 = 0
    16'b01111111_11010001 : OUT <= 0;  //127 / 209 = 0
    16'b01111111_11010010 : OUT <= 0;  //127 / 210 = 0
    16'b01111111_11010011 : OUT <= 0;  //127 / 211 = 0
    16'b01111111_11010100 : OUT <= 0;  //127 / 212 = 0
    16'b01111111_11010101 : OUT <= 0;  //127 / 213 = 0
    16'b01111111_11010110 : OUT <= 0;  //127 / 214 = 0
    16'b01111111_11010111 : OUT <= 0;  //127 / 215 = 0
    16'b01111111_11011000 : OUT <= 0;  //127 / 216 = 0
    16'b01111111_11011001 : OUT <= 0;  //127 / 217 = 0
    16'b01111111_11011010 : OUT <= 0;  //127 / 218 = 0
    16'b01111111_11011011 : OUT <= 0;  //127 / 219 = 0
    16'b01111111_11011100 : OUT <= 0;  //127 / 220 = 0
    16'b01111111_11011101 : OUT <= 0;  //127 / 221 = 0
    16'b01111111_11011110 : OUT <= 0;  //127 / 222 = 0
    16'b01111111_11011111 : OUT <= 0;  //127 / 223 = 0
    16'b01111111_11100000 : OUT <= 0;  //127 / 224 = 0
    16'b01111111_11100001 : OUT <= 0;  //127 / 225 = 0
    16'b01111111_11100010 : OUT <= 0;  //127 / 226 = 0
    16'b01111111_11100011 : OUT <= 0;  //127 / 227 = 0
    16'b01111111_11100100 : OUT <= 0;  //127 / 228 = 0
    16'b01111111_11100101 : OUT <= 0;  //127 / 229 = 0
    16'b01111111_11100110 : OUT <= 0;  //127 / 230 = 0
    16'b01111111_11100111 : OUT <= 0;  //127 / 231 = 0
    16'b01111111_11101000 : OUT <= 0;  //127 / 232 = 0
    16'b01111111_11101001 : OUT <= 0;  //127 / 233 = 0
    16'b01111111_11101010 : OUT <= 0;  //127 / 234 = 0
    16'b01111111_11101011 : OUT <= 0;  //127 / 235 = 0
    16'b01111111_11101100 : OUT <= 0;  //127 / 236 = 0
    16'b01111111_11101101 : OUT <= 0;  //127 / 237 = 0
    16'b01111111_11101110 : OUT <= 0;  //127 / 238 = 0
    16'b01111111_11101111 : OUT <= 0;  //127 / 239 = 0
    16'b01111111_11110000 : OUT <= 0;  //127 / 240 = 0
    16'b01111111_11110001 : OUT <= 0;  //127 / 241 = 0
    16'b01111111_11110010 : OUT <= 0;  //127 / 242 = 0
    16'b01111111_11110011 : OUT <= 0;  //127 / 243 = 0
    16'b01111111_11110100 : OUT <= 0;  //127 / 244 = 0
    16'b01111111_11110101 : OUT <= 0;  //127 / 245 = 0
    16'b01111111_11110110 : OUT <= 0;  //127 / 246 = 0
    16'b01111111_11110111 : OUT <= 0;  //127 / 247 = 0
    16'b01111111_11111000 : OUT <= 0;  //127 / 248 = 0
    16'b01111111_11111001 : OUT <= 0;  //127 / 249 = 0
    16'b01111111_11111010 : OUT <= 0;  //127 / 250 = 0
    16'b01111111_11111011 : OUT <= 0;  //127 / 251 = 0
    16'b01111111_11111100 : OUT <= 0;  //127 / 252 = 0
    16'b01111111_11111101 : OUT <= 0;  //127 / 253 = 0
    16'b01111111_11111110 : OUT <= 0;  //127 / 254 = 0
    16'b01111111_11111111 : OUT <= 0;  //127 / 255 = 0
    16'b10000000_00000000 : OUT <= 0;  //128 / 0 = 0
    16'b10000000_00000001 : OUT <= 128;  //128 / 1 = 128
    16'b10000000_00000010 : OUT <= 64;  //128 / 2 = 64
    16'b10000000_00000011 : OUT <= 42;  //128 / 3 = 42
    16'b10000000_00000100 : OUT <= 32;  //128 / 4 = 32
    16'b10000000_00000101 : OUT <= 25;  //128 / 5 = 25
    16'b10000000_00000110 : OUT <= 21;  //128 / 6 = 21
    16'b10000000_00000111 : OUT <= 18;  //128 / 7 = 18
    16'b10000000_00001000 : OUT <= 16;  //128 / 8 = 16
    16'b10000000_00001001 : OUT <= 14;  //128 / 9 = 14
    16'b10000000_00001010 : OUT <= 12;  //128 / 10 = 12
    16'b10000000_00001011 : OUT <= 11;  //128 / 11 = 11
    16'b10000000_00001100 : OUT <= 10;  //128 / 12 = 10
    16'b10000000_00001101 : OUT <= 9;  //128 / 13 = 9
    16'b10000000_00001110 : OUT <= 9;  //128 / 14 = 9
    16'b10000000_00001111 : OUT <= 8;  //128 / 15 = 8
    16'b10000000_00010000 : OUT <= 8;  //128 / 16 = 8
    16'b10000000_00010001 : OUT <= 7;  //128 / 17 = 7
    16'b10000000_00010010 : OUT <= 7;  //128 / 18 = 7
    16'b10000000_00010011 : OUT <= 6;  //128 / 19 = 6
    16'b10000000_00010100 : OUT <= 6;  //128 / 20 = 6
    16'b10000000_00010101 : OUT <= 6;  //128 / 21 = 6
    16'b10000000_00010110 : OUT <= 5;  //128 / 22 = 5
    16'b10000000_00010111 : OUT <= 5;  //128 / 23 = 5
    16'b10000000_00011000 : OUT <= 5;  //128 / 24 = 5
    16'b10000000_00011001 : OUT <= 5;  //128 / 25 = 5
    16'b10000000_00011010 : OUT <= 4;  //128 / 26 = 4
    16'b10000000_00011011 : OUT <= 4;  //128 / 27 = 4
    16'b10000000_00011100 : OUT <= 4;  //128 / 28 = 4
    16'b10000000_00011101 : OUT <= 4;  //128 / 29 = 4
    16'b10000000_00011110 : OUT <= 4;  //128 / 30 = 4
    16'b10000000_00011111 : OUT <= 4;  //128 / 31 = 4
    16'b10000000_00100000 : OUT <= 4;  //128 / 32 = 4
    16'b10000000_00100001 : OUT <= 3;  //128 / 33 = 3
    16'b10000000_00100010 : OUT <= 3;  //128 / 34 = 3
    16'b10000000_00100011 : OUT <= 3;  //128 / 35 = 3
    16'b10000000_00100100 : OUT <= 3;  //128 / 36 = 3
    16'b10000000_00100101 : OUT <= 3;  //128 / 37 = 3
    16'b10000000_00100110 : OUT <= 3;  //128 / 38 = 3
    16'b10000000_00100111 : OUT <= 3;  //128 / 39 = 3
    16'b10000000_00101000 : OUT <= 3;  //128 / 40 = 3
    16'b10000000_00101001 : OUT <= 3;  //128 / 41 = 3
    16'b10000000_00101010 : OUT <= 3;  //128 / 42 = 3
    16'b10000000_00101011 : OUT <= 2;  //128 / 43 = 2
    16'b10000000_00101100 : OUT <= 2;  //128 / 44 = 2
    16'b10000000_00101101 : OUT <= 2;  //128 / 45 = 2
    16'b10000000_00101110 : OUT <= 2;  //128 / 46 = 2
    16'b10000000_00101111 : OUT <= 2;  //128 / 47 = 2
    16'b10000000_00110000 : OUT <= 2;  //128 / 48 = 2
    16'b10000000_00110001 : OUT <= 2;  //128 / 49 = 2
    16'b10000000_00110010 : OUT <= 2;  //128 / 50 = 2
    16'b10000000_00110011 : OUT <= 2;  //128 / 51 = 2
    16'b10000000_00110100 : OUT <= 2;  //128 / 52 = 2
    16'b10000000_00110101 : OUT <= 2;  //128 / 53 = 2
    16'b10000000_00110110 : OUT <= 2;  //128 / 54 = 2
    16'b10000000_00110111 : OUT <= 2;  //128 / 55 = 2
    16'b10000000_00111000 : OUT <= 2;  //128 / 56 = 2
    16'b10000000_00111001 : OUT <= 2;  //128 / 57 = 2
    16'b10000000_00111010 : OUT <= 2;  //128 / 58 = 2
    16'b10000000_00111011 : OUT <= 2;  //128 / 59 = 2
    16'b10000000_00111100 : OUT <= 2;  //128 / 60 = 2
    16'b10000000_00111101 : OUT <= 2;  //128 / 61 = 2
    16'b10000000_00111110 : OUT <= 2;  //128 / 62 = 2
    16'b10000000_00111111 : OUT <= 2;  //128 / 63 = 2
    16'b10000000_01000000 : OUT <= 2;  //128 / 64 = 2
    16'b10000000_01000001 : OUT <= 1;  //128 / 65 = 1
    16'b10000000_01000010 : OUT <= 1;  //128 / 66 = 1
    16'b10000000_01000011 : OUT <= 1;  //128 / 67 = 1
    16'b10000000_01000100 : OUT <= 1;  //128 / 68 = 1
    16'b10000000_01000101 : OUT <= 1;  //128 / 69 = 1
    16'b10000000_01000110 : OUT <= 1;  //128 / 70 = 1
    16'b10000000_01000111 : OUT <= 1;  //128 / 71 = 1
    16'b10000000_01001000 : OUT <= 1;  //128 / 72 = 1
    16'b10000000_01001001 : OUT <= 1;  //128 / 73 = 1
    16'b10000000_01001010 : OUT <= 1;  //128 / 74 = 1
    16'b10000000_01001011 : OUT <= 1;  //128 / 75 = 1
    16'b10000000_01001100 : OUT <= 1;  //128 / 76 = 1
    16'b10000000_01001101 : OUT <= 1;  //128 / 77 = 1
    16'b10000000_01001110 : OUT <= 1;  //128 / 78 = 1
    16'b10000000_01001111 : OUT <= 1;  //128 / 79 = 1
    16'b10000000_01010000 : OUT <= 1;  //128 / 80 = 1
    16'b10000000_01010001 : OUT <= 1;  //128 / 81 = 1
    16'b10000000_01010010 : OUT <= 1;  //128 / 82 = 1
    16'b10000000_01010011 : OUT <= 1;  //128 / 83 = 1
    16'b10000000_01010100 : OUT <= 1;  //128 / 84 = 1
    16'b10000000_01010101 : OUT <= 1;  //128 / 85 = 1
    16'b10000000_01010110 : OUT <= 1;  //128 / 86 = 1
    16'b10000000_01010111 : OUT <= 1;  //128 / 87 = 1
    16'b10000000_01011000 : OUT <= 1;  //128 / 88 = 1
    16'b10000000_01011001 : OUT <= 1;  //128 / 89 = 1
    16'b10000000_01011010 : OUT <= 1;  //128 / 90 = 1
    16'b10000000_01011011 : OUT <= 1;  //128 / 91 = 1
    16'b10000000_01011100 : OUT <= 1;  //128 / 92 = 1
    16'b10000000_01011101 : OUT <= 1;  //128 / 93 = 1
    16'b10000000_01011110 : OUT <= 1;  //128 / 94 = 1
    16'b10000000_01011111 : OUT <= 1;  //128 / 95 = 1
    16'b10000000_01100000 : OUT <= 1;  //128 / 96 = 1
    16'b10000000_01100001 : OUT <= 1;  //128 / 97 = 1
    16'b10000000_01100010 : OUT <= 1;  //128 / 98 = 1
    16'b10000000_01100011 : OUT <= 1;  //128 / 99 = 1
    16'b10000000_01100100 : OUT <= 1;  //128 / 100 = 1
    16'b10000000_01100101 : OUT <= 1;  //128 / 101 = 1
    16'b10000000_01100110 : OUT <= 1;  //128 / 102 = 1
    16'b10000000_01100111 : OUT <= 1;  //128 / 103 = 1
    16'b10000000_01101000 : OUT <= 1;  //128 / 104 = 1
    16'b10000000_01101001 : OUT <= 1;  //128 / 105 = 1
    16'b10000000_01101010 : OUT <= 1;  //128 / 106 = 1
    16'b10000000_01101011 : OUT <= 1;  //128 / 107 = 1
    16'b10000000_01101100 : OUT <= 1;  //128 / 108 = 1
    16'b10000000_01101101 : OUT <= 1;  //128 / 109 = 1
    16'b10000000_01101110 : OUT <= 1;  //128 / 110 = 1
    16'b10000000_01101111 : OUT <= 1;  //128 / 111 = 1
    16'b10000000_01110000 : OUT <= 1;  //128 / 112 = 1
    16'b10000000_01110001 : OUT <= 1;  //128 / 113 = 1
    16'b10000000_01110010 : OUT <= 1;  //128 / 114 = 1
    16'b10000000_01110011 : OUT <= 1;  //128 / 115 = 1
    16'b10000000_01110100 : OUT <= 1;  //128 / 116 = 1
    16'b10000000_01110101 : OUT <= 1;  //128 / 117 = 1
    16'b10000000_01110110 : OUT <= 1;  //128 / 118 = 1
    16'b10000000_01110111 : OUT <= 1;  //128 / 119 = 1
    16'b10000000_01111000 : OUT <= 1;  //128 / 120 = 1
    16'b10000000_01111001 : OUT <= 1;  //128 / 121 = 1
    16'b10000000_01111010 : OUT <= 1;  //128 / 122 = 1
    16'b10000000_01111011 : OUT <= 1;  //128 / 123 = 1
    16'b10000000_01111100 : OUT <= 1;  //128 / 124 = 1
    16'b10000000_01111101 : OUT <= 1;  //128 / 125 = 1
    16'b10000000_01111110 : OUT <= 1;  //128 / 126 = 1
    16'b10000000_01111111 : OUT <= 1;  //128 / 127 = 1
    16'b10000000_10000000 : OUT <= 1;  //128 / 128 = 1
    16'b10000000_10000001 : OUT <= 0;  //128 / 129 = 0
    16'b10000000_10000010 : OUT <= 0;  //128 / 130 = 0
    16'b10000000_10000011 : OUT <= 0;  //128 / 131 = 0
    16'b10000000_10000100 : OUT <= 0;  //128 / 132 = 0
    16'b10000000_10000101 : OUT <= 0;  //128 / 133 = 0
    16'b10000000_10000110 : OUT <= 0;  //128 / 134 = 0
    16'b10000000_10000111 : OUT <= 0;  //128 / 135 = 0
    16'b10000000_10001000 : OUT <= 0;  //128 / 136 = 0
    16'b10000000_10001001 : OUT <= 0;  //128 / 137 = 0
    16'b10000000_10001010 : OUT <= 0;  //128 / 138 = 0
    16'b10000000_10001011 : OUT <= 0;  //128 / 139 = 0
    16'b10000000_10001100 : OUT <= 0;  //128 / 140 = 0
    16'b10000000_10001101 : OUT <= 0;  //128 / 141 = 0
    16'b10000000_10001110 : OUT <= 0;  //128 / 142 = 0
    16'b10000000_10001111 : OUT <= 0;  //128 / 143 = 0
    16'b10000000_10010000 : OUT <= 0;  //128 / 144 = 0
    16'b10000000_10010001 : OUT <= 0;  //128 / 145 = 0
    16'b10000000_10010010 : OUT <= 0;  //128 / 146 = 0
    16'b10000000_10010011 : OUT <= 0;  //128 / 147 = 0
    16'b10000000_10010100 : OUT <= 0;  //128 / 148 = 0
    16'b10000000_10010101 : OUT <= 0;  //128 / 149 = 0
    16'b10000000_10010110 : OUT <= 0;  //128 / 150 = 0
    16'b10000000_10010111 : OUT <= 0;  //128 / 151 = 0
    16'b10000000_10011000 : OUT <= 0;  //128 / 152 = 0
    16'b10000000_10011001 : OUT <= 0;  //128 / 153 = 0
    16'b10000000_10011010 : OUT <= 0;  //128 / 154 = 0
    16'b10000000_10011011 : OUT <= 0;  //128 / 155 = 0
    16'b10000000_10011100 : OUT <= 0;  //128 / 156 = 0
    16'b10000000_10011101 : OUT <= 0;  //128 / 157 = 0
    16'b10000000_10011110 : OUT <= 0;  //128 / 158 = 0
    16'b10000000_10011111 : OUT <= 0;  //128 / 159 = 0
    16'b10000000_10100000 : OUT <= 0;  //128 / 160 = 0
    16'b10000000_10100001 : OUT <= 0;  //128 / 161 = 0
    16'b10000000_10100010 : OUT <= 0;  //128 / 162 = 0
    16'b10000000_10100011 : OUT <= 0;  //128 / 163 = 0
    16'b10000000_10100100 : OUT <= 0;  //128 / 164 = 0
    16'b10000000_10100101 : OUT <= 0;  //128 / 165 = 0
    16'b10000000_10100110 : OUT <= 0;  //128 / 166 = 0
    16'b10000000_10100111 : OUT <= 0;  //128 / 167 = 0
    16'b10000000_10101000 : OUT <= 0;  //128 / 168 = 0
    16'b10000000_10101001 : OUT <= 0;  //128 / 169 = 0
    16'b10000000_10101010 : OUT <= 0;  //128 / 170 = 0
    16'b10000000_10101011 : OUT <= 0;  //128 / 171 = 0
    16'b10000000_10101100 : OUT <= 0;  //128 / 172 = 0
    16'b10000000_10101101 : OUT <= 0;  //128 / 173 = 0
    16'b10000000_10101110 : OUT <= 0;  //128 / 174 = 0
    16'b10000000_10101111 : OUT <= 0;  //128 / 175 = 0
    16'b10000000_10110000 : OUT <= 0;  //128 / 176 = 0
    16'b10000000_10110001 : OUT <= 0;  //128 / 177 = 0
    16'b10000000_10110010 : OUT <= 0;  //128 / 178 = 0
    16'b10000000_10110011 : OUT <= 0;  //128 / 179 = 0
    16'b10000000_10110100 : OUT <= 0;  //128 / 180 = 0
    16'b10000000_10110101 : OUT <= 0;  //128 / 181 = 0
    16'b10000000_10110110 : OUT <= 0;  //128 / 182 = 0
    16'b10000000_10110111 : OUT <= 0;  //128 / 183 = 0
    16'b10000000_10111000 : OUT <= 0;  //128 / 184 = 0
    16'b10000000_10111001 : OUT <= 0;  //128 / 185 = 0
    16'b10000000_10111010 : OUT <= 0;  //128 / 186 = 0
    16'b10000000_10111011 : OUT <= 0;  //128 / 187 = 0
    16'b10000000_10111100 : OUT <= 0;  //128 / 188 = 0
    16'b10000000_10111101 : OUT <= 0;  //128 / 189 = 0
    16'b10000000_10111110 : OUT <= 0;  //128 / 190 = 0
    16'b10000000_10111111 : OUT <= 0;  //128 / 191 = 0
    16'b10000000_11000000 : OUT <= 0;  //128 / 192 = 0
    16'b10000000_11000001 : OUT <= 0;  //128 / 193 = 0
    16'b10000000_11000010 : OUT <= 0;  //128 / 194 = 0
    16'b10000000_11000011 : OUT <= 0;  //128 / 195 = 0
    16'b10000000_11000100 : OUT <= 0;  //128 / 196 = 0
    16'b10000000_11000101 : OUT <= 0;  //128 / 197 = 0
    16'b10000000_11000110 : OUT <= 0;  //128 / 198 = 0
    16'b10000000_11000111 : OUT <= 0;  //128 / 199 = 0
    16'b10000000_11001000 : OUT <= 0;  //128 / 200 = 0
    16'b10000000_11001001 : OUT <= 0;  //128 / 201 = 0
    16'b10000000_11001010 : OUT <= 0;  //128 / 202 = 0
    16'b10000000_11001011 : OUT <= 0;  //128 / 203 = 0
    16'b10000000_11001100 : OUT <= 0;  //128 / 204 = 0
    16'b10000000_11001101 : OUT <= 0;  //128 / 205 = 0
    16'b10000000_11001110 : OUT <= 0;  //128 / 206 = 0
    16'b10000000_11001111 : OUT <= 0;  //128 / 207 = 0
    16'b10000000_11010000 : OUT <= 0;  //128 / 208 = 0
    16'b10000000_11010001 : OUT <= 0;  //128 / 209 = 0
    16'b10000000_11010010 : OUT <= 0;  //128 / 210 = 0
    16'b10000000_11010011 : OUT <= 0;  //128 / 211 = 0
    16'b10000000_11010100 : OUT <= 0;  //128 / 212 = 0
    16'b10000000_11010101 : OUT <= 0;  //128 / 213 = 0
    16'b10000000_11010110 : OUT <= 0;  //128 / 214 = 0
    16'b10000000_11010111 : OUT <= 0;  //128 / 215 = 0
    16'b10000000_11011000 : OUT <= 0;  //128 / 216 = 0
    16'b10000000_11011001 : OUT <= 0;  //128 / 217 = 0
    16'b10000000_11011010 : OUT <= 0;  //128 / 218 = 0
    16'b10000000_11011011 : OUT <= 0;  //128 / 219 = 0
    16'b10000000_11011100 : OUT <= 0;  //128 / 220 = 0
    16'b10000000_11011101 : OUT <= 0;  //128 / 221 = 0
    16'b10000000_11011110 : OUT <= 0;  //128 / 222 = 0
    16'b10000000_11011111 : OUT <= 0;  //128 / 223 = 0
    16'b10000000_11100000 : OUT <= 0;  //128 / 224 = 0
    16'b10000000_11100001 : OUT <= 0;  //128 / 225 = 0
    16'b10000000_11100010 : OUT <= 0;  //128 / 226 = 0
    16'b10000000_11100011 : OUT <= 0;  //128 / 227 = 0
    16'b10000000_11100100 : OUT <= 0;  //128 / 228 = 0
    16'b10000000_11100101 : OUT <= 0;  //128 / 229 = 0
    16'b10000000_11100110 : OUT <= 0;  //128 / 230 = 0
    16'b10000000_11100111 : OUT <= 0;  //128 / 231 = 0
    16'b10000000_11101000 : OUT <= 0;  //128 / 232 = 0
    16'b10000000_11101001 : OUT <= 0;  //128 / 233 = 0
    16'b10000000_11101010 : OUT <= 0;  //128 / 234 = 0
    16'b10000000_11101011 : OUT <= 0;  //128 / 235 = 0
    16'b10000000_11101100 : OUT <= 0;  //128 / 236 = 0
    16'b10000000_11101101 : OUT <= 0;  //128 / 237 = 0
    16'b10000000_11101110 : OUT <= 0;  //128 / 238 = 0
    16'b10000000_11101111 : OUT <= 0;  //128 / 239 = 0
    16'b10000000_11110000 : OUT <= 0;  //128 / 240 = 0
    16'b10000000_11110001 : OUT <= 0;  //128 / 241 = 0
    16'b10000000_11110010 : OUT <= 0;  //128 / 242 = 0
    16'b10000000_11110011 : OUT <= 0;  //128 / 243 = 0
    16'b10000000_11110100 : OUT <= 0;  //128 / 244 = 0
    16'b10000000_11110101 : OUT <= 0;  //128 / 245 = 0
    16'b10000000_11110110 : OUT <= 0;  //128 / 246 = 0
    16'b10000000_11110111 : OUT <= 0;  //128 / 247 = 0
    16'b10000000_11111000 : OUT <= 0;  //128 / 248 = 0
    16'b10000000_11111001 : OUT <= 0;  //128 / 249 = 0
    16'b10000000_11111010 : OUT <= 0;  //128 / 250 = 0
    16'b10000000_11111011 : OUT <= 0;  //128 / 251 = 0
    16'b10000000_11111100 : OUT <= 0;  //128 / 252 = 0
    16'b10000000_11111101 : OUT <= 0;  //128 / 253 = 0
    16'b10000000_11111110 : OUT <= 0;  //128 / 254 = 0
    16'b10000000_11111111 : OUT <= 0;  //128 / 255 = 0
    16'b10000001_00000000 : OUT <= 0;  //129 / 0 = 0
    16'b10000001_00000001 : OUT <= 129;  //129 / 1 = 129
    16'b10000001_00000010 : OUT <= 64;  //129 / 2 = 64
    16'b10000001_00000011 : OUT <= 43;  //129 / 3 = 43
    16'b10000001_00000100 : OUT <= 32;  //129 / 4 = 32
    16'b10000001_00000101 : OUT <= 25;  //129 / 5 = 25
    16'b10000001_00000110 : OUT <= 21;  //129 / 6 = 21
    16'b10000001_00000111 : OUT <= 18;  //129 / 7 = 18
    16'b10000001_00001000 : OUT <= 16;  //129 / 8 = 16
    16'b10000001_00001001 : OUT <= 14;  //129 / 9 = 14
    16'b10000001_00001010 : OUT <= 12;  //129 / 10 = 12
    16'b10000001_00001011 : OUT <= 11;  //129 / 11 = 11
    16'b10000001_00001100 : OUT <= 10;  //129 / 12 = 10
    16'b10000001_00001101 : OUT <= 9;  //129 / 13 = 9
    16'b10000001_00001110 : OUT <= 9;  //129 / 14 = 9
    16'b10000001_00001111 : OUT <= 8;  //129 / 15 = 8
    16'b10000001_00010000 : OUT <= 8;  //129 / 16 = 8
    16'b10000001_00010001 : OUT <= 7;  //129 / 17 = 7
    16'b10000001_00010010 : OUT <= 7;  //129 / 18 = 7
    16'b10000001_00010011 : OUT <= 6;  //129 / 19 = 6
    16'b10000001_00010100 : OUT <= 6;  //129 / 20 = 6
    16'b10000001_00010101 : OUT <= 6;  //129 / 21 = 6
    16'b10000001_00010110 : OUT <= 5;  //129 / 22 = 5
    16'b10000001_00010111 : OUT <= 5;  //129 / 23 = 5
    16'b10000001_00011000 : OUT <= 5;  //129 / 24 = 5
    16'b10000001_00011001 : OUT <= 5;  //129 / 25 = 5
    16'b10000001_00011010 : OUT <= 4;  //129 / 26 = 4
    16'b10000001_00011011 : OUT <= 4;  //129 / 27 = 4
    16'b10000001_00011100 : OUT <= 4;  //129 / 28 = 4
    16'b10000001_00011101 : OUT <= 4;  //129 / 29 = 4
    16'b10000001_00011110 : OUT <= 4;  //129 / 30 = 4
    16'b10000001_00011111 : OUT <= 4;  //129 / 31 = 4
    16'b10000001_00100000 : OUT <= 4;  //129 / 32 = 4
    16'b10000001_00100001 : OUT <= 3;  //129 / 33 = 3
    16'b10000001_00100010 : OUT <= 3;  //129 / 34 = 3
    16'b10000001_00100011 : OUT <= 3;  //129 / 35 = 3
    16'b10000001_00100100 : OUT <= 3;  //129 / 36 = 3
    16'b10000001_00100101 : OUT <= 3;  //129 / 37 = 3
    16'b10000001_00100110 : OUT <= 3;  //129 / 38 = 3
    16'b10000001_00100111 : OUT <= 3;  //129 / 39 = 3
    16'b10000001_00101000 : OUT <= 3;  //129 / 40 = 3
    16'b10000001_00101001 : OUT <= 3;  //129 / 41 = 3
    16'b10000001_00101010 : OUT <= 3;  //129 / 42 = 3
    16'b10000001_00101011 : OUT <= 3;  //129 / 43 = 3
    16'b10000001_00101100 : OUT <= 2;  //129 / 44 = 2
    16'b10000001_00101101 : OUT <= 2;  //129 / 45 = 2
    16'b10000001_00101110 : OUT <= 2;  //129 / 46 = 2
    16'b10000001_00101111 : OUT <= 2;  //129 / 47 = 2
    16'b10000001_00110000 : OUT <= 2;  //129 / 48 = 2
    16'b10000001_00110001 : OUT <= 2;  //129 / 49 = 2
    16'b10000001_00110010 : OUT <= 2;  //129 / 50 = 2
    16'b10000001_00110011 : OUT <= 2;  //129 / 51 = 2
    16'b10000001_00110100 : OUT <= 2;  //129 / 52 = 2
    16'b10000001_00110101 : OUT <= 2;  //129 / 53 = 2
    16'b10000001_00110110 : OUT <= 2;  //129 / 54 = 2
    16'b10000001_00110111 : OUT <= 2;  //129 / 55 = 2
    16'b10000001_00111000 : OUT <= 2;  //129 / 56 = 2
    16'b10000001_00111001 : OUT <= 2;  //129 / 57 = 2
    16'b10000001_00111010 : OUT <= 2;  //129 / 58 = 2
    16'b10000001_00111011 : OUT <= 2;  //129 / 59 = 2
    16'b10000001_00111100 : OUT <= 2;  //129 / 60 = 2
    16'b10000001_00111101 : OUT <= 2;  //129 / 61 = 2
    16'b10000001_00111110 : OUT <= 2;  //129 / 62 = 2
    16'b10000001_00111111 : OUT <= 2;  //129 / 63 = 2
    16'b10000001_01000000 : OUT <= 2;  //129 / 64 = 2
    16'b10000001_01000001 : OUT <= 1;  //129 / 65 = 1
    16'b10000001_01000010 : OUT <= 1;  //129 / 66 = 1
    16'b10000001_01000011 : OUT <= 1;  //129 / 67 = 1
    16'b10000001_01000100 : OUT <= 1;  //129 / 68 = 1
    16'b10000001_01000101 : OUT <= 1;  //129 / 69 = 1
    16'b10000001_01000110 : OUT <= 1;  //129 / 70 = 1
    16'b10000001_01000111 : OUT <= 1;  //129 / 71 = 1
    16'b10000001_01001000 : OUT <= 1;  //129 / 72 = 1
    16'b10000001_01001001 : OUT <= 1;  //129 / 73 = 1
    16'b10000001_01001010 : OUT <= 1;  //129 / 74 = 1
    16'b10000001_01001011 : OUT <= 1;  //129 / 75 = 1
    16'b10000001_01001100 : OUT <= 1;  //129 / 76 = 1
    16'b10000001_01001101 : OUT <= 1;  //129 / 77 = 1
    16'b10000001_01001110 : OUT <= 1;  //129 / 78 = 1
    16'b10000001_01001111 : OUT <= 1;  //129 / 79 = 1
    16'b10000001_01010000 : OUT <= 1;  //129 / 80 = 1
    16'b10000001_01010001 : OUT <= 1;  //129 / 81 = 1
    16'b10000001_01010010 : OUT <= 1;  //129 / 82 = 1
    16'b10000001_01010011 : OUT <= 1;  //129 / 83 = 1
    16'b10000001_01010100 : OUT <= 1;  //129 / 84 = 1
    16'b10000001_01010101 : OUT <= 1;  //129 / 85 = 1
    16'b10000001_01010110 : OUT <= 1;  //129 / 86 = 1
    16'b10000001_01010111 : OUT <= 1;  //129 / 87 = 1
    16'b10000001_01011000 : OUT <= 1;  //129 / 88 = 1
    16'b10000001_01011001 : OUT <= 1;  //129 / 89 = 1
    16'b10000001_01011010 : OUT <= 1;  //129 / 90 = 1
    16'b10000001_01011011 : OUT <= 1;  //129 / 91 = 1
    16'b10000001_01011100 : OUT <= 1;  //129 / 92 = 1
    16'b10000001_01011101 : OUT <= 1;  //129 / 93 = 1
    16'b10000001_01011110 : OUT <= 1;  //129 / 94 = 1
    16'b10000001_01011111 : OUT <= 1;  //129 / 95 = 1
    16'b10000001_01100000 : OUT <= 1;  //129 / 96 = 1
    16'b10000001_01100001 : OUT <= 1;  //129 / 97 = 1
    16'b10000001_01100010 : OUT <= 1;  //129 / 98 = 1
    16'b10000001_01100011 : OUT <= 1;  //129 / 99 = 1
    16'b10000001_01100100 : OUT <= 1;  //129 / 100 = 1
    16'b10000001_01100101 : OUT <= 1;  //129 / 101 = 1
    16'b10000001_01100110 : OUT <= 1;  //129 / 102 = 1
    16'b10000001_01100111 : OUT <= 1;  //129 / 103 = 1
    16'b10000001_01101000 : OUT <= 1;  //129 / 104 = 1
    16'b10000001_01101001 : OUT <= 1;  //129 / 105 = 1
    16'b10000001_01101010 : OUT <= 1;  //129 / 106 = 1
    16'b10000001_01101011 : OUT <= 1;  //129 / 107 = 1
    16'b10000001_01101100 : OUT <= 1;  //129 / 108 = 1
    16'b10000001_01101101 : OUT <= 1;  //129 / 109 = 1
    16'b10000001_01101110 : OUT <= 1;  //129 / 110 = 1
    16'b10000001_01101111 : OUT <= 1;  //129 / 111 = 1
    16'b10000001_01110000 : OUT <= 1;  //129 / 112 = 1
    16'b10000001_01110001 : OUT <= 1;  //129 / 113 = 1
    16'b10000001_01110010 : OUT <= 1;  //129 / 114 = 1
    16'b10000001_01110011 : OUT <= 1;  //129 / 115 = 1
    16'b10000001_01110100 : OUT <= 1;  //129 / 116 = 1
    16'b10000001_01110101 : OUT <= 1;  //129 / 117 = 1
    16'b10000001_01110110 : OUT <= 1;  //129 / 118 = 1
    16'b10000001_01110111 : OUT <= 1;  //129 / 119 = 1
    16'b10000001_01111000 : OUT <= 1;  //129 / 120 = 1
    16'b10000001_01111001 : OUT <= 1;  //129 / 121 = 1
    16'b10000001_01111010 : OUT <= 1;  //129 / 122 = 1
    16'b10000001_01111011 : OUT <= 1;  //129 / 123 = 1
    16'b10000001_01111100 : OUT <= 1;  //129 / 124 = 1
    16'b10000001_01111101 : OUT <= 1;  //129 / 125 = 1
    16'b10000001_01111110 : OUT <= 1;  //129 / 126 = 1
    16'b10000001_01111111 : OUT <= 1;  //129 / 127 = 1
    16'b10000001_10000000 : OUT <= 1;  //129 / 128 = 1
    16'b10000001_10000001 : OUT <= 1;  //129 / 129 = 1
    16'b10000001_10000010 : OUT <= 0;  //129 / 130 = 0
    16'b10000001_10000011 : OUT <= 0;  //129 / 131 = 0
    16'b10000001_10000100 : OUT <= 0;  //129 / 132 = 0
    16'b10000001_10000101 : OUT <= 0;  //129 / 133 = 0
    16'b10000001_10000110 : OUT <= 0;  //129 / 134 = 0
    16'b10000001_10000111 : OUT <= 0;  //129 / 135 = 0
    16'b10000001_10001000 : OUT <= 0;  //129 / 136 = 0
    16'b10000001_10001001 : OUT <= 0;  //129 / 137 = 0
    16'b10000001_10001010 : OUT <= 0;  //129 / 138 = 0
    16'b10000001_10001011 : OUT <= 0;  //129 / 139 = 0
    16'b10000001_10001100 : OUT <= 0;  //129 / 140 = 0
    16'b10000001_10001101 : OUT <= 0;  //129 / 141 = 0
    16'b10000001_10001110 : OUT <= 0;  //129 / 142 = 0
    16'b10000001_10001111 : OUT <= 0;  //129 / 143 = 0
    16'b10000001_10010000 : OUT <= 0;  //129 / 144 = 0
    16'b10000001_10010001 : OUT <= 0;  //129 / 145 = 0
    16'b10000001_10010010 : OUT <= 0;  //129 / 146 = 0
    16'b10000001_10010011 : OUT <= 0;  //129 / 147 = 0
    16'b10000001_10010100 : OUT <= 0;  //129 / 148 = 0
    16'b10000001_10010101 : OUT <= 0;  //129 / 149 = 0
    16'b10000001_10010110 : OUT <= 0;  //129 / 150 = 0
    16'b10000001_10010111 : OUT <= 0;  //129 / 151 = 0
    16'b10000001_10011000 : OUT <= 0;  //129 / 152 = 0
    16'b10000001_10011001 : OUT <= 0;  //129 / 153 = 0
    16'b10000001_10011010 : OUT <= 0;  //129 / 154 = 0
    16'b10000001_10011011 : OUT <= 0;  //129 / 155 = 0
    16'b10000001_10011100 : OUT <= 0;  //129 / 156 = 0
    16'b10000001_10011101 : OUT <= 0;  //129 / 157 = 0
    16'b10000001_10011110 : OUT <= 0;  //129 / 158 = 0
    16'b10000001_10011111 : OUT <= 0;  //129 / 159 = 0
    16'b10000001_10100000 : OUT <= 0;  //129 / 160 = 0
    16'b10000001_10100001 : OUT <= 0;  //129 / 161 = 0
    16'b10000001_10100010 : OUT <= 0;  //129 / 162 = 0
    16'b10000001_10100011 : OUT <= 0;  //129 / 163 = 0
    16'b10000001_10100100 : OUT <= 0;  //129 / 164 = 0
    16'b10000001_10100101 : OUT <= 0;  //129 / 165 = 0
    16'b10000001_10100110 : OUT <= 0;  //129 / 166 = 0
    16'b10000001_10100111 : OUT <= 0;  //129 / 167 = 0
    16'b10000001_10101000 : OUT <= 0;  //129 / 168 = 0
    16'b10000001_10101001 : OUT <= 0;  //129 / 169 = 0
    16'b10000001_10101010 : OUT <= 0;  //129 / 170 = 0
    16'b10000001_10101011 : OUT <= 0;  //129 / 171 = 0
    16'b10000001_10101100 : OUT <= 0;  //129 / 172 = 0
    16'b10000001_10101101 : OUT <= 0;  //129 / 173 = 0
    16'b10000001_10101110 : OUT <= 0;  //129 / 174 = 0
    16'b10000001_10101111 : OUT <= 0;  //129 / 175 = 0
    16'b10000001_10110000 : OUT <= 0;  //129 / 176 = 0
    16'b10000001_10110001 : OUT <= 0;  //129 / 177 = 0
    16'b10000001_10110010 : OUT <= 0;  //129 / 178 = 0
    16'b10000001_10110011 : OUT <= 0;  //129 / 179 = 0
    16'b10000001_10110100 : OUT <= 0;  //129 / 180 = 0
    16'b10000001_10110101 : OUT <= 0;  //129 / 181 = 0
    16'b10000001_10110110 : OUT <= 0;  //129 / 182 = 0
    16'b10000001_10110111 : OUT <= 0;  //129 / 183 = 0
    16'b10000001_10111000 : OUT <= 0;  //129 / 184 = 0
    16'b10000001_10111001 : OUT <= 0;  //129 / 185 = 0
    16'b10000001_10111010 : OUT <= 0;  //129 / 186 = 0
    16'b10000001_10111011 : OUT <= 0;  //129 / 187 = 0
    16'b10000001_10111100 : OUT <= 0;  //129 / 188 = 0
    16'b10000001_10111101 : OUT <= 0;  //129 / 189 = 0
    16'b10000001_10111110 : OUT <= 0;  //129 / 190 = 0
    16'b10000001_10111111 : OUT <= 0;  //129 / 191 = 0
    16'b10000001_11000000 : OUT <= 0;  //129 / 192 = 0
    16'b10000001_11000001 : OUT <= 0;  //129 / 193 = 0
    16'b10000001_11000010 : OUT <= 0;  //129 / 194 = 0
    16'b10000001_11000011 : OUT <= 0;  //129 / 195 = 0
    16'b10000001_11000100 : OUT <= 0;  //129 / 196 = 0
    16'b10000001_11000101 : OUT <= 0;  //129 / 197 = 0
    16'b10000001_11000110 : OUT <= 0;  //129 / 198 = 0
    16'b10000001_11000111 : OUT <= 0;  //129 / 199 = 0
    16'b10000001_11001000 : OUT <= 0;  //129 / 200 = 0
    16'b10000001_11001001 : OUT <= 0;  //129 / 201 = 0
    16'b10000001_11001010 : OUT <= 0;  //129 / 202 = 0
    16'b10000001_11001011 : OUT <= 0;  //129 / 203 = 0
    16'b10000001_11001100 : OUT <= 0;  //129 / 204 = 0
    16'b10000001_11001101 : OUT <= 0;  //129 / 205 = 0
    16'b10000001_11001110 : OUT <= 0;  //129 / 206 = 0
    16'b10000001_11001111 : OUT <= 0;  //129 / 207 = 0
    16'b10000001_11010000 : OUT <= 0;  //129 / 208 = 0
    16'b10000001_11010001 : OUT <= 0;  //129 / 209 = 0
    16'b10000001_11010010 : OUT <= 0;  //129 / 210 = 0
    16'b10000001_11010011 : OUT <= 0;  //129 / 211 = 0
    16'b10000001_11010100 : OUT <= 0;  //129 / 212 = 0
    16'b10000001_11010101 : OUT <= 0;  //129 / 213 = 0
    16'b10000001_11010110 : OUT <= 0;  //129 / 214 = 0
    16'b10000001_11010111 : OUT <= 0;  //129 / 215 = 0
    16'b10000001_11011000 : OUT <= 0;  //129 / 216 = 0
    16'b10000001_11011001 : OUT <= 0;  //129 / 217 = 0
    16'b10000001_11011010 : OUT <= 0;  //129 / 218 = 0
    16'b10000001_11011011 : OUT <= 0;  //129 / 219 = 0
    16'b10000001_11011100 : OUT <= 0;  //129 / 220 = 0
    16'b10000001_11011101 : OUT <= 0;  //129 / 221 = 0
    16'b10000001_11011110 : OUT <= 0;  //129 / 222 = 0
    16'b10000001_11011111 : OUT <= 0;  //129 / 223 = 0
    16'b10000001_11100000 : OUT <= 0;  //129 / 224 = 0
    16'b10000001_11100001 : OUT <= 0;  //129 / 225 = 0
    16'b10000001_11100010 : OUT <= 0;  //129 / 226 = 0
    16'b10000001_11100011 : OUT <= 0;  //129 / 227 = 0
    16'b10000001_11100100 : OUT <= 0;  //129 / 228 = 0
    16'b10000001_11100101 : OUT <= 0;  //129 / 229 = 0
    16'b10000001_11100110 : OUT <= 0;  //129 / 230 = 0
    16'b10000001_11100111 : OUT <= 0;  //129 / 231 = 0
    16'b10000001_11101000 : OUT <= 0;  //129 / 232 = 0
    16'b10000001_11101001 : OUT <= 0;  //129 / 233 = 0
    16'b10000001_11101010 : OUT <= 0;  //129 / 234 = 0
    16'b10000001_11101011 : OUT <= 0;  //129 / 235 = 0
    16'b10000001_11101100 : OUT <= 0;  //129 / 236 = 0
    16'b10000001_11101101 : OUT <= 0;  //129 / 237 = 0
    16'b10000001_11101110 : OUT <= 0;  //129 / 238 = 0
    16'b10000001_11101111 : OUT <= 0;  //129 / 239 = 0
    16'b10000001_11110000 : OUT <= 0;  //129 / 240 = 0
    16'b10000001_11110001 : OUT <= 0;  //129 / 241 = 0
    16'b10000001_11110010 : OUT <= 0;  //129 / 242 = 0
    16'b10000001_11110011 : OUT <= 0;  //129 / 243 = 0
    16'b10000001_11110100 : OUT <= 0;  //129 / 244 = 0
    16'b10000001_11110101 : OUT <= 0;  //129 / 245 = 0
    16'b10000001_11110110 : OUT <= 0;  //129 / 246 = 0
    16'b10000001_11110111 : OUT <= 0;  //129 / 247 = 0
    16'b10000001_11111000 : OUT <= 0;  //129 / 248 = 0
    16'b10000001_11111001 : OUT <= 0;  //129 / 249 = 0
    16'b10000001_11111010 : OUT <= 0;  //129 / 250 = 0
    16'b10000001_11111011 : OUT <= 0;  //129 / 251 = 0
    16'b10000001_11111100 : OUT <= 0;  //129 / 252 = 0
    16'b10000001_11111101 : OUT <= 0;  //129 / 253 = 0
    16'b10000001_11111110 : OUT <= 0;  //129 / 254 = 0
    16'b10000001_11111111 : OUT <= 0;  //129 / 255 = 0
    16'b10000010_00000000 : OUT <= 0;  //130 / 0 = 0
    16'b10000010_00000001 : OUT <= 130;  //130 / 1 = 130
    16'b10000010_00000010 : OUT <= 65;  //130 / 2 = 65
    16'b10000010_00000011 : OUT <= 43;  //130 / 3 = 43
    16'b10000010_00000100 : OUT <= 32;  //130 / 4 = 32
    16'b10000010_00000101 : OUT <= 26;  //130 / 5 = 26
    16'b10000010_00000110 : OUT <= 21;  //130 / 6 = 21
    16'b10000010_00000111 : OUT <= 18;  //130 / 7 = 18
    16'b10000010_00001000 : OUT <= 16;  //130 / 8 = 16
    16'b10000010_00001001 : OUT <= 14;  //130 / 9 = 14
    16'b10000010_00001010 : OUT <= 13;  //130 / 10 = 13
    16'b10000010_00001011 : OUT <= 11;  //130 / 11 = 11
    16'b10000010_00001100 : OUT <= 10;  //130 / 12 = 10
    16'b10000010_00001101 : OUT <= 10;  //130 / 13 = 10
    16'b10000010_00001110 : OUT <= 9;  //130 / 14 = 9
    16'b10000010_00001111 : OUT <= 8;  //130 / 15 = 8
    16'b10000010_00010000 : OUT <= 8;  //130 / 16 = 8
    16'b10000010_00010001 : OUT <= 7;  //130 / 17 = 7
    16'b10000010_00010010 : OUT <= 7;  //130 / 18 = 7
    16'b10000010_00010011 : OUT <= 6;  //130 / 19 = 6
    16'b10000010_00010100 : OUT <= 6;  //130 / 20 = 6
    16'b10000010_00010101 : OUT <= 6;  //130 / 21 = 6
    16'b10000010_00010110 : OUT <= 5;  //130 / 22 = 5
    16'b10000010_00010111 : OUT <= 5;  //130 / 23 = 5
    16'b10000010_00011000 : OUT <= 5;  //130 / 24 = 5
    16'b10000010_00011001 : OUT <= 5;  //130 / 25 = 5
    16'b10000010_00011010 : OUT <= 5;  //130 / 26 = 5
    16'b10000010_00011011 : OUT <= 4;  //130 / 27 = 4
    16'b10000010_00011100 : OUT <= 4;  //130 / 28 = 4
    16'b10000010_00011101 : OUT <= 4;  //130 / 29 = 4
    16'b10000010_00011110 : OUT <= 4;  //130 / 30 = 4
    16'b10000010_00011111 : OUT <= 4;  //130 / 31 = 4
    16'b10000010_00100000 : OUT <= 4;  //130 / 32 = 4
    16'b10000010_00100001 : OUT <= 3;  //130 / 33 = 3
    16'b10000010_00100010 : OUT <= 3;  //130 / 34 = 3
    16'b10000010_00100011 : OUT <= 3;  //130 / 35 = 3
    16'b10000010_00100100 : OUT <= 3;  //130 / 36 = 3
    16'b10000010_00100101 : OUT <= 3;  //130 / 37 = 3
    16'b10000010_00100110 : OUT <= 3;  //130 / 38 = 3
    16'b10000010_00100111 : OUT <= 3;  //130 / 39 = 3
    16'b10000010_00101000 : OUT <= 3;  //130 / 40 = 3
    16'b10000010_00101001 : OUT <= 3;  //130 / 41 = 3
    16'b10000010_00101010 : OUT <= 3;  //130 / 42 = 3
    16'b10000010_00101011 : OUT <= 3;  //130 / 43 = 3
    16'b10000010_00101100 : OUT <= 2;  //130 / 44 = 2
    16'b10000010_00101101 : OUT <= 2;  //130 / 45 = 2
    16'b10000010_00101110 : OUT <= 2;  //130 / 46 = 2
    16'b10000010_00101111 : OUT <= 2;  //130 / 47 = 2
    16'b10000010_00110000 : OUT <= 2;  //130 / 48 = 2
    16'b10000010_00110001 : OUT <= 2;  //130 / 49 = 2
    16'b10000010_00110010 : OUT <= 2;  //130 / 50 = 2
    16'b10000010_00110011 : OUT <= 2;  //130 / 51 = 2
    16'b10000010_00110100 : OUT <= 2;  //130 / 52 = 2
    16'b10000010_00110101 : OUT <= 2;  //130 / 53 = 2
    16'b10000010_00110110 : OUT <= 2;  //130 / 54 = 2
    16'b10000010_00110111 : OUT <= 2;  //130 / 55 = 2
    16'b10000010_00111000 : OUT <= 2;  //130 / 56 = 2
    16'b10000010_00111001 : OUT <= 2;  //130 / 57 = 2
    16'b10000010_00111010 : OUT <= 2;  //130 / 58 = 2
    16'b10000010_00111011 : OUT <= 2;  //130 / 59 = 2
    16'b10000010_00111100 : OUT <= 2;  //130 / 60 = 2
    16'b10000010_00111101 : OUT <= 2;  //130 / 61 = 2
    16'b10000010_00111110 : OUT <= 2;  //130 / 62 = 2
    16'b10000010_00111111 : OUT <= 2;  //130 / 63 = 2
    16'b10000010_01000000 : OUT <= 2;  //130 / 64 = 2
    16'b10000010_01000001 : OUT <= 2;  //130 / 65 = 2
    16'b10000010_01000010 : OUT <= 1;  //130 / 66 = 1
    16'b10000010_01000011 : OUT <= 1;  //130 / 67 = 1
    16'b10000010_01000100 : OUT <= 1;  //130 / 68 = 1
    16'b10000010_01000101 : OUT <= 1;  //130 / 69 = 1
    16'b10000010_01000110 : OUT <= 1;  //130 / 70 = 1
    16'b10000010_01000111 : OUT <= 1;  //130 / 71 = 1
    16'b10000010_01001000 : OUT <= 1;  //130 / 72 = 1
    16'b10000010_01001001 : OUT <= 1;  //130 / 73 = 1
    16'b10000010_01001010 : OUT <= 1;  //130 / 74 = 1
    16'b10000010_01001011 : OUT <= 1;  //130 / 75 = 1
    16'b10000010_01001100 : OUT <= 1;  //130 / 76 = 1
    16'b10000010_01001101 : OUT <= 1;  //130 / 77 = 1
    16'b10000010_01001110 : OUT <= 1;  //130 / 78 = 1
    16'b10000010_01001111 : OUT <= 1;  //130 / 79 = 1
    16'b10000010_01010000 : OUT <= 1;  //130 / 80 = 1
    16'b10000010_01010001 : OUT <= 1;  //130 / 81 = 1
    16'b10000010_01010010 : OUT <= 1;  //130 / 82 = 1
    16'b10000010_01010011 : OUT <= 1;  //130 / 83 = 1
    16'b10000010_01010100 : OUT <= 1;  //130 / 84 = 1
    16'b10000010_01010101 : OUT <= 1;  //130 / 85 = 1
    16'b10000010_01010110 : OUT <= 1;  //130 / 86 = 1
    16'b10000010_01010111 : OUT <= 1;  //130 / 87 = 1
    16'b10000010_01011000 : OUT <= 1;  //130 / 88 = 1
    16'b10000010_01011001 : OUT <= 1;  //130 / 89 = 1
    16'b10000010_01011010 : OUT <= 1;  //130 / 90 = 1
    16'b10000010_01011011 : OUT <= 1;  //130 / 91 = 1
    16'b10000010_01011100 : OUT <= 1;  //130 / 92 = 1
    16'b10000010_01011101 : OUT <= 1;  //130 / 93 = 1
    16'b10000010_01011110 : OUT <= 1;  //130 / 94 = 1
    16'b10000010_01011111 : OUT <= 1;  //130 / 95 = 1
    16'b10000010_01100000 : OUT <= 1;  //130 / 96 = 1
    16'b10000010_01100001 : OUT <= 1;  //130 / 97 = 1
    16'b10000010_01100010 : OUT <= 1;  //130 / 98 = 1
    16'b10000010_01100011 : OUT <= 1;  //130 / 99 = 1
    16'b10000010_01100100 : OUT <= 1;  //130 / 100 = 1
    16'b10000010_01100101 : OUT <= 1;  //130 / 101 = 1
    16'b10000010_01100110 : OUT <= 1;  //130 / 102 = 1
    16'b10000010_01100111 : OUT <= 1;  //130 / 103 = 1
    16'b10000010_01101000 : OUT <= 1;  //130 / 104 = 1
    16'b10000010_01101001 : OUT <= 1;  //130 / 105 = 1
    16'b10000010_01101010 : OUT <= 1;  //130 / 106 = 1
    16'b10000010_01101011 : OUT <= 1;  //130 / 107 = 1
    16'b10000010_01101100 : OUT <= 1;  //130 / 108 = 1
    16'b10000010_01101101 : OUT <= 1;  //130 / 109 = 1
    16'b10000010_01101110 : OUT <= 1;  //130 / 110 = 1
    16'b10000010_01101111 : OUT <= 1;  //130 / 111 = 1
    16'b10000010_01110000 : OUT <= 1;  //130 / 112 = 1
    16'b10000010_01110001 : OUT <= 1;  //130 / 113 = 1
    16'b10000010_01110010 : OUT <= 1;  //130 / 114 = 1
    16'b10000010_01110011 : OUT <= 1;  //130 / 115 = 1
    16'b10000010_01110100 : OUT <= 1;  //130 / 116 = 1
    16'b10000010_01110101 : OUT <= 1;  //130 / 117 = 1
    16'b10000010_01110110 : OUT <= 1;  //130 / 118 = 1
    16'b10000010_01110111 : OUT <= 1;  //130 / 119 = 1
    16'b10000010_01111000 : OUT <= 1;  //130 / 120 = 1
    16'b10000010_01111001 : OUT <= 1;  //130 / 121 = 1
    16'b10000010_01111010 : OUT <= 1;  //130 / 122 = 1
    16'b10000010_01111011 : OUT <= 1;  //130 / 123 = 1
    16'b10000010_01111100 : OUT <= 1;  //130 / 124 = 1
    16'b10000010_01111101 : OUT <= 1;  //130 / 125 = 1
    16'b10000010_01111110 : OUT <= 1;  //130 / 126 = 1
    16'b10000010_01111111 : OUT <= 1;  //130 / 127 = 1
    16'b10000010_10000000 : OUT <= 1;  //130 / 128 = 1
    16'b10000010_10000001 : OUT <= 1;  //130 / 129 = 1
    16'b10000010_10000010 : OUT <= 1;  //130 / 130 = 1
    16'b10000010_10000011 : OUT <= 0;  //130 / 131 = 0
    16'b10000010_10000100 : OUT <= 0;  //130 / 132 = 0
    16'b10000010_10000101 : OUT <= 0;  //130 / 133 = 0
    16'b10000010_10000110 : OUT <= 0;  //130 / 134 = 0
    16'b10000010_10000111 : OUT <= 0;  //130 / 135 = 0
    16'b10000010_10001000 : OUT <= 0;  //130 / 136 = 0
    16'b10000010_10001001 : OUT <= 0;  //130 / 137 = 0
    16'b10000010_10001010 : OUT <= 0;  //130 / 138 = 0
    16'b10000010_10001011 : OUT <= 0;  //130 / 139 = 0
    16'b10000010_10001100 : OUT <= 0;  //130 / 140 = 0
    16'b10000010_10001101 : OUT <= 0;  //130 / 141 = 0
    16'b10000010_10001110 : OUT <= 0;  //130 / 142 = 0
    16'b10000010_10001111 : OUT <= 0;  //130 / 143 = 0
    16'b10000010_10010000 : OUT <= 0;  //130 / 144 = 0
    16'b10000010_10010001 : OUT <= 0;  //130 / 145 = 0
    16'b10000010_10010010 : OUT <= 0;  //130 / 146 = 0
    16'b10000010_10010011 : OUT <= 0;  //130 / 147 = 0
    16'b10000010_10010100 : OUT <= 0;  //130 / 148 = 0
    16'b10000010_10010101 : OUT <= 0;  //130 / 149 = 0
    16'b10000010_10010110 : OUT <= 0;  //130 / 150 = 0
    16'b10000010_10010111 : OUT <= 0;  //130 / 151 = 0
    16'b10000010_10011000 : OUT <= 0;  //130 / 152 = 0
    16'b10000010_10011001 : OUT <= 0;  //130 / 153 = 0
    16'b10000010_10011010 : OUT <= 0;  //130 / 154 = 0
    16'b10000010_10011011 : OUT <= 0;  //130 / 155 = 0
    16'b10000010_10011100 : OUT <= 0;  //130 / 156 = 0
    16'b10000010_10011101 : OUT <= 0;  //130 / 157 = 0
    16'b10000010_10011110 : OUT <= 0;  //130 / 158 = 0
    16'b10000010_10011111 : OUT <= 0;  //130 / 159 = 0
    16'b10000010_10100000 : OUT <= 0;  //130 / 160 = 0
    16'b10000010_10100001 : OUT <= 0;  //130 / 161 = 0
    16'b10000010_10100010 : OUT <= 0;  //130 / 162 = 0
    16'b10000010_10100011 : OUT <= 0;  //130 / 163 = 0
    16'b10000010_10100100 : OUT <= 0;  //130 / 164 = 0
    16'b10000010_10100101 : OUT <= 0;  //130 / 165 = 0
    16'b10000010_10100110 : OUT <= 0;  //130 / 166 = 0
    16'b10000010_10100111 : OUT <= 0;  //130 / 167 = 0
    16'b10000010_10101000 : OUT <= 0;  //130 / 168 = 0
    16'b10000010_10101001 : OUT <= 0;  //130 / 169 = 0
    16'b10000010_10101010 : OUT <= 0;  //130 / 170 = 0
    16'b10000010_10101011 : OUT <= 0;  //130 / 171 = 0
    16'b10000010_10101100 : OUT <= 0;  //130 / 172 = 0
    16'b10000010_10101101 : OUT <= 0;  //130 / 173 = 0
    16'b10000010_10101110 : OUT <= 0;  //130 / 174 = 0
    16'b10000010_10101111 : OUT <= 0;  //130 / 175 = 0
    16'b10000010_10110000 : OUT <= 0;  //130 / 176 = 0
    16'b10000010_10110001 : OUT <= 0;  //130 / 177 = 0
    16'b10000010_10110010 : OUT <= 0;  //130 / 178 = 0
    16'b10000010_10110011 : OUT <= 0;  //130 / 179 = 0
    16'b10000010_10110100 : OUT <= 0;  //130 / 180 = 0
    16'b10000010_10110101 : OUT <= 0;  //130 / 181 = 0
    16'b10000010_10110110 : OUT <= 0;  //130 / 182 = 0
    16'b10000010_10110111 : OUT <= 0;  //130 / 183 = 0
    16'b10000010_10111000 : OUT <= 0;  //130 / 184 = 0
    16'b10000010_10111001 : OUT <= 0;  //130 / 185 = 0
    16'b10000010_10111010 : OUT <= 0;  //130 / 186 = 0
    16'b10000010_10111011 : OUT <= 0;  //130 / 187 = 0
    16'b10000010_10111100 : OUT <= 0;  //130 / 188 = 0
    16'b10000010_10111101 : OUT <= 0;  //130 / 189 = 0
    16'b10000010_10111110 : OUT <= 0;  //130 / 190 = 0
    16'b10000010_10111111 : OUT <= 0;  //130 / 191 = 0
    16'b10000010_11000000 : OUT <= 0;  //130 / 192 = 0
    16'b10000010_11000001 : OUT <= 0;  //130 / 193 = 0
    16'b10000010_11000010 : OUT <= 0;  //130 / 194 = 0
    16'b10000010_11000011 : OUT <= 0;  //130 / 195 = 0
    16'b10000010_11000100 : OUT <= 0;  //130 / 196 = 0
    16'b10000010_11000101 : OUT <= 0;  //130 / 197 = 0
    16'b10000010_11000110 : OUT <= 0;  //130 / 198 = 0
    16'b10000010_11000111 : OUT <= 0;  //130 / 199 = 0
    16'b10000010_11001000 : OUT <= 0;  //130 / 200 = 0
    16'b10000010_11001001 : OUT <= 0;  //130 / 201 = 0
    16'b10000010_11001010 : OUT <= 0;  //130 / 202 = 0
    16'b10000010_11001011 : OUT <= 0;  //130 / 203 = 0
    16'b10000010_11001100 : OUT <= 0;  //130 / 204 = 0
    16'b10000010_11001101 : OUT <= 0;  //130 / 205 = 0
    16'b10000010_11001110 : OUT <= 0;  //130 / 206 = 0
    16'b10000010_11001111 : OUT <= 0;  //130 / 207 = 0
    16'b10000010_11010000 : OUT <= 0;  //130 / 208 = 0
    16'b10000010_11010001 : OUT <= 0;  //130 / 209 = 0
    16'b10000010_11010010 : OUT <= 0;  //130 / 210 = 0
    16'b10000010_11010011 : OUT <= 0;  //130 / 211 = 0
    16'b10000010_11010100 : OUT <= 0;  //130 / 212 = 0
    16'b10000010_11010101 : OUT <= 0;  //130 / 213 = 0
    16'b10000010_11010110 : OUT <= 0;  //130 / 214 = 0
    16'b10000010_11010111 : OUT <= 0;  //130 / 215 = 0
    16'b10000010_11011000 : OUT <= 0;  //130 / 216 = 0
    16'b10000010_11011001 : OUT <= 0;  //130 / 217 = 0
    16'b10000010_11011010 : OUT <= 0;  //130 / 218 = 0
    16'b10000010_11011011 : OUT <= 0;  //130 / 219 = 0
    16'b10000010_11011100 : OUT <= 0;  //130 / 220 = 0
    16'b10000010_11011101 : OUT <= 0;  //130 / 221 = 0
    16'b10000010_11011110 : OUT <= 0;  //130 / 222 = 0
    16'b10000010_11011111 : OUT <= 0;  //130 / 223 = 0
    16'b10000010_11100000 : OUT <= 0;  //130 / 224 = 0
    16'b10000010_11100001 : OUT <= 0;  //130 / 225 = 0
    16'b10000010_11100010 : OUT <= 0;  //130 / 226 = 0
    16'b10000010_11100011 : OUT <= 0;  //130 / 227 = 0
    16'b10000010_11100100 : OUT <= 0;  //130 / 228 = 0
    16'b10000010_11100101 : OUT <= 0;  //130 / 229 = 0
    16'b10000010_11100110 : OUT <= 0;  //130 / 230 = 0
    16'b10000010_11100111 : OUT <= 0;  //130 / 231 = 0
    16'b10000010_11101000 : OUT <= 0;  //130 / 232 = 0
    16'b10000010_11101001 : OUT <= 0;  //130 / 233 = 0
    16'b10000010_11101010 : OUT <= 0;  //130 / 234 = 0
    16'b10000010_11101011 : OUT <= 0;  //130 / 235 = 0
    16'b10000010_11101100 : OUT <= 0;  //130 / 236 = 0
    16'b10000010_11101101 : OUT <= 0;  //130 / 237 = 0
    16'b10000010_11101110 : OUT <= 0;  //130 / 238 = 0
    16'b10000010_11101111 : OUT <= 0;  //130 / 239 = 0
    16'b10000010_11110000 : OUT <= 0;  //130 / 240 = 0
    16'b10000010_11110001 : OUT <= 0;  //130 / 241 = 0
    16'b10000010_11110010 : OUT <= 0;  //130 / 242 = 0
    16'b10000010_11110011 : OUT <= 0;  //130 / 243 = 0
    16'b10000010_11110100 : OUT <= 0;  //130 / 244 = 0
    16'b10000010_11110101 : OUT <= 0;  //130 / 245 = 0
    16'b10000010_11110110 : OUT <= 0;  //130 / 246 = 0
    16'b10000010_11110111 : OUT <= 0;  //130 / 247 = 0
    16'b10000010_11111000 : OUT <= 0;  //130 / 248 = 0
    16'b10000010_11111001 : OUT <= 0;  //130 / 249 = 0
    16'b10000010_11111010 : OUT <= 0;  //130 / 250 = 0
    16'b10000010_11111011 : OUT <= 0;  //130 / 251 = 0
    16'b10000010_11111100 : OUT <= 0;  //130 / 252 = 0
    16'b10000010_11111101 : OUT <= 0;  //130 / 253 = 0
    16'b10000010_11111110 : OUT <= 0;  //130 / 254 = 0
    16'b10000010_11111111 : OUT <= 0;  //130 / 255 = 0
    16'b10000011_00000000 : OUT <= 0;  //131 / 0 = 0
    16'b10000011_00000001 : OUT <= 131;  //131 / 1 = 131
    16'b10000011_00000010 : OUT <= 65;  //131 / 2 = 65
    16'b10000011_00000011 : OUT <= 43;  //131 / 3 = 43
    16'b10000011_00000100 : OUT <= 32;  //131 / 4 = 32
    16'b10000011_00000101 : OUT <= 26;  //131 / 5 = 26
    16'b10000011_00000110 : OUT <= 21;  //131 / 6 = 21
    16'b10000011_00000111 : OUT <= 18;  //131 / 7 = 18
    16'b10000011_00001000 : OUT <= 16;  //131 / 8 = 16
    16'b10000011_00001001 : OUT <= 14;  //131 / 9 = 14
    16'b10000011_00001010 : OUT <= 13;  //131 / 10 = 13
    16'b10000011_00001011 : OUT <= 11;  //131 / 11 = 11
    16'b10000011_00001100 : OUT <= 10;  //131 / 12 = 10
    16'b10000011_00001101 : OUT <= 10;  //131 / 13 = 10
    16'b10000011_00001110 : OUT <= 9;  //131 / 14 = 9
    16'b10000011_00001111 : OUT <= 8;  //131 / 15 = 8
    16'b10000011_00010000 : OUT <= 8;  //131 / 16 = 8
    16'b10000011_00010001 : OUT <= 7;  //131 / 17 = 7
    16'b10000011_00010010 : OUT <= 7;  //131 / 18 = 7
    16'b10000011_00010011 : OUT <= 6;  //131 / 19 = 6
    16'b10000011_00010100 : OUT <= 6;  //131 / 20 = 6
    16'b10000011_00010101 : OUT <= 6;  //131 / 21 = 6
    16'b10000011_00010110 : OUT <= 5;  //131 / 22 = 5
    16'b10000011_00010111 : OUT <= 5;  //131 / 23 = 5
    16'b10000011_00011000 : OUT <= 5;  //131 / 24 = 5
    16'b10000011_00011001 : OUT <= 5;  //131 / 25 = 5
    16'b10000011_00011010 : OUT <= 5;  //131 / 26 = 5
    16'b10000011_00011011 : OUT <= 4;  //131 / 27 = 4
    16'b10000011_00011100 : OUT <= 4;  //131 / 28 = 4
    16'b10000011_00011101 : OUT <= 4;  //131 / 29 = 4
    16'b10000011_00011110 : OUT <= 4;  //131 / 30 = 4
    16'b10000011_00011111 : OUT <= 4;  //131 / 31 = 4
    16'b10000011_00100000 : OUT <= 4;  //131 / 32 = 4
    16'b10000011_00100001 : OUT <= 3;  //131 / 33 = 3
    16'b10000011_00100010 : OUT <= 3;  //131 / 34 = 3
    16'b10000011_00100011 : OUT <= 3;  //131 / 35 = 3
    16'b10000011_00100100 : OUT <= 3;  //131 / 36 = 3
    16'b10000011_00100101 : OUT <= 3;  //131 / 37 = 3
    16'b10000011_00100110 : OUT <= 3;  //131 / 38 = 3
    16'b10000011_00100111 : OUT <= 3;  //131 / 39 = 3
    16'b10000011_00101000 : OUT <= 3;  //131 / 40 = 3
    16'b10000011_00101001 : OUT <= 3;  //131 / 41 = 3
    16'b10000011_00101010 : OUT <= 3;  //131 / 42 = 3
    16'b10000011_00101011 : OUT <= 3;  //131 / 43 = 3
    16'b10000011_00101100 : OUT <= 2;  //131 / 44 = 2
    16'b10000011_00101101 : OUT <= 2;  //131 / 45 = 2
    16'b10000011_00101110 : OUT <= 2;  //131 / 46 = 2
    16'b10000011_00101111 : OUT <= 2;  //131 / 47 = 2
    16'b10000011_00110000 : OUT <= 2;  //131 / 48 = 2
    16'b10000011_00110001 : OUT <= 2;  //131 / 49 = 2
    16'b10000011_00110010 : OUT <= 2;  //131 / 50 = 2
    16'b10000011_00110011 : OUT <= 2;  //131 / 51 = 2
    16'b10000011_00110100 : OUT <= 2;  //131 / 52 = 2
    16'b10000011_00110101 : OUT <= 2;  //131 / 53 = 2
    16'b10000011_00110110 : OUT <= 2;  //131 / 54 = 2
    16'b10000011_00110111 : OUT <= 2;  //131 / 55 = 2
    16'b10000011_00111000 : OUT <= 2;  //131 / 56 = 2
    16'b10000011_00111001 : OUT <= 2;  //131 / 57 = 2
    16'b10000011_00111010 : OUT <= 2;  //131 / 58 = 2
    16'b10000011_00111011 : OUT <= 2;  //131 / 59 = 2
    16'b10000011_00111100 : OUT <= 2;  //131 / 60 = 2
    16'b10000011_00111101 : OUT <= 2;  //131 / 61 = 2
    16'b10000011_00111110 : OUT <= 2;  //131 / 62 = 2
    16'b10000011_00111111 : OUT <= 2;  //131 / 63 = 2
    16'b10000011_01000000 : OUT <= 2;  //131 / 64 = 2
    16'b10000011_01000001 : OUT <= 2;  //131 / 65 = 2
    16'b10000011_01000010 : OUT <= 1;  //131 / 66 = 1
    16'b10000011_01000011 : OUT <= 1;  //131 / 67 = 1
    16'b10000011_01000100 : OUT <= 1;  //131 / 68 = 1
    16'b10000011_01000101 : OUT <= 1;  //131 / 69 = 1
    16'b10000011_01000110 : OUT <= 1;  //131 / 70 = 1
    16'b10000011_01000111 : OUT <= 1;  //131 / 71 = 1
    16'b10000011_01001000 : OUT <= 1;  //131 / 72 = 1
    16'b10000011_01001001 : OUT <= 1;  //131 / 73 = 1
    16'b10000011_01001010 : OUT <= 1;  //131 / 74 = 1
    16'b10000011_01001011 : OUT <= 1;  //131 / 75 = 1
    16'b10000011_01001100 : OUT <= 1;  //131 / 76 = 1
    16'b10000011_01001101 : OUT <= 1;  //131 / 77 = 1
    16'b10000011_01001110 : OUT <= 1;  //131 / 78 = 1
    16'b10000011_01001111 : OUT <= 1;  //131 / 79 = 1
    16'b10000011_01010000 : OUT <= 1;  //131 / 80 = 1
    16'b10000011_01010001 : OUT <= 1;  //131 / 81 = 1
    16'b10000011_01010010 : OUT <= 1;  //131 / 82 = 1
    16'b10000011_01010011 : OUT <= 1;  //131 / 83 = 1
    16'b10000011_01010100 : OUT <= 1;  //131 / 84 = 1
    16'b10000011_01010101 : OUT <= 1;  //131 / 85 = 1
    16'b10000011_01010110 : OUT <= 1;  //131 / 86 = 1
    16'b10000011_01010111 : OUT <= 1;  //131 / 87 = 1
    16'b10000011_01011000 : OUT <= 1;  //131 / 88 = 1
    16'b10000011_01011001 : OUT <= 1;  //131 / 89 = 1
    16'b10000011_01011010 : OUT <= 1;  //131 / 90 = 1
    16'b10000011_01011011 : OUT <= 1;  //131 / 91 = 1
    16'b10000011_01011100 : OUT <= 1;  //131 / 92 = 1
    16'b10000011_01011101 : OUT <= 1;  //131 / 93 = 1
    16'b10000011_01011110 : OUT <= 1;  //131 / 94 = 1
    16'b10000011_01011111 : OUT <= 1;  //131 / 95 = 1
    16'b10000011_01100000 : OUT <= 1;  //131 / 96 = 1
    16'b10000011_01100001 : OUT <= 1;  //131 / 97 = 1
    16'b10000011_01100010 : OUT <= 1;  //131 / 98 = 1
    16'b10000011_01100011 : OUT <= 1;  //131 / 99 = 1
    16'b10000011_01100100 : OUT <= 1;  //131 / 100 = 1
    16'b10000011_01100101 : OUT <= 1;  //131 / 101 = 1
    16'b10000011_01100110 : OUT <= 1;  //131 / 102 = 1
    16'b10000011_01100111 : OUT <= 1;  //131 / 103 = 1
    16'b10000011_01101000 : OUT <= 1;  //131 / 104 = 1
    16'b10000011_01101001 : OUT <= 1;  //131 / 105 = 1
    16'b10000011_01101010 : OUT <= 1;  //131 / 106 = 1
    16'b10000011_01101011 : OUT <= 1;  //131 / 107 = 1
    16'b10000011_01101100 : OUT <= 1;  //131 / 108 = 1
    16'b10000011_01101101 : OUT <= 1;  //131 / 109 = 1
    16'b10000011_01101110 : OUT <= 1;  //131 / 110 = 1
    16'b10000011_01101111 : OUT <= 1;  //131 / 111 = 1
    16'b10000011_01110000 : OUT <= 1;  //131 / 112 = 1
    16'b10000011_01110001 : OUT <= 1;  //131 / 113 = 1
    16'b10000011_01110010 : OUT <= 1;  //131 / 114 = 1
    16'b10000011_01110011 : OUT <= 1;  //131 / 115 = 1
    16'b10000011_01110100 : OUT <= 1;  //131 / 116 = 1
    16'b10000011_01110101 : OUT <= 1;  //131 / 117 = 1
    16'b10000011_01110110 : OUT <= 1;  //131 / 118 = 1
    16'b10000011_01110111 : OUT <= 1;  //131 / 119 = 1
    16'b10000011_01111000 : OUT <= 1;  //131 / 120 = 1
    16'b10000011_01111001 : OUT <= 1;  //131 / 121 = 1
    16'b10000011_01111010 : OUT <= 1;  //131 / 122 = 1
    16'b10000011_01111011 : OUT <= 1;  //131 / 123 = 1
    16'b10000011_01111100 : OUT <= 1;  //131 / 124 = 1
    16'b10000011_01111101 : OUT <= 1;  //131 / 125 = 1
    16'b10000011_01111110 : OUT <= 1;  //131 / 126 = 1
    16'b10000011_01111111 : OUT <= 1;  //131 / 127 = 1
    16'b10000011_10000000 : OUT <= 1;  //131 / 128 = 1
    16'b10000011_10000001 : OUT <= 1;  //131 / 129 = 1
    16'b10000011_10000010 : OUT <= 1;  //131 / 130 = 1
    16'b10000011_10000011 : OUT <= 1;  //131 / 131 = 1
    16'b10000011_10000100 : OUT <= 0;  //131 / 132 = 0
    16'b10000011_10000101 : OUT <= 0;  //131 / 133 = 0
    16'b10000011_10000110 : OUT <= 0;  //131 / 134 = 0
    16'b10000011_10000111 : OUT <= 0;  //131 / 135 = 0
    16'b10000011_10001000 : OUT <= 0;  //131 / 136 = 0
    16'b10000011_10001001 : OUT <= 0;  //131 / 137 = 0
    16'b10000011_10001010 : OUT <= 0;  //131 / 138 = 0
    16'b10000011_10001011 : OUT <= 0;  //131 / 139 = 0
    16'b10000011_10001100 : OUT <= 0;  //131 / 140 = 0
    16'b10000011_10001101 : OUT <= 0;  //131 / 141 = 0
    16'b10000011_10001110 : OUT <= 0;  //131 / 142 = 0
    16'b10000011_10001111 : OUT <= 0;  //131 / 143 = 0
    16'b10000011_10010000 : OUT <= 0;  //131 / 144 = 0
    16'b10000011_10010001 : OUT <= 0;  //131 / 145 = 0
    16'b10000011_10010010 : OUT <= 0;  //131 / 146 = 0
    16'b10000011_10010011 : OUT <= 0;  //131 / 147 = 0
    16'b10000011_10010100 : OUT <= 0;  //131 / 148 = 0
    16'b10000011_10010101 : OUT <= 0;  //131 / 149 = 0
    16'b10000011_10010110 : OUT <= 0;  //131 / 150 = 0
    16'b10000011_10010111 : OUT <= 0;  //131 / 151 = 0
    16'b10000011_10011000 : OUT <= 0;  //131 / 152 = 0
    16'b10000011_10011001 : OUT <= 0;  //131 / 153 = 0
    16'b10000011_10011010 : OUT <= 0;  //131 / 154 = 0
    16'b10000011_10011011 : OUT <= 0;  //131 / 155 = 0
    16'b10000011_10011100 : OUT <= 0;  //131 / 156 = 0
    16'b10000011_10011101 : OUT <= 0;  //131 / 157 = 0
    16'b10000011_10011110 : OUT <= 0;  //131 / 158 = 0
    16'b10000011_10011111 : OUT <= 0;  //131 / 159 = 0
    16'b10000011_10100000 : OUT <= 0;  //131 / 160 = 0
    16'b10000011_10100001 : OUT <= 0;  //131 / 161 = 0
    16'b10000011_10100010 : OUT <= 0;  //131 / 162 = 0
    16'b10000011_10100011 : OUT <= 0;  //131 / 163 = 0
    16'b10000011_10100100 : OUT <= 0;  //131 / 164 = 0
    16'b10000011_10100101 : OUT <= 0;  //131 / 165 = 0
    16'b10000011_10100110 : OUT <= 0;  //131 / 166 = 0
    16'b10000011_10100111 : OUT <= 0;  //131 / 167 = 0
    16'b10000011_10101000 : OUT <= 0;  //131 / 168 = 0
    16'b10000011_10101001 : OUT <= 0;  //131 / 169 = 0
    16'b10000011_10101010 : OUT <= 0;  //131 / 170 = 0
    16'b10000011_10101011 : OUT <= 0;  //131 / 171 = 0
    16'b10000011_10101100 : OUT <= 0;  //131 / 172 = 0
    16'b10000011_10101101 : OUT <= 0;  //131 / 173 = 0
    16'b10000011_10101110 : OUT <= 0;  //131 / 174 = 0
    16'b10000011_10101111 : OUT <= 0;  //131 / 175 = 0
    16'b10000011_10110000 : OUT <= 0;  //131 / 176 = 0
    16'b10000011_10110001 : OUT <= 0;  //131 / 177 = 0
    16'b10000011_10110010 : OUT <= 0;  //131 / 178 = 0
    16'b10000011_10110011 : OUT <= 0;  //131 / 179 = 0
    16'b10000011_10110100 : OUT <= 0;  //131 / 180 = 0
    16'b10000011_10110101 : OUT <= 0;  //131 / 181 = 0
    16'b10000011_10110110 : OUT <= 0;  //131 / 182 = 0
    16'b10000011_10110111 : OUT <= 0;  //131 / 183 = 0
    16'b10000011_10111000 : OUT <= 0;  //131 / 184 = 0
    16'b10000011_10111001 : OUT <= 0;  //131 / 185 = 0
    16'b10000011_10111010 : OUT <= 0;  //131 / 186 = 0
    16'b10000011_10111011 : OUT <= 0;  //131 / 187 = 0
    16'b10000011_10111100 : OUT <= 0;  //131 / 188 = 0
    16'b10000011_10111101 : OUT <= 0;  //131 / 189 = 0
    16'b10000011_10111110 : OUT <= 0;  //131 / 190 = 0
    16'b10000011_10111111 : OUT <= 0;  //131 / 191 = 0
    16'b10000011_11000000 : OUT <= 0;  //131 / 192 = 0
    16'b10000011_11000001 : OUT <= 0;  //131 / 193 = 0
    16'b10000011_11000010 : OUT <= 0;  //131 / 194 = 0
    16'b10000011_11000011 : OUT <= 0;  //131 / 195 = 0
    16'b10000011_11000100 : OUT <= 0;  //131 / 196 = 0
    16'b10000011_11000101 : OUT <= 0;  //131 / 197 = 0
    16'b10000011_11000110 : OUT <= 0;  //131 / 198 = 0
    16'b10000011_11000111 : OUT <= 0;  //131 / 199 = 0
    16'b10000011_11001000 : OUT <= 0;  //131 / 200 = 0
    16'b10000011_11001001 : OUT <= 0;  //131 / 201 = 0
    16'b10000011_11001010 : OUT <= 0;  //131 / 202 = 0
    16'b10000011_11001011 : OUT <= 0;  //131 / 203 = 0
    16'b10000011_11001100 : OUT <= 0;  //131 / 204 = 0
    16'b10000011_11001101 : OUT <= 0;  //131 / 205 = 0
    16'b10000011_11001110 : OUT <= 0;  //131 / 206 = 0
    16'b10000011_11001111 : OUT <= 0;  //131 / 207 = 0
    16'b10000011_11010000 : OUT <= 0;  //131 / 208 = 0
    16'b10000011_11010001 : OUT <= 0;  //131 / 209 = 0
    16'b10000011_11010010 : OUT <= 0;  //131 / 210 = 0
    16'b10000011_11010011 : OUT <= 0;  //131 / 211 = 0
    16'b10000011_11010100 : OUT <= 0;  //131 / 212 = 0
    16'b10000011_11010101 : OUT <= 0;  //131 / 213 = 0
    16'b10000011_11010110 : OUT <= 0;  //131 / 214 = 0
    16'b10000011_11010111 : OUT <= 0;  //131 / 215 = 0
    16'b10000011_11011000 : OUT <= 0;  //131 / 216 = 0
    16'b10000011_11011001 : OUT <= 0;  //131 / 217 = 0
    16'b10000011_11011010 : OUT <= 0;  //131 / 218 = 0
    16'b10000011_11011011 : OUT <= 0;  //131 / 219 = 0
    16'b10000011_11011100 : OUT <= 0;  //131 / 220 = 0
    16'b10000011_11011101 : OUT <= 0;  //131 / 221 = 0
    16'b10000011_11011110 : OUT <= 0;  //131 / 222 = 0
    16'b10000011_11011111 : OUT <= 0;  //131 / 223 = 0
    16'b10000011_11100000 : OUT <= 0;  //131 / 224 = 0
    16'b10000011_11100001 : OUT <= 0;  //131 / 225 = 0
    16'b10000011_11100010 : OUT <= 0;  //131 / 226 = 0
    16'b10000011_11100011 : OUT <= 0;  //131 / 227 = 0
    16'b10000011_11100100 : OUT <= 0;  //131 / 228 = 0
    16'b10000011_11100101 : OUT <= 0;  //131 / 229 = 0
    16'b10000011_11100110 : OUT <= 0;  //131 / 230 = 0
    16'b10000011_11100111 : OUT <= 0;  //131 / 231 = 0
    16'b10000011_11101000 : OUT <= 0;  //131 / 232 = 0
    16'b10000011_11101001 : OUT <= 0;  //131 / 233 = 0
    16'b10000011_11101010 : OUT <= 0;  //131 / 234 = 0
    16'b10000011_11101011 : OUT <= 0;  //131 / 235 = 0
    16'b10000011_11101100 : OUT <= 0;  //131 / 236 = 0
    16'b10000011_11101101 : OUT <= 0;  //131 / 237 = 0
    16'b10000011_11101110 : OUT <= 0;  //131 / 238 = 0
    16'b10000011_11101111 : OUT <= 0;  //131 / 239 = 0
    16'b10000011_11110000 : OUT <= 0;  //131 / 240 = 0
    16'b10000011_11110001 : OUT <= 0;  //131 / 241 = 0
    16'b10000011_11110010 : OUT <= 0;  //131 / 242 = 0
    16'b10000011_11110011 : OUT <= 0;  //131 / 243 = 0
    16'b10000011_11110100 : OUT <= 0;  //131 / 244 = 0
    16'b10000011_11110101 : OUT <= 0;  //131 / 245 = 0
    16'b10000011_11110110 : OUT <= 0;  //131 / 246 = 0
    16'b10000011_11110111 : OUT <= 0;  //131 / 247 = 0
    16'b10000011_11111000 : OUT <= 0;  //131 / 248 = 0
    16'b10000011_11111001 : OUT <= 0;  //131 / 249 = 0
    16'b10000011_11111010 : OUT <= 0;  //131 / 250 = 0
    16'b10000011_11111011 : OUT <= 0;  //131 / 251 = 0
    16'b10000011_11111100 : OUT <= 0;  //131 / 252 = 0
    16'b10000011_11111101 : OUT <= 0;  //131 / 253 = 0
    16'b10000011_11111110 : OUT <= 0;  //131 / 254 = 0
    16'b10000011_11111111 : OUT <= 0;  //131 / 255 = 0
    16'b10000100_00000000 : OUT <= 0;  //132 / 0 = 0
    16'b10000100_00000001 : OUT <= 132;  //132 / 1 = 132
    16'b10000100_00000010 : OUT <= 66;  //132 / 2 = 66
    16'b10000100_00000011 : OUT <= 44;  //132 / 3 = 44
    16'b10000100_00000100 : OUT <= 33;  //132 / 4 = 33
    16'b10000100_00000101 : OUT <= 26;  //132 / 5 = 26
    16'b10000100_00000110 : OUT <= 22;  //132 / 6 = 22
    16'b10000100_00000111 : OUT <= 18;  //132 / 7 = 18
    16'b10000100_00001000 : OUT <= 16;  //132 / 8 = 16
    16'b10000100_00001001 : OUT <= 14;  //132 / 9 = 14
    16'b10000100_00001010 : OUT <= 13;  //132 / 10 = 13
    16'b10000100_00001011 : OUT <= 12;  //132 / 11 = 12
    16'b10000100_00001100 : OUT <= 11;  //132 / 12 = 11
    16'b10000100_00001101 : OUT <= 10;  //132 / 13 = 10
    16'b10000100_00001110 : OUT <= 9;  //132 / 14 = 9
    16'b10000100_00001111 : OUT <= 8;  //132 / 15 = 8
    16'b10000100_00010000 : OUT <= 8;  //132 / 16 = 8
    16'b10000100_00010001 : OUT <= 7;  //132 / 17 = 7
    16'b10000100_00010010 : OUT <= 7;  //132 / 18 = 7
    16'b10000100_00010011 : OUT <= 6;  //132 / 19 = 6
    16'b10000100_00010100 : OUT <= 6;  //132 / 20 = 6
    16'b10000100_00010101 : OUT <= 6;  //132 / 21 = 6
    16'b10000100_00010110 : OUT <= 6;  //132 / 22 = 6
    16'b10000100_00010111 : OUT <= 5;  //132 / 23 = 5
    16'b10000100_00011000 : OUT <= 5;  //132 / 24 = 5
    16'b10000100_00011001 : OUT <= 5;  //132 / 25 = 5
    16'b10000100_00011010 : OUT <= 5;  //132 / 26 = 5
    16'b10000100_00011011 : OUT <= 4;  //132 / 27 = 4
    16'b10000100_00011100 : OUT <= 4;  //132 / 28 = 4
    16'b10000100_00011101 : OUT <= 4;  //132 / 29 = 4
    16'b10000100_00011110 : OUT <= 4;  //132 / 30 = 4
    16'b10000100_00011111 : OUT <= 4;  //132 / 31 = 4
    16'b10000100_00100000 : OUT <= 4;  //132 / 32 = 4
    16'b10000100_00100001 : OUT <= 4;  //132 / 33 = 4
    16'b10000100_00100010 : OUT <= 3;  //132 / 34 = 3
    16'b10000100_00100011 : OUT <= 3;  //132 / 35 = 3
    16'b10000100_00100100 : OUT <= 3;  //132 / 36 = 3
    16'b10000100_00100101 : OUT <= 3;  //132 / 37 = 3
    16'b10000100_00100110 : OUT <= 3;  //132 / 38 = 3
    16'b10000100_00100111 : OUT <= 3;  //132 / 39 = 3
    16'b10000100_00101000 : OUT <= 3;  //132 / 40 = 3
    16'b10000100_00101001 : OUT <= 3;  //132 / 41 = 3
    16'b10000100_00101010 : OUT <= 3;  //132 / 42 = 3
    16'b10000100_00101011 : OUT <= 3;  //132 / 43 = 3
    16'b10000100_00101100 : OUT <= 3;  //132 / 44 = 3
    16'b10000100_00101101 : OUT <= 2;  //132 / 45 = 2
    16'b10000100_00101110 : OUT <= 2;  //132 / 46 = 2
    16'b10000100_00101111 : OUT <= 2;  //132 / 47 = 2
    16'b10000100_00110000 : OUT <= 2;  //132 / 48 = 2
    16'b10000100_00110001 : OUT <= 2;  //132 / 49 = 2
    16'b10000100_00110010 : OUT <= 2;  //132 / 50 = 2
    16'b10000100_00110011 : OUT <= 2;  //132 / 51 = 2
    16'b10000100_00110100 : OUT <= 2;  //132 / 52 = 2
    16'b10000100_00110101 : OUT <= 2;  //132 / 53 = 2
    16'b10000100_00110110 : OUT <= 2;  //132 / 54 = 2
    16'b10000100_00110111 : OUT <= 2;  //132 / 55 = 2
    16'b10000100_00111000 : OUT <= 2;  //132 / 56 = 2
    16'b10000100_00111001 : OUT <= 2;  //132 / 57 = 2
    16'b10000100_00111010 : OUT <= 2;  //132 / 58 = 2
    16'b10000100_00111011 : OUT <= 2;  //132 / 59 = 2
    16'b10000100_00111100 : OUT <= 2;  //132 / 60 = 2
    16'b10000100_00111101 : OUT <= 2;  //132 / 61 = 2
    16'b10000100_00111110 : OUT <= 2;  //132 / 62 = 2
    16'b10000100_00111111 : OUT <= 2;  //132 / 63 = 2
    16'b10000100_01000000 : OUT <= 2;  //132 / 64 = 2
    16'b10000100_01000001 : OUT <= 2;  //132 / 65 = 2
    16'b10000100_01000010 : OUT <= 2;  //132 / 66 = 2
    16'b10000100_01000011 : OUT <= 1;  //132 / 67 = 1
    16'b10000100_01000100 : OUT <= 1;  //132 / 68 = 1
    16'b10000100_01000101 : OUT <= 1;  //132 / 69 = 1
    16'b10000100_01000110 : OUT <= 1;  //132 / 70 = 1
    16'b10000100_01000111 : OUT <= 1;  //132 / 71 = 1
    16'b10000100_01001000 : OUT <= 1;  //132 / 72 = 1
    16'b10000100_01001001 : OUT <= 1;  //132 / 73 = 1
    16'b10000100_01001010 : OUT <= 1;  //132 / 74 = 1
    16'b10000100_01001011 : OUT <= 1;  //132 / 75 = 1
    16'b10000100_01001100 : OUT <= 1;  //132 / 76 = 1
    16'b10000100_01001101 : OUT <= 1;  //132 / 77 = 1
    16'b10000100_01001110 : OUT <= 1;  //132 / 78 = 1
    16'b10000100_01001111 : OUT <= 1;  //132 / 79 = 1
    16'b10000100_01010000 : OUT <= 1;  //132 / 80 = 1
    16'b10000100_01010001 : OUT <= 1;  //132 / 81 = 1
    16'b10000100_01010010 : OUT <= 1;  //132 / 82 = 1
    16'b10000100_01010011 : OUT <= 1;  //132 / 83 = 1
    16'b10000100_01010100 : OUT <= 1;  //132 / 84 = 1
    16'b10000100_01010101 : OUT <= 1;  //132 / 85 = 1
    16'b10000100_01010110 : OUT <= 1;  //132 / 86 = 1
    16'b10000100_01010111 : OUT <= 1;  //132 / 87 = 1
    16'b10000100_01011000 : OUT <= 1;  //132 / 88 = 1
    16'b10000100_01011001 : OUT <= 1;  //132 / 89 = 1
    16'b10000100_01011010 : OUT <= 1;  //132 / 90 = 1
    16'b10000100_01011011 : OUT <= 1;  //132 / 91 = 1
    16'b10000100_01011100 : OUT <= 1;  //132 / 92 = 1
    16'b10000100_01011101 : OUT <= 1;  //132 / 93 = 1
    16'b10000100_01011110 : OUT <= 1;  //132 / 94 = 1
    16'b10000100_01011111 : OUT <= 1;  //132 / 95 = 1
    16'b10000100_01100000 : OUT <= 1;  //132 / 96 = 1
    16'b10000100_01100001 : OUT <= 1;  //132 / 97 = 1
    16'b10000100_01100010 : OUT <= 1;  //132 / 98 = 1
    16'b10000100_01100011 : OUT <= 1;  //132 / 99 = 1
    16'b10000100_01100100 : OUT <= 1;  //132 / 100 = 1
    16'b10000100_01100101 : OUT <= 1;  //132 / 101 = 1
    16'b10000100_01100110 : OUT <= 1;  //132 / 102 = 1
    16'b10000100_01100111 : OUT <= 1;  //132 / 103 = 1
    16'b10000100_01101000 : OUT <= 1;  //132 / 104 = 1
    16'b10000100_01101001 : OUT <= 1;  //132 / 105 = 1
    16'b10000100_01101010 : OUT <= 1;  //132 / 106 = 1
    16'b10000100_01101011 : OUT <= 1;  //132 / 107 = 1
    16'b10000100_01101100 : OUT <= 1;  //132 / 108 = 1
    16'b10000100_01101101 : OUT <= 1;  //132 / 109 = 1
    16'b10000100_01101110 : OUT <= 1;  //132 / 110 = 1
    16'b10000100_01101111 : OUT <= 1;  //132 / 111 = 1
    16'b10000100_01110000 : OUT <= 1;  //132 / 112 = 1
    16'b10000100_01110001 : OUT <= 1;  //132 / 113 = 1
    16'b10000100_01110010 : OUT <= 1;  //132 / 114 = 1
    16'b10000100_01110011 : OUT <= 1;  //132 / 115 = 1
    16'b10000100_01110100 : OUT <= 1;  //132 / 116 = 1
    16'b10000100_01110101 : OUT <= 1;  //132 / 117 = 1
    16'b10000100_01110110 : OUT <= 1;  //132 / 118 = 1
    16'b10000100_01110111 : OUT <= 1;  //132 / 119 = 1
    16'b10000100_01111000 : OUT <= 1;  //132 / 120 = 1
    16'b10000100_01111001 : OUT <= 1;  //132 / 121 = 1
    16'b10000100_01111010 : OUT <= 1;  //132 / 122 = 1
    16'b10000100_01111011 : OUT <= 1;  //132 / 123 = 1
    16'b10000100_01111100 : OUT <= 1;  //132 / 124 = 1
    16'b10000100_01111101 : OUT <= 1;  //132 / 125 = 1
    16'b10000100_01111110 : OUT <= 1;  //132 / 126 = 1
    16'b10000100_01111111 : OUT <= 1;  //132 / 127 = 1
    16'b10000100_10000000 : OUT <= 1;  //132 / 128 = 1
    16'b10000100_10000001 : OUT <= 1;  //132 / 129 = 1
    16'b10000100_10000010 : OUT <= 1;  //132 / 130 = 1
    16'b10000100_10000011 : OUT <= 1;  //132 / 131 = 1
    16'b10000100_10000100 : OUT <= 1;  //132 / 132 = 1
    16'b10000100_10000101 : OUT <= 0;  //132 / 133 = 0
    16'b10000100_10000110 : OUT <= 0;  //132 / 134 = 0
    16'b10000100_10000111 : OUT <= 0;  //132 / 135 = 0
    16'b10000100_10001000 : OUT <= 0;  //132 / 136 = 0
    16'b10000100_10001001 : OUT <= 0;  //132 / 137 = 0
    16'b10000100_10001010 : OUT <= 0;  //132 / 138 = 0
    16'b10000100_10001011 : OUT <= 0;  //132 / 139 = 0
    16'b10000100_10001100 : OUT <= 0;  //132 / 140 = 0
    16'b10000100_10001101 : OUT <= 0;  //132 / 141 = 0
    16'b10000100_10001110 : OUT <= 0;  //132 / 142 = 0
    16'b10000100_10001111 : OUT <= 0;  //132 / 143 = 0
    16'b10000100_10010000 : OUT <= 0;  //132 / 144 = 0
    16'b10000100_10010001 : OUT <= 0;  //132 / 145 = 0
    16'b10000100_10010010 : OUT <= 0;  //132 / 146 = 0
    16'b10000100_10010011 : OUT <= 0;  //132 / 147 = 0
    16'b10000100_10010100 : OUT <= 0;  //132 / 148 = 0
    16'b10000100_10010101 : OUT <= 0;  //132 / 149 = 0
    16'b10000100_10010110 : OUT <= 0;  //132 / 150 = 0
    16'b10000100_10010111 : OUT <= 0;  //132 / 151 = 0
    16'b10000100_10011000 : OUT <= 0;  //132 / 152 = 0
    16'b10000100_10011001 : OUT <= 0;  //132 / 153 = 0
    16'b10000100_10011010 : OUT <= 0;  //132 / 154 = 0
    16'b10000100_10011011 : OUT <= 0;  //132 / 155 = 0
    16'b10000100_10011100 : OUT <= 0;  //132 / 156 = 0
    16'b10000100_10011101 : OUT <= 0;  //132 / 157 = 0
    16'b10000100_10011110 : OUT <= 0;  //132 / 158 = 0
    16'b10000100_10011111 : OUT <= 0;  //132 / 159 = 0
    16'b10000100_10100000 : OUT <= 0;  //132 / 160 = 0
    16'b10000100_10100001 : OUT <= 0;  //132 / 161 = 0
    16'b10000100_10100010 : OUT <= 0;  //132 / 162 = 0
    16'b10000100_10100011 : OUT <= 0;  //132 / 163 = 0
    16'b10000100_10100100 : OUT <= 0;  //132 / 164 = 0
    16'b10000100_10100101 : OUT <= 0;  //132 / 165 = 0
    16'b10000100_10100110 : OUT <= 0;  //132 / 166 = 0
    16'b10000100_10100111 : OUT <= 0;  //132 / 167 = 0
    16'b10000100_10101000 : OUT <= 0;  //132 / 168 = 0
    16'b10000100_10101001 : OUT <= 0;  //132 / 169 = 0
    16'b10000100_10101010 : OUT <= 0;  //132 / 170 = 0
    16'b10000100_10101011 : OUT <= 0;  //132 / 171 = 0
    16'b10000100_10101100 : OUT <= 0;  //132 / 172 = 0
    16'b10000100_10101101 : OUT <= 0;  //132 / 173 = 0
    16'b10000100_10101110 : OUT <= 0;  //132 / 174 = 0
    16'b10000100_10101111 : OUT <= 0;  //132 / 175 = 0
    16'b10000100_10110000 : OUT <= 0;  //132 / 176 = 0
    16'b10000100_10110001 : OUT <= 0;  //132 / 177 = 0
    16'b10000100_10110010 : OUT <= 0;  //132 / 178 = 0
    16'b10000100_10110011 : OUT <= 0;  //132 / 179 = 0
    16'b10000100_10110100 : OUT <= 0;  //132 / 180 = 0
    16'b10000100_10110101 : OUT <= 0;  //132 / 181 = 0
    16'b10000100_10110110 : OUT <= 0;  //132 / 182 = 0
    16'b10000100_10110111 : OUT <= 0;  //132 / 183 = 0
    16'b10000100_10111000 : OUT <= 0;  //132 / 184 = 0
    16'b10000100_10111001 : OUT <= 0;  //132 / 185 = 0
    16'b10000100_10111010 : OUT <= 0;  //132 / 186 = 0
    16'b10000100_10111011 : OUT <= 0;  //132 / 187 = 0
    16'b10000100_10111100 : OUT <= 0;  //132 / 188 = 0
    16'b10000100_10111101 : OUT <= 0;  //132 / 189 = 0
    16'b10000100_10111110 : OUT <= 0;  //132 / 190 = 0
    16'b10000100_10111111 : OUT <= 0;  //132 / 191 = 0
    16'b10000100_11000000 : OUT <= 0;  //132 / 192 = 0
    16'b10000100_11000001 : OUT <= 0;  //132 / 193 = 0
    16'b10000100_11000010 : OUT <= 0;  //132 / 194 = 0
    16'b10000100_11000011 : OUT <= 0;  //132 / 195 = 0
    16'b10000100_11000100 : OUT <= 0;  //132 / 196 = 0
    16'b10000100_11000101 : OUT <= 0;  //132 / 197 = 0
    16'b10000100_11000110 : OUT <= 0;  //132 / 198 = 0
    16'b10000100_11000111 : OUT <= 0;  //132 / 199 = 0
    16'b10000100_11001000 : OUT <= 0;  //132 / 200 = 0
    16'b10000100_11001001 : OUT <= 0;  //132 / 201 = 0
    16'b10000100_11001010 : OUT <= 0;  //132 / 202 = 0
    16'b10000100_11001011 : OUT <= 0;  //132 / 203 = 0
    16'b10000100_11001100 : OUT <= 0;  //132 / 204 = 0
    16'b10000100_11001101 : OUT <= 0;  //132 / 205 = 0
    16'b10000100_11001110 : OUT <= 0;  //132 / 206 = 0
    16'b10000100_11001111 : OUT <= 0;  //132 / 207 = 0
    16'b10000100_11010000 : OUT <= 0;  //132 / 208 = 0
    16'b10000100_11010001 : OUT <= 0;  //132 / 209 = 0
    16'b10000100_11010010 : OUT <= 0;  //132 / 210 = 0
    16'b10000100_11010011 : OUT <= 0;  //132 / 211 = 0
    16'b10000100_11010100 : OUT <= 0;  //132 / 212 = 0
    16'b10000100_11010101 : OUT <= 0;  //132 / 213 = 0
    16'b10000100_11010110 : OUT <= 0;  //132 / 214 = 0
    16'b10000100_11010111 : OUT <= 0;  //132 / 215 = 0
    16'b10000100_11011000 : OUT <= 0;  //132 / 216 = 0
    16'b10000100_11011001 : OUT <= 0;  //132 / 217 = 0
    16'b10000100_11011010 : OUT <= 0;  //132 / 218 = 0
    16'b10000100_11011011 : OUT <= 0;  //132 / 219 = 0
    16'b10000100_11011100 : OUT <= 0;  //132 / 220 = 0
    16'b10000100_11011101 : OUT <= 0;  //132 / 221 = 0
    16'b10000100_11011110 : OUT <= 0;  //132 / 222 = 0
    16'b10000100_11011111 : OUT <= 0;  //132 / 223 = 0
    16'b10000100_11100000 : OUT <= 0;  //132 / 224 = 0
    16'b10000100_11100001 : OUT <= 0;  //132 / 225 = 0
    16'b10000100_11100010 : OUT <= 0;  //132 / 226 = 0
    16'b10000100_11100011 : OUT <= 0;  //132 / 227 = 0
    16'b10000100_11100100 : OUT <= 0;  //132 / 228 = 0
    16'b10000100_11100101 : OUT <= 0;  //132 / 229 = 0
    16'b10000100_11100110 : OUT <= 0;  //132 / 230 = 0
    16'b10000100_11100111 : OUT <= 0;  //132 / 231 = 0
    16'b10000100_11101000 : OUT <= 0;  //132 / 232 = 0
    16'b10000100_11101001 : OUT <= 0;  //132 / 233 = 0
    16'b10000100_11101010 : OUT <= 0;  //132 / 234 = 0
    16'b10000100_11101011 : OUT <= 0;  //132 / 235 = 0
    16'b10000100_11101100 : OUT <= 0;  //132 / 236 = 0
    16'b10000100_11101101 : OUT <= 0;  //132 / 237 = 0
    16'b10000100_11101110 : OUT <= 0;  //132 / 238 = 0
    16'b10000100_11101111 : OUT <= 0;  //132 / 239 = 0
    16'b10000100_11110000 : OUT <= 0;  //132 / 240 = 0
    16'b10000100_11110001 : OUT <= 0;  //132 / 241 = 0
    16'b10000100_11110010 : OUT <= 0;  //132 / 242 = 0
    16'b10000100_11110011 : OUT <= 0;  //132 / 243 = 0
    16'b10000100_11110100 : OUT <= 0;  //132 / 244 = 0
    16'b10000100_11110101 : OUT <= 0;  //132 / 245 = 0
    16'b10000100_11110110 : OUT <= 0;  //132 / 246 = 0
    16'b10000100_11110111 : OUT <= 0;  //132 / 247 = 0
    16'b10000100_11111000 : OUT <= 0;  //132 / 248 = 0
    16'b10000100_11111001 : OUT <= 0;  //132 / 249 = 0
    16'b10000100_11111010 : OUT <= 0;  //132 / 250 = 0
    16'b10000100_11111011 : OUT <= 0;  //132 / 251 = 0
    16'b10000100_11111100 : OUT <= 0;  //132 / 252 = 0
    16'b10000100_11111101 : OUT <= 0;  //132 / 253 = 0
    16'b10000100_11111110 : OUT <= 0;  //132 / 254 = 0
    16'b10000100_11111111 : OUT <= 0;  //132 / 255 = 0
    16'b10000101_00000000 : OUT <= 0;  //133 / 0 = 0
    16'b10000101_00000001 : OUT <= 133;  //133 / 1 = 133
    16'b10000101_00000010 : OUT <= 66;  //133 / 2 = 66
    16'b10000101_00000011 : OUT <= 44;  //133 / 3 = 44
    16'b10000101_00000100 : OUT <= 33;  //133 / 4 = 33
    16'b10000101_00000101 : OUT <= 26;  //133 / 5 = 26
    16'b10000101_00000110 : OUT <= 22;  //133 / 6 = 22
    16'b10000101_00000111 : OUT <= 19;  //133 / 7 = 19
    16'b10000101_00001000 : OUT <= 16;  //133 / 8 = 16
    16'b10000101_00001001 : OUT <= 14;  //133 / 9 = 14
    16'b10000101_00001010 : OUT <= 13;  //133 / 10 = 13
    16'b10000101_00001011 : OUT <= 12;  //133 / 11 = 12
    16'b10000101_00001100 : OUT <= 11;  //133 / 12 = 11
    16'b10000101_00001101 : OUT <= 10;  //133 / 13 = 10
    16'b10000101_00001110 : OUT <= 9;  //133 / 14 = 9
    16'b10000101_00001111 : OUT <= 8;  //133 / 15 = 8
    16'b10000101_00010000 : OUT <= 8;  //133 / 16 = 8
    16'b10000101_00010001 : OUT <= 7;  //133 / 17 = 7
    16'b10000101_00010010 : OUT <= 7;  //133 / 18 = 7
    16'b10000101_00010011 : OUT <= 7;  //133 / 19 = 7
    16'b10000101_00010100 : OUT <= 6;  //133 / 20 = 6
    16'b10000101_00010101 : OUT <= 6;  //133 / 21 = 6
    16'b10000101_00010110 : OUT <= 6;  //133 / 22 = 6
    16'b10000101_00010111 : OUT <= 5;  //133 / 23 = 5
    16'b10000101_00011000 : OUT <= 5;  //133 / 24 = 5
    16'b10000101_00011001 : OUT <= 5;  //133 / 25 = 5
    16'b10000101_00011010 : OUT <= 5;  //133 / 26 = 5
    16'b10000101_00011011 : OUT <= 4;  //133 / 27 = 4
    16'b10000101_00011100 : OUT <= 4;  //133 / 28 = 4
    16'b10000101_00011101 : OUT <= 4;  //133 / 29 = 4
    16'b10000101_00011110 : OUT <= 4;  //133 / 30 = 4
    16'b10000101_00011111 : OUT <= 4;  //133 / 31 = 4
    16'b10000101_00100000 : OUT <= 4;  //133 / 32 = 4
    16'b10000101_00100001 : OUT <= 4;  //133 / 33 = 4
    16'b10000101_00100010 : OUT <= 3;  //133 / 34 = 3
    16'b10000101_00100011 : OUT <= 3;  //133 / 35 = 3
    16'b10000101_00100100 : OUT <= 3;  //133 / 36 = 3
    16'b10000101_00100101 : OUT <= 3;  //133 / 37 = 3
    16'b10000101_00100110 : OUT <= 3;  //133 / 38 = 3
    16'b10000101_00100111 : OUT <= 3;  //133 / 39 = 3
    16'b10000101_00101000 : OUT <= 3;  //133 / 40 = 3
    16'b10000101_00101001 : OUT <= 3;  //133 / 41 = 3
    16'b10000101_00101010 : OUT <= 3;  //133 / 42 = 3
    16'b10000101_00101011 : OUT <= 3;  //133 / 43 = 3
    16'b10000101_00101100 : OUT <= 3;  //133 / 44 = 3
    16'b10000101_00101101 : OUT <= 2;  //133 / 45 = 2
    16'b10000101_00101110 : OUT <= 2;  //133 / 46 = 2
    16'b10000101_00101111 : OUT <= 2;  //133 / 47 = 2
    16'b10000101_00110000 : OUT <= 2;  //133 / 48 = 2
    16'b10000101_00110001 : OUT <= 2;  //133 / 49 = 2
    16'b10000101_00110010 : OUT <= 2;  //133 / 50 = 2
    16'b10000101_00110011 : OUT <= 2;  //133 / 51 = 2
    16'b10000101_00110100 : OUT <= 2;  //133 / 52 = 2
    16'b10000101_00110101 : OUT <= 2;  //133 / 53 = 2
    16'b10000101_00110110 : OUT <= 2;  //133 / 54 = 2
    16'b10000101_00110111 : OUT <= 2;  //133 / 55 = 2
    16'b10000101_00111000 : OUT <= 2;  //133 / 56 = 2
    16'b10000101_00111001 : OUT <= 2;  //133 / 57 = 2
    16'b10000101_00111010 : OUT <= 2;  //133 / 58 = 2
    16'b10000101_00111011 : OUT <= 2;  //133 / 59 = 2
    16'b10000101_00111100 : OUT <= 2;  //133 / 60 = 2
    16'b10000101_00111101 : OUT <= 2;  //133 / 61 = 2
    16'b10000101_00111110 : OUT <= 2;  //133 / 62 = 2
    16'b10000101_00111111 : OUT <= 2;  //133 / 63 = 2
    16'b10000101_01000000 : OUT <= 2;  //133 / 64 = 2
    16'b10000101_01000001 : OUT <= 2;  //133 / 65 = 2
    16'b10000101_01000010 : OUT <= 2;  //133 / 66 = 2
    16'b10000101_01000011 : OUT <= 1;  //133 / 67 = 1
    16'b10000101_01000100 : OUT <= 1;  //133 / 68 = 1
    16'b10000101_01000101 : OUT <= 1;  //133 / 69 = 1
    16'b10000101_01000110 : OUT <= 1;  //133 / 70 = 1
    16'b10000101_01000111 : OUT <= 1;  //133 / 71 = 1
    16'b10000101_01001000 : OUT <= 1;  //133 / 72 = 1
    16'b10000101_01001001 : OUT <= 1;  //133 / 73 = 1
    16'b10000101_01001010 : OUT <= 1;  //133 / 74 = 1
    16'b10000101_01001011 : OUT <= 1;  //133 / 75 = 1
    16'b10000101_01001100 : OUT <= 1;  //133 / 76 = 1
    16'b10000101_01001101 : OUT <= 1;  //133 / 77 = 1
    16'b10000101_01001110 : OUT <= 1;  //133 / 78 = 1
    16'b10000101_01001111 : OUT <= 1;  //133 / 79 = 1
    16'b10000101_01010000 : OUT <= 1;  //133 / 80 = 1
    16'b10000101_01010001 : OUT <= 1;  //133 / 81 = 1
    16'b10000101_01010010 : OUT <= 1;  //133 / 82 = 1
    16'b10000101_01010011 : OUT <= 1;  //133 / 83 = 1
    16'b10000101_01010100 : OUT <= 1;  //133 / 84 = 1
    16'b10000101_01010101 : OUT <= 1;  //133 / 85 = 1
    16'b10000101_01010110 : OUT <= 1;  //133 / 86 = 1
    16'b10000101_01010111 : OUT <= 1;  //133 / 87 = 1
    16'b10000101_01011000 : OUT <= 1;  //133 / 88 = 1
    16'b10000101_01011001 : OUT <= 1;  //133 / 89 = 1
    16'b10000101_01011010 : OUT <= 1;  //133 / 90 = 1
    16'b10000101_01011011 : OUT <= 1;  //133 / 91 = 1
    16'b10000101_01011100 : OUT <= 1;  //133 / 92 = 1
    16'b10000101_01011101 : OUT <= 1;  //133 / 93 = 1
    16'b10000101_01011110 : OUT <= 1;  //133 / 94 = 1
    16'b10000101_01011111 : OUT <= 1;  //133 / 95 = 1
    16'b10000101_01100000 : OUT <= 1;  //133 / 96 = 1
    16'b10000101_01100001 : OUT <= 1;  //133 / 97 = 1
    16'b10000101_01100010 : OUT <= 1;  //133 / 98 = 1
    16'b10000101_01100011 : OUT <= 1;  //133 / 99 = 1
    16'b10000101_01100100 : OUT <= 1;  //133 / 100 = 1
    16'b10000101_01100101 : OUT <= 1;  //133 / 101 = 1
    16'b10000101_01100110 : OUT <= 1;  //133 / 102 = 1
    16'b10000101_01100111 : OUT <= 1;  //133 / 103 = 1
    16'b10000101_01101000 : OUT <= 1;  //133 / 104 = 1
    16'b10000101_01101001 : OUT <= 1;  //133 / 105 = 1
    16'b10000101_01101010 : OUT <= 1;  //133 / 106 = 1
    16'b10000101_01101011 : OUT <= 1;  //133 / 107 = 1
    16'b10000101_01101100 : OUT <= 1;  //133 / 108 = 1
    16'b10000101_01101101 : OUT <= 1;  //133 / 109 = 1
    16'b10000101_01101110 : OUT <= 1;  //133 / 110 = 1
    16'b10000101_01101111 : OUT <= 1;  //133 / 111 = 1
    16'b10000101_01110000 : OUT <= 1;  //133 / 112 = 1
    16'b10000101_01110001 : OUT <= 1;  //133 / 113 = 1
    16'b10000101_01110010 : OUT <= 1;  //133 / 114 = 1
    16'b10000101_01110011 : OUT <= 1;  //133 / 115 = 1
    16'b10000101_01110100 : OUT <= 1;  //133 / 116 = 1
    16'b10000101_01110101 : OUT <= 1;  //133 / 117 = 1
    16'b10000101_01110110 : OUT <= 1;  //133 / 118 = 1
    16'b10000101_01110111 : OUT <= 1;  //133 / 119 = 1
    16'b10000101_01111000 : OUT <= 1;  //133 / 120 = 1
    16'b10000101_01111001 : OUT <= 1;  //133 / 121 = 1
    16'b10000101_01111010 : OUT <= 1;  //133 / 122 = 1
    16'b10000101_01111011 : OUT <= 1;  //133 / 123 = 1
    16'b10000101_01111100 : OUT <= 1;  //133 / 124 = 1
    16'b10000101_01111101 : OUT <= 1;  //133 / 125 = 1
    16'b10000101_01111110 : OUT <= 1;  //133 / 126 = 1
    16'b10000101_01111111 : OUT <= 1;  //133 / 127 = 1
    16'b10000101_10000000 : OUT <= 1;  //133 / 128 = 1
    16'b10000101_10000001 : OUT <= 1;  //133 / 129 = 1
    16'b10000101_10000010 : OUT <= 1;  //133 / 130 = 1
    16'b10000101_10000011 : OUT <= 1;  //133 / 131 = 1
    16'b10000101_10000100 : OUT <= 1;  //133 / 132 = 1
    16'b10000101_10000101 : OUT <= 1;  //133 / 133 = 1
    16'b10000101_10000110 : OUT <= 0;  //133 / 134 = 0
    16'b10000101_10000111 : OUT <= 0;  //133 / 135 = 0
    16'b10000101_10001000 : OUT <= 0;  //133 / 136 = 0
    16'b10000101_10001001 : OUT <= 0;  //133 / 137 = 0
    16'b10000101_10001010 : OUT <= 0;  //133 / 138 = 0
    16'b10000101_10001011 : OUT <= 0;  //133 / 139 = 0
    16'b10000101_10001100 : OUT <= 0;  //133 / 140 = 0
    16'b10000101_10001101 : OUT <= 0;  //133 / 141 = 0
    16'b10000101_10001110 : OUT <= 0;  //133 / 142 = 0
    16'b10000101_10001111 : OUT <= 0;  //133 / 143 = 0
    16'b10000101_10010000 : OUT <= 0;  //133 / 144 = 0
    16'b10000101_10010001 : OUT <= 0;  //133 / 145 = 0
    16'b10000101_10010010 : OUT <= 0;  //133 / 146 = 0
    16'b10000101_10010011 : OUT <= 0;  //133 / 147 = 0
    16'b10000101_10010100 : OUT <= 0;  //133 / 148 = 0
    16'b10000101_10010101 : OUT <= 0;  //133 / 149 = 0
    16'b10000101_10010110 : OUT <= 0;  //133 / 150 = 0
    16'b10000101_10010111 : OUT <= 0;  //133 / 151 = 0
    16'b10000101_10011000 : OUT <= 0;  //133 / 152 = 0
    16'b10000101_10011001 : OUT <= 0;  //133 / 153 = 0
    16'b10000101_10011010 : OUT <= 0;  //133 / 154 = 0
    16'b10000101_10011011 : OUT <= 0;  //133 / 155 = 0
    16'b10000101_10011100 : OUT <= 0;  //133 / 156 = 0
    16'b10000101_10011101 : OUT <= 0;  //133 / 157 = 0
    16'b10000101_10011110 : OUT <= 0;  //133 / 158 = 0
    16'b10000101_10011111 : OUT <= 0;  //133 / 159 = 0
    16'b10000101_10100000 : OUT <= 0;  //133 / 160 = 0
    16'b10000101_10100001 : OUT <= 0;  //133 / 161 = 0
    16'b10000101_10100010 : OUT <= 0;  //133 / 162 = 0
    16'b10000101_10100011 : OUT <= 0;  //133 / 163 = 0
    16'b10000101_10100100 : OUT <= 0;  //133 / 164 = 0
    16'b10000101_10100101 : OUT <= 0;  //133 / 165 = 0
    16'b10000101_10100110 : OUT <= 0;  //133 / 166 = 0
    16'b10000101_10100111 : OUT <= 0;  //133 / 167 = 0
    16'b10000101_10101000 : OUT <= 0;  //133 / 168 = 0
    16'b10000101_10101001 : OUT <= 0;  //133 / 169 = 0
    16'b10000101_10101010 : OUT <= 0;  //133 / 170 = 0
    16'b10000101_10101011 : OUT <= 0;  //133 / 171 = 0
    16'b10000101_10101100 : OUT <= 0;  //133 / 172 = 0
    16'b10000101_10101101 : OUT <= 0;  //133 / 173 = 0
    16'b10000101_10101110 : OUT <= 0;  //133 / 174 = 0
    16'b10000101_10101111 : OUT <= 0;  //133 / 175 = 0
    16'b10000101_10110000 : OUT <= 0;  //133 / 176 = 0
    16'b10000101_10110001 : OUT <= 0;  //133 / 177 = 0
    16'b10000101_10110010 : OUT <= 0;  //133 / 178 = 0
    16'b10000101_10110011 : OUT <= 0;  //133 / 179 = 0
    16'b10000101_10110100 : OUT <= 0;  //133 / 180 = 0
    16'b10000101_10110101 : OUT <= 0;  //133 / 181 = 0
    16'b10000101_10110110 : OUT <= 0;  //133 / 182 = 0
    16'b10000101_10110111 : OUT <= 0;  //133 / 183 = 0
    16'b10000101_10111000 : OUT <= 0;  //133 / 184 = 0
    16'b10000101_10111001 : OUT <= 0;  //133 / 185 = 0
    16'b10000101_10111010 : OUT <= 0;  //133 / 186 = 0
    16'b10000101_10111011 : OUT <= 0;  //133 / 187 = 0
    16'b10000101_10111100 : OUT <= 0;  //133 / 188 = 0
    16'b10000101_10111101 : OUT <= 0;  //133 / 189 = 0
    16'b10000101_10111110 : OUT <= 0;  //133 / 190 = 0
    16'b10000101_10111111 : OUT <= 0;  //133 / 191 = 0
    16'b10000101_11000000 : OUT <= 0;  //133 / 192 = 0
    16'b10000101_11000001 : OUT <= 0;  //133 / 193 = 0
    16'b10000101_11000010 : OUT <= 0;  //133 / 194 = 0
    16'b10000101_11000011 : OUT <= 0;  //133 / 195 = 0
    16'b10000101_11000100 : OUT <= 0;  //133 / 196 = 0
    16'b10000101_11000101 : OUT <= 0;  //133 / 197 = 0
    16'b10000101_11000110 : OUT <= 0;  //133 / 198 = 0
    16'b10000101_11000111 : OUT <= 0;  //133 / 199 = 0
    16'b10000101_11001000 : OUT <= 0;  //133 / 200 = 0
    16'b10000101_11001001 : OUT <= 0;  //133 / 201 = 0
    16'b10000101_11001010 : OUT <= 0;  //133 / 202 = 0
    16'b10000101_11001011 : OUT <= 0;  //133 / 203 = 0
    16'b10000101_11001100 : OUT <= 0;  //133 / 204 = 0
    16'b10000101_11001101 : OUT <= 0;  //133 / 205 = 0
    16'b10000101_11001110 : OUT <= 0;  //133 / 206 = 0
    16'b10000101_11001111 : OUT <= 0;  //133 / 207 = 0
    16'b10000101_11010000 : OUT <= 0;  //133 / 208 = 0
    16'b10000101_11010001 : OUT <= 0;  //133 / 209 = 0
    16'b10000101_11010010 : OUT <= 0;  //133 / 210 = 0
    16'b10000101_11010011 : OUT <= 0;  //133 / 211 = 0
    16'b10000101_11010100 : OUT <= 0;  //133 / 212 = 0
    16'b10000101_11010101 : OUT <= 0;  //133 / 213 = 0
    16'b10000101_11010110 : OUT <= 0;  //133 / 214 = 0
    16'b10000101_11010111 : OUT <= 0;  //133 / 215 = 0
    16'b10000101_11011000 : OUT <= 0;  //133 / 216 = 0
    16'b10000101_11011001 : OUT <= 0;  //133 / 217 = 0
    16'b10000101_11011010 : OUT <= 0;  //133 / 218 = 0
    16'b10000101_11011011 : OUT <= 0;  //133 / 219 = 0
    16'b10000101_11011100 : OUT <= 0;  //133 / 220 = 0
    16'b10000101_11011101 : OUT <= 0;  //133 / 221 = 0
    16'b10000101_11011110 : OUT <= 0;  //133 / 222 = 0
    16'b10000101_11011111 : OUT <= 0;  //133 / 223 = 0
    16'b10000101_11100000 : OUT <= 0;  //133 / 224 = 0
    16'b10000101_11100001 : OUT <= 0;  //133 / 225 = 0
    16'b10000101_11100010 : OUT <= 0;  //133 / 226 = 0
    16'b10000101_11100011 : OUT <= 0;  //133 / 227 = 0
    16'b10000101_11100100 : OUT <= 0;  //133 / 228 = 0
    16'b10000101_11100101 : OUT <= 0;  //133 / 229 = 0
    16'b10000101_11100110 : OUT <= 0;  //133 / 230 = 0
    16'b10000101_11100111 : OUT <= 0;  //133 / 231 = 0
    16'b10000101_11101000 : OUT <= 0;  //133 / 232 = 0
    16'b10000101_11101001 : OUT <= 0;  //133 / 233 = 0
    16'b10000101_11101010 : OUT <= 0;  //133 / 234 = 0
    16'b10000101_11101011 : OUT <= 0;  //133 / 235 = 0
    16'b10000101_11101100 : OUT <= 0;  //133 / 236 = 0
    16'b10000101_11101101 : OUT <= 0;  //133 / 237 = 0
    16'b10000101_11101110 : OUT <= 0;  //133 / 238 = 0
    16'b10000101_11101111 : OUT <= 0;  //133 / 239 = 0
    16'b10000101_11110000 : OUT <= 0;  //133 / 240 = 0
    16'b10000101_11110001 : OUT <= 0;  //133 / 241 = 0
    16'b10000101_11110010 : OUT <= 0;  //133 / 242 = 0
    16'b10000101_11110011 : OUT <= 0;  //133 / 243 = 0
    16'b10000101_11110100 : OUT <= 0;  //133 / 244 = 0
    16'b10000101_11110101 : OUT <= 0;  //133 / 245 = 0
    16'b10000101_11110110 : OUT <= 0;  //133 / 246 = 0
    16'b10000101_11110111 : OUT <= 0;  //133 / 247 = 0
    16'b10000101_11111000 : OUT <= 0;  //133 / 248 = 0
    16'b10000101_11111001 : OUT <= 0;  //133 / 249 = 0
    16'b10000101_11111010 : OUT <= 0;  //133 / 250 = 0
    16'b10000101_11111011 : OUT <= 0;  //133 / 251 = 0
    16'b10000101_11111100 : OUT <= 0;  //133 / 252 = 0
    16'b10000101_11111101 : OUT <= 0;  //133 / 253 = 0
    16'b10000101_11111110 : OUT <= 0;  //133 / 254 = 0
    16'b10000101_11111111 : OUT <= 0;  //133 / 255 = 0
    16'b10000110_00000000 : OUT <= 0;  //134 / 0 = 0
    16'b10000110_00000001 : OUT <= 134;  //134 / 1 = 134
    16'b10000110_00000010 : OUT <= 67;  //134 / 2 = 67
    16'b10000110_00000011 : OUT <= 44;  //134 / 3 = 44
    16'b10000110_00000100 : OUT <= 33;  //134 / 4 = 33
    16'b10000110_00000101 : OUT <= 26;  //134 / 5 = 26
    16'b10000110_00000110 : OUT <= 22;  //134 / 6 = 22
    16'b10000110_00000111 : OUT <= 19;  //134 / 7 = 19
    16'b10000110_00001000 : OUT <= 16;  //134 / 8 = 16
    16'b10000110_00001001 : OUT <= 14;  //134 / 9 = 14
    16'b10000110_00001010 : OUT <= 13;  //134 / 10 = 13
    16'b10000110_00001011 : OUT <= 12;  //134 / 11 = 12
    16'b10000110_00001100 : OUT <= 11;  //134 / 12 = 11
    16'b10000110_00001101 : OUT <= 10;  //134 / 13 = 10
    16'b10000110_00001110 : OUT <= 9;  //134 / 14 = 9
    16'b10000110_00001111 : OUT <= 8;  //134 / 15 = 8
    16'b10000110_00010000 : OUT <= 8;  //134 / 16 = 8
    16'b10000110_00010001 : OUT <= 7;  //134 / 17 = 7
    16'b10000110_00010010 : OUT <= 7;  //134 / 18 = 7
    16'b10000110_00010011 : OUT <= 7;  //134 / 19 = 7
    16'b10000110_00010100 : OUT <= 6;  //134 / 20 = 6
    16'b10000110_00010101 : OUT <= 6;  //134 / 21 = 6
    16'b10000110_00010110 : OUT <= 6;  //134 / 22 = 6
    16'b10000110_00010111 : OUT <= 5;  //134 / 23 = 5
    16'b10000110_00011000 : OUT <= 5;  //134 / 24 = 5
    16'b10000110_00011001 : OUT <= 5;  //134 / 25 = 5
    16'b10000110_00011010 : OUT <= 5;  //134 / 26 = 5
    16'b10000110_00011011 : OUT <= 4;  //134 / 27 = 4
    16'b10000110_00011100 : OUT <= 4;  //134 / 28 = 4
    16'b10000110_00011101 : OUT <= 4;  //134 / 29 = 4
    16'b10000110_00011110 : OUT <= 4;  //134 / 30 = 4
    16'b10000110_00011111 : OUT <= 4;  //134 / 31 = 4
    16'b10000110_00100000 : OUT <= 4;  //134 / 32 = 4
    16'b10000110_00100001 : OUT <= 4;  //134 / 33 = 4
    16'b10000110_00100010 : OUT <= 3;  //134 / 34 = 3
    16'b10000110_00100011 : OUT <= 3;  //134 / 35 = 3
    16'b10000110_00100100 : OUT <= 3;  //134 / 36 = 3
    16'b10000110_00100101 : OUT <= 3;  //134 / 37 = 3
    16'b10000110_00100110 : OUT <= 3;  //134 / 38 = 3
    16'b10000110_00100111 : OUT <= 3;  //134 / 39 = 3
    16'b10000110_00101000 : OUT <= 3;  //134 / 40 = 3
    16'b10000110_00101001 : OUT <= 3;  //134 / 41 = 3
    16'b10000110_00101010 : OUT <= 3;  //134 / 42 = 3
    16'b10000110_00101011 : OUT <= 3;  //134 / 43 = 3
    16'b10000110_00101100 : OUT <= 3;  //134 / 44 = 3
    16'b10000110_00101101 : OUT <= 2;  //134 / 45 = 2
    16'b10000110_00101110 : OUT <= 2;  //134 / 46 = 2
    16'b10000110_00101111 : OUT <= 2;  //134 / 47 = 2
    16'b10000110_00110000 : OUT <= 2;  //134 / 48 = 2
    16'b10000110_00110001 : OUT <= 2;  //134 / 49 = 2
    16'b10000110_00110010 : OUT <= 2;  //134 / 50 = 2
    16'b10000110_00110011 : OUT <= 2;  //134 / 51 = 2
    16'b10000110_00110100 : OUT <= 2;  //134 / 52 = 2
    16'b10000110_00110101 : OUT <= 2;  //134 / 53 = 2
    16'b10000110_00110110 : OUT <= 2;  //134 / 54 = 2
    16'b10000110_00110111 : OUT <= 2;  //134 / 55 = 2
    16'b10000110_00111000 : OUT <= 2;  //134 / 56 = 2
    16'b10000110_00111001 : OUT <= 2;  //134 / 57 = 2
    16'b10000110_00111010 : OUT <= 2;  //134 / 58 = 2
    16'b10000110_00111011 : OUT <= 2;  //134 / 59 = 2
    16'b10000110_00111100 : OUT <= 2;  //134 / 60 = 2
    16'b10000110_00111101 : OUT <= 2;  //134 / 61 = 2
    16'b10000110_00111110 : OUT <= 2;  //134 / 62 = 2
    16'b10000110_00111111 : OUT <= 2;  //134 / 63 = 2
    16'b10000110_01000000 : OUT <= 2;  //134 / 64 = 2
    16'b10000110_01000001 : OUT <= 2;  //134 / 65 = 2
    16'b10000110_01000010 : OUT <= 2;  //134 / 66 = 2
    16'b10000110_01000011 : OUT <= 2;  //134 / 67 = 2
    16'b10000110_01000100 : OUT <= 1;  //134 / 68 = 1
    16'b10000110_01000101 : OUT <= 1;  //134 / 69 = 1
    16'b10000110_01000110 : OUT <= 1;  //134 / 70 = 1
    16'b10000110_01000111 : OUT <= 1;  //134 / 71 = 1
    16'b10000110_01001000 : OUT <= 1;  //134 / 72 = 1
    16'b10000110_01001001 : OUT <= 1;  //134 / 73 = 1
    16'b10000110_01001010 : OUT <= 1;  //134 / 74 = 1
    16'b10000110_01001011 : OUT <= 1;  //134 / 75 = 1
    16'b10000110_01001100 : OUT <= 1;  //134 / 76 = 1
    16'b10000110_01001101 : OUT <= 1;  //134 / 77 = 1
    16'b10000110_01001110 : OUT <= 1;  //134 / 78 = 1
    16'b10000110_01001111 : OUT <= 1;  //134 / 79 = 1
    16'b10000110_01010000 : OUT <= 1;  //134 / 80 = 1
    16'b10000110_01010001 : OUT <= 1;  //134 / 81 = 1
    16'b10000110_01010010 : OUT <= 1;  //134 / 82 = 1
    16'b10000110_01010011 : OUT <= 1;  //134 / 83 = 1
    16'b10000110_01010100 : OUT <= 1;  //134 / 84 = 1
    16'b10000110_01010101 : OUT <= 1;  //134 / 85 = 1
    16'b10000110_01010110 : OUT <= 1;  //134 / 86 = 1
    16'b10000110_01010111 : OUT <= 1;  //134 / 87 = 1
    16'b10000110_01011000 : OUT <= 1;  //134 / 88 = 1
    16'b10000110_01011001 : OUT <= 1;  //134 / 89 = 1
    16'b10000110_01011010 : OUT <= 1;  //134 / 90 = 1
    16'b10000110_01011011 : OUT <= 1;  //134 / 91 = 1
    16'b10000110_01011100 : OUT <= 1;  //134 / 92 = 1
    16'b10000110_01011101 : OUT <= 1;  //134 / 93 = 1
    16'b10000110_01011110 : OUT <= 1;  //134 / 94 = 1
    16'b10000110_01011111 : OUT <= 1;  //134 / 95 = 1
    16'b10000110_01100000 : OUT <= 1;  //134 / 96 = 1
    16'b10000110_01100001 : OUT <= 1;  //134 / 97 = 1
    16'b10000110_01100010 : OUT <= 1;  //134 / 98 = 1
    16'b10000110_01100011 : OUT <= 1;  //134 / 99 = 1
    16'b10000110_01100100 : OUT <= 1;  //134 / 100 = 1
    16'b10000110_01100101 : OUT <= 1;  //134 / 101 = 1
    16'b10000110_01100110 : OUT <= 1;  //134 / 102 = 1
    16'b10000110_01100111 : OUT <= 1;  //134 / 103 = 1
    16'b10000110_01101000 : OUT <= 1;  //134 / 104 = 1
    16'b10000110_01101001 : OUT <= 1;  //134 / 105 = 1
    16'b10000110_01101010 : OUT <= 1;  //134 / 106 = 1
    16'b10000110_01101011 : OUT <= 1;  //134 / 107 = 1
    16'b10000110_01101100 : OUT <= 1;  //134 / 108 = 1
    16'b10000110_01101101 : OUT <= 1;  //134 / 109 = 1
    16'b10000110_01101110 : OUT <= 1;  //134 / 110 = 1
    16'b10000110_01101111 : OUT <= 1;  //134 / 111 = 1
    16'b10000110_01110000 : OUT <= 1;  //134 / 112 = 1
    16'b10000110_01110001 : OUT <= 1;  //134 / 113 = 1
    16'b10000110_01110010 : OUT <= 1;  //134 / 114 = 1
    16'b10000110_01110011 : OUT <= 1;  //134 / 115 = 1
    16'b10000110_01110100 : OUT <= 1;  //134 / 116 = 1
    16'b10000110_01110101 : OUT <= 1;  //134 / 117 = 1
    16'b10000110_01110110 : OUT <= 1;  //134 / 118 = 1
    16'b10000110_01110111 : OUT <= 1;  //134 / 119 = 1
    16'b10000110_01111000 : OUT <= 1;  //134 / 120 = 1
    16'b10000110_01111001 : OUT <= 1;  //134 / 121 = 1
    16'b10000110_01111010 : OUT <= 1;  //134 / 122 = 1
    16'b10000110_01111011 : OUT <= 1;  //134 / 123 = 1
    16'b10000110_01111100 : OUT <= 1;  //134 / 124 = 1
    16'b10000110_01111101 : OUT <= 1;  //134 / 125 = 1
    16'b10000110_01111110 : OUT <= 1;  //134 / 126 = 1
    16'b10000110_01111111 : OUT <= 1;  //134 / 127 = 1
    16'b10000110_10000000 : OUT <= 1;  //134 / 128 = 1
    16'b10000110_10000001 : OUT <= 1;  //134 / 129 = 1
    16'b10000110_10000010 : OUT <= 1;  //134 / 130 = 1
    16'b10000110_10000011 : OUT <= 1;  //134 / 131 = 1
    16'b10000110_10000100 : OUT <= 1;  //134 / 132 = 1
    16'b10000110_10000101 : OUT <= 1;  //134 / 133 = 1
    16'b10000110_10000110 : OUT <= 1;  //134 / 134 = 1
    16'b10000110_10000111 : OUT <= 0;  //134 / 135 = 0
    16'b10000110_10001000 : OUT <= 0;  //134 / 136 = 0
    16'b10000110_10001001 : OUT <= 0;  //134 / 137 = 0
    16'b10000110_10001010 : OUT <= 0;  //134 / 138 = 0
    16'b10000110_10001011 : OUT <= 0;  //134 / 139 = 0
    16'b10000110_10001100 : OUT <= 0;  //134 / 140 = 0
    16'b10000110_10001101 : OUT <= 0;  //134 / 141 = 0
    16'b10000110_10001110 : OUT <= 0;  //134 / 142 = 0
    16'b10000110_10001111 : OUT <= 0;  //134 / 143 = 0
    16'b10000110_10010000 : OUT <= 0;  //134 / 144 = 0
    16'b10000110_10010001 : OUT <= 0;  //134 / 145 = 0
    16'b10000110_10010010 : OUT <= 0;  //134 / 146 = 0
    16'b10000110_10010011 : OUT <= 0;  //134 / 147 = 0
    16'b10000110_10010100 : OUT <= 0;  //134 / 148 = 0
    16'b10000110_10010101 : OUT <= 0;  //134 / 149 = 0
    16'b10000110_10010110 : OUT <= 0;  //134 / 150 = 0
    16'b10000110_10010111 : OUT <= 0;  //134 / 151 = 0
    16'b10000110_10011000 : OUT <= 0;  //134 / 152 = 0
    16'b10000110_10011001 : OUT <= 0;  //134 / 153 = 0
    16'b10000110_10011010 : OUT <= 0;  //134 / 154 = 0
    16'b10000110_10011011 : OUT <= 0;  //134 / 155 = 0
    16'b10000110_10011100 : OUT <= 0;  //134 / 156 = 0
    16'b10000110_10011101 : OUT <= 0;  //134 / 157 = 0
    16'b10000110_10011110 : OUT <= 0;  //134 / 158 = 0
    16'b10000110_10011111 : OUT <= 0;  //134 / 159 = 0
    16'b10000110_10100000 : OUT <= 0;  //134 / 160 = 0
    16'b10000110_10100001 : OUT <= 0;  //134 / 161 = 0
    16'b10000110_10100010 : OUT <= 0;  //134 / 162 = 0
    16'b10000110_10100011 : OUT <= 0;  //134 / 163 = 0
    16'b10000110_10100100 : OUT <= 0;  //134 / 164 = 0
    16'b10000110_10100101 : OUT <= 0;  //134 / 165 = 0
    16'b10000110_10100110 : OUT <= 0;  //134 / 166 = 0
    16'b10000110_10100111 : OUT <= 0;  //134 / 167 = 0
    16'b10000110_10101000 : OUT <= 0;  //134 / 168 = 0
    16'b10000110_10101001 : OUT <= 0;  //134 / 169 = 0
    16'b10000110_10101010 : OUT <= 0;  //134 / 170 = 0
    16'b10000110_10101011 : OUT <= 0;  //134 / 171 = 0
    16'b10000110_10101100 : OUT <= 0;  //134 / 172 = 0
    16'b10000110_10101101 : OUT <= 0;  //134 / 173 = 0
    16'b10000110_10101110 : OUT <= 0;  //134 / 174 = 0
    16'b10000110_10101111 : OUT <= 0;  //134 / 175 = 0
    16'b10000110_10110000 : OUT <= 0;  //134 / 176 = 0
    16'b10000110_10110001 : OUT <= 0;  //134 / 177 = 0
    16'b10000110_10110010 : OUT <= 0;  //134 / 178 = 0
    16'b10000110_10110011 : OUT <= 0;  //134 / 179 = 0
    16'b10000110_10110100 : OUT <= 0;  //134 / 180 = 0
    16'b10000110_10110101 : OUT <= 0;  //134 / 181 = 0
    16'b10000110_10110110 : OUT <= 0;  //134 / 182 = 0
    16'b10000110_10110111 : OUT <= 0;  //134 / 183 = 0
    16'b10000110_10111000 : OUT <= 0;  //134 / 184 = 0
    16'b10000110_10111001 : OUT <= 0;  //134 / 185 = 0
    16'b10000110_10111010 : OUT <= 0;  //134 / 186 = 0
    16'b10000110_10111011 : OUT <= 0;  //134 / 187 = 0
    16'b10000110_10111100 : OUT <= 0;  //134 / 188 = 0
    16'b10000110_10111101 : OUT <= 0;  //134 / 189 = 0
    16'b10000110_10111110 : OUT <= 0;  //134 / 190 = 0
    16'b10000110_10111111 : OUT <= 0;  //134 / 191 = 0
    16'b10000110_11000000 : OUT <= 0;  //134 / 192 = 0
    16'b10000110_11000001 : OUT <= 0;  //134 / 193 = 0
    16'b10000110_11000010 : OUT <= 0;  //134 / 194 = 0
    16'b10000110_11000011 : OUT <= 0;  //134 / 195 = 0
    16'b10000110_11000100 : OUT <= 0;  //134 / 196 = 0
    16'b10000110_11000101 : OUT <= 0;  //134 / 197 = 0
    16'b10000110_11000110 : OUT <= 0;  //134 / 198 = 0
    16'b10000110_11000111 : OUT <= 0;  //134 / 199 = 0
    16'b10000110_11001000 : OUT <= 0;  //134 / 200 = 0
    16'b10000110_11001001 : OUT <= 0;  //134 / 201 = 0
    16'b10000110_11001010 : OUT <= 0;  //134 / 202 = 0
    16'b10000110_11001011 : OUT <= 0;  //134 / 203 = 0
    16'b10000110_11001100 : OUT <= 0;  //134 / 204 = 0
    16'b10000110_11001101 : OUT <= 0;  //134 / 205 = 0
    16'b10000110_11001110 : OUT <= 0;  //134 / 206 = 0
    16'b10000110_11001111 : OUT <= 0;  //134 / 207 = 0
    16'b10000110_11010000 : OUT <= 0;  //134 / 208 = 0
    16'b10000110_11010001 : OUT <= 0;  //134 / 209 = 0
    16'b10000110_11010010 : OUT <= 0;  //134 / 210 = 0
    16'b10000110_11010011 : OUT <= 0;  //134 / 211 = 0
    16'b10000110_11010100 : OUT <= 0;  //134 / 212 = 0
    16'b10000110_11010101 : OUT <= 0;  //134 / 213 = 0
    16'b10000110_11010110 : OUT <= 0;  //134 / 214 = 0
    16'b10000110_11010111 : OUT <= 0;  //134 / 215 = 0
    16'b10000110_11011000 : OUT <= 0;  //134 / 216 = 0
    16'b10000110_11011001 : OUT <= 0;  //134 / 217 = 0
    16'b10000110_11011010 : OUT <= 0;  //134 / 218 = 0
    16'b10000110_11011011 : OUT <= 0;  //134 / 219 = 0
    16'b10000110_11011100 : OUT <= 0;  //134 / 220 = 0
    16'b10000110_11011101 : OUT <= 0;  //134 / 221 = 0
    16'b10000110_11011110 : OUT <= 0;  //134 / 222 = 0
    16'b10000110_11011111 : OUT <= 0;  //134 / 223 = 0
    16'b10000110_11100000 : OUT <= 0;  //134 / 224 = 0
    16'b10000110_11100001 : OUT <= 0;  //134 / 225 = 0
    16'b10000110_11100010 : OUT <= 0;  //134 / 226 = 0
    16'b10000110_11100011 : OUT <= 0;  //134 / 227 = 0
    16'b10000110_11100100 : OUT <= 0;  //134 / 228 = 0
    16'b10000110_11100101 : OUT <= 0;  //134 / 229 = 0
    16'b10000110_11100110 : OUT <= 0;  //134 / 230 = 0
    16'b10000110_11100111 : OUT <= 0;  //134 / 231 = 0
    16'b10000110_11101000 : OUT <= 0;  //134 / 232 = 0
    16'b10000110_11101001 : OUT <= 0;  //134 / 233 = 0
    16'b10000110_11101010 : OUT <= 0;  //134 / 234 = 0
    16'b10000110_11101011 : OUT <= 0;  //134 / 235 = 0
    16'b10000110_11101100 : OUT <= 0;  //134 / 236 = 0
    16'b10000110_11101101 : OUT <= 0;  //134 / 237 = 0
    16'b10000110_11101110 : OUT <= 0;  //134 / 238 = 0
    16'b10000110_11101111 : OUT <= 0;  //134 / 239 = 0
    16'b10000110_11110000 : OUT <= 0;  //134 / 240 = 0
    16'b10000110_11110001 : OUT <= 0;  //134 / 241 = 0
    16'b10000110_11110010 : OUT <= 0;  //134 / 242 = 0
    16'b10000110_11110011 : OUT <= 0;  //134 / 243 = 0
    16'b10000110_11110100 : OUT <= 0;  //134 / 244 = 0
    16'b10000110_11110101 : OUT <= 0;  //134 / 245 = 0
    16'b10000110_11110110 : OUT <= 0;  //134 / 246 = 0
    16'b10000110_11110111 : OUT <= 0;  //134 / 247 = 0
    16'b10000110_11111000 : OUT <= 0;  //134 / 248 = 0
    16'b10000110_11111001 : OUT <= 0;  //134 / 249 = 0
    16'b10000110_11111010 : OUT <= 0;  //134 / 250 = 0
    16'b10000110_11111011 : OUT <= 0;  //134 / 251 = 0
    16'b10000110_11111100 : OUT <= 0;  //134 / 252 = 0
    16'b10000110_11111101 : OUT <= 0;  //134 / 253 = 0
    16'b10000110_11111110 : OUT <= 0;  //134 / 254 = 0
    16'b10000110_11111111 : OUT <= 0;  //134 / 255 = 0
    16'b10000111_00000000 : OUT <= 0;  //135 / 0 = 0
    16'b10000111_00000001 : OUT <= 135;  //135 / 1 = 135
    16'b10000111_00000010 : OUT <= 67;  //135 / 2 = 67
    16'b10000111_00000011 : OUT <= 45;  //135 / 3 = 45
    16'b10000111_00000100 : OUT <= 33;  //135 / 4 = 33
    16'b10000111_00000101 : OUT <= 27;  //135 / 5 = 27
    16'b10000111_00000110 : OUT <= 22;  //135 / 6 = 22
    16'b10000111_00000111 : OUT <= 19;  //135 / 7 = 19
    16'b10000111_00001000 : OUT <= 16;  //135 / 8 = 16
    16'b10000111_00001001 : OUT <= 15;  //135 / 9 = 15
    16'b10000111_00001010 : OUT <= 13;  //135 / 10 = 13
    16'b10000111_00001011 : OUT <= 12;  //135 / 11 = 12
    16'b10000111_00001100 : OUT <= 11;  //135 / 12 = 11
    16'b10000111_00001101 : OUT <= 10;  //135 / 13 = 10
    16'b10000111_00001110 : OUT <= 9;  //135 / 14 = 9
    16'b10000111_00001111 : OUT <= 9;  //135 / 15 = 9
    16'b10000111_00010000 : OUT <= 8;  //135 / 16 = 8
    16'b10000111_00010001 : OUT <= 7;  //135 / 17 = 7
    16'b10000111_00010010 : OUT <= 7;  //135 / 18 = 7
    16'b10000111_00010011 : OUT <= 7;  //135 / 19 = 7
    16'b10000111_00010100 : OUT <= 6;  //135 / 20 = 6
    16'b10000111_00010101 : OUT <= 6;  //135 / 21 = 6
    16'b10000111_00010110 : OUT <= 6;  //135 / 22 = 6
    16'b10000111_00010111 : OUT <= 5;  //135 / 23 = 5
    16'b10000111_00011000 : OUT <= 5;  //135 / 24 = 5
    16'b10000111_00011001 : OUT <= 5;  //135 / 25 = 5
    16'b10000111_00011010 : OUT <= 5;  //135 / 26 = 5
    16'b10000111_00011011 : OUT <= 5;  //135 / 27 = 5
    16'b10000111_00011100 : OUT <= 4;  //135 / 28 = 4
    16'b10000111_00011101 : OUT <= 4;  //135 / 29 = 4
    16'b10000111_00011110 : OUT <= 4;  //135 / 30 = 4
    16'b10000111_00011111 : OUT <= 4;  //135 / 31 = 4
    16'b10000111_00100000 : OUT <= 4;  //135 / 32 = 4
    16'b10000111_00100001 : OUT <= 4;  //135 / 33 = 4
    16'b10000111_00100010 : OUT <= 3;  //135 / 34 = 3
    16'b10000111_00100011 : OUT <= 3;  //135 / 35 = 3
    16'b10000111_00100100 : OUT <= 3;  //135 / 36 = 3
    16'b10000111_00100101 : OUT <= 3;  //135 / 37 = 3
    16'b10000111_00100110 : OUT <= 3;  //135 / 38 = 3
    16'b10000111_00100111 : OUT <= 3;  //135 / 39 = 3
    16'b10000111_00101000 : OUT <= 3;  //135 / 40 = 3
    16'b10000111_00101001 : OUT <= 3;  //135 / 41 = 3
    16'b10000111_00101010 : OUT <= 3;  //135 / 42 = 3
    16'b10000111_00101011 : OUT <= 3;  //135 / 43 = 3
    16'b10000111_00101100 : OUT <= 3;  //135 / 44 = 3
    16'b10000111_00101101 : OUT <= 3;  //135 / 45 = 3
    16'b10000111_00101110 : OUT <= 2;  //135 / 46 = 2
    16'b10000111_00101111 : OUT <= 2;  //135 / 47 = 2
    16'b10000111_00110000 : OUT <= 2;  //135 / 48 = 2
    16'b10000111_00110001 : OUT <= 2;  //135 / 49 = 2
    16'b10000111_00110010 : OUT <= 2;  //135 / 50 = 2
    16'b10000111_00110011 : OUT <= 2;  //135 / 51 = 2
    16'b10000111_00110100 : OUT <= 2;  //135 / 52 = 2
    16'b10000111_00110101 : OUT <= 2;  //135 / 53 = 2
    16'b10000111_00110110 : OUT <= 2;  //135 / 54 = 2
    16'b10000111_00110111 : OUT <= 2;  //135 / 55 = 2
    16'b10000111_00111000 : OUT <= 2;  //135 / 56 = 2
    16'b10000111_00111001 : OUT <= 2;  //135 / 57 = 2
    16'b10000111_00111010 : OUT <= 2;  //135 / 58 = 2
    16'b10000111_00111011 : OUT <= 2;  //135 / 59 = 2
    16'b10000111_00111100 : OUT <= 2;  //135 / 60 = 2
    16'b10000111_00111101 : OUT <= 2;  //135 / 61 = 2
    16'b10000111_00111110 : OUT <= 2;  //135 / 62 = 2
    16'b10000111_00111111 : OUT <= 2;  //135 / 63 = 2
    16'b10000111_01000000 : OUT <= 2;  //135 / 64 = 2
    16'b10000111_01000001 : OUT <= 2;  //135 / 65 = 2
    16'b10000111_01000010 : OUT <= 2;  //135 / 66 = 2
    16'b10000111_01000011 : OUT <= 2;  //135 / 67 = 2
    16'b10000111_01000100 : OUT <= 1;  //135 / 68 = 1
    16'b10000111_01000101 : OUT <= 1;  //135 / 69 = 1
    16'b10000111_01000110 : OUT <= 1;  //135 / 70 = 1
    16'b10000111_01000111 : OUT <= 1;  //135 / 71 = 1
    16'b10000111_01001000 : OUT <= 1;  //135 / 72 = 1
    16'b10000111_01001001 : OUT <= 1;  //135 / 73 = 1
    16'b10000111_01001010 : OUT <= 1;  //135 / 74 = 1
    16'b10000111_01001011 : OUT <= 1;  //135 / 75 = 1
    16'b10000111_01001100 : OUT <= 1;  //135 / 76 = 1
    16'b10000111_01001101 : OUT <= 1;  //135 / 77 = 1
    16'b10000111_01001110 : OUT <= 1;  //135 / 78 = 1
    16'b10000111_01001111 : OUT <= 1;  //135 / 79 = 1
    16'b10000111_01010000 : OUT <= 1;  //135 / 80 = 1
    16'b10000111_01010001 : OUT <= 1;  //135 / 81 = 1
    16'b10000111_01010010 : OUT <= 1;  //135 / 82 = 1
    16'b10000111_01010011 : OUT <= 1;  //135 / 83 = 1
    16'b10000111_01010100 : OUT <= 1;  //135 / 84 = 1
    16'b10000111_01010101 : OUT <= 1;  //135 / 85 = 1
    16'b10000111_01010110 : OUT <= 1;  //135 / 86 = 1
    16'b10000111_01010111 : OUT <= 1;  //135 / 87 = 1
    16'b10000111_01011000 : OUT <= 1;  //135 / 88 = 1
    16'b10000111_01011001 : OUT <= 1;  //135 / 89 = 1
    16'b10000111_01011010 : OUT <= 1;  //135 / 90 = 1
    16'b10000111_01011011 : OUT <= 1;  //135 / 91 = 1
    16'b10000111_01011100 : OUT <= 1;  //135 / 92 = 1
    16'b10000111_01011101 : OUT <= 1;  //135 / 93 = 1
    16'b10000111_01011110 : OUT <= 1;  //135 / 94 = 1
    16'b10000111_01011111 : OUT <= 1;  //135 / 95 = 1
    16'b10000111_01100000 : OUT <= 1;  //135 / 96 = 1
    16'b10000111_01100001 : OUT <= 1;  //135 / 97 = 1
    16'b10000111_01100010 : OUT <= 1;  //135 / 98 = 1
    16'b10000111_01100011 : OUT <= 1;  //135 / 99 = 1
    16'b10000111_01100100 : OUT <= 1;  //135 / 100 = 1
    16'b10000111_01100101 : OUT <= 1;  //135 / 101 = 1
    16'b10000111_01100110 : OUT <= 1;  //135 / 102 = 1
    16'b10000111_01100111 : OUT <= 1;  //135 / 103 = 1
    16'b10000111_01101000 : OUT <= 1;  //135 / 104 = 1
    16'b10000111_01101001 : OUT <= 1;  //135 / 105 = 1
    16'b10000111_01101010 : OUT <= 1;  //135 / 106 = 1
    16'b10000111_01101011 : OUT <= 1;  //135 / 107 = 1
    16'b10000111_01101100 : OUT <= 1;  //135 / 108 = 1
    16'b10000111_01101101 : OUT <= 1;  //135 / 109 = 1
    16'b10000111_01101110 : OUT <= 1;  //135 / 110 = 1
    16'b10000111_01101111 : OUT <= 1;  //135 / 111 = 1
    16'b10000111_01110000 : OUT <= 1;  //135 / 112 = 1
    16'b10000111_01110001 : OUT <= 1;  //135 / 113 = 1
    16'b10000111_01110010 : OUT <= 1;  //135 / 114 = 1
    16'b10000111_01110011 : OUT <= 1;  //135 / 115 = 1
    16'b10000111_01110100 : OUT <= 1;  //135 / 116 = 1
    16'b10000111_01110101 : OUT <= 1;  //135 / 117 = 1
    16'b10000111_01110110 : OUT <= 1;  //135 / 118 = 1
    16'b10000111_01110111 : OUT <= 1;  //135 / 119 = 1
    16'b10000111_01111000 : OUT <= 1;  //135 / 120 = 1
    16'b10000111_01111001 : OUT <= 1;  //135 / 121 = 1
    16'b10000111_01111010 : OUT <= 1;  //135 / 122 = 1
    16'b10000111_01111011 : OUT <= 1;  //135 / 123 = 1
    16'b10000111_01111100 : OUT <= 1;  //135 / 124 = 1
    16'b10000111_01111101 : OUT <= 1;  //135 / 125 = 1
    16'b10000111_01111110 : OUT <= 1;  //135 / 126 = 1
    16'b10000111_01111111 : OUT <= 1;  //135 / 127 = 1
    16'b10000111_10000000 : OUT <= 1;  //135 / 128 = 1
    16'b10000111_10000001 : OUT <= 1;  //135 / 129 = 1
    16'b10000111_10000010 : OUT <= 1;  //135 / 130 = 1
    16'b10000111_10000011 : OUT <= 1;  //135 / 131 = 1
    16'b10000111_10000100 : OUT <= 1;  //135 / 132 = 1
    16'b10000111_10000101 : OUT <= 1;  //135 / 133 = 1
    16'b10000111_10000110 : OUT <= 1;  //135 / 134 = 1
    16'b10000111_10000111 : OUT <= 1;  //135 / 135 = 1
    16'b10000111_10001000 : OUT <= 0;  //135 / 136 = 0
    16'b10000111_10001001 : OUT <= 0;  //135 / 137 = 0
    16'b10000111_10001010 : OUT <= 0;  //135 / 138 = 0
    16'b10000111_10001011 : OUT <= 0;  //135 / 139 = 0
    16'b10000111_10001100 : OUT <= 0;  //135 / 140 = 0
    16'b10000111_10001101 : OUT <= 0;  //135 / 141 = 0
    16'b10000111_10001110 : OUT <= 0;  //135 / 142 = 0
    16'b10000111_10001111 : OUT <= 0;  //135 / 143 = 0
    16'b10000111_10010000 : OUT <= 0;  //135 / 144 = 0
    16'b10000111_10010001 : OUT <= 0;  //135 / 145 = 0
    16'b10000111_10010010 : OUT <= 0;  //135 / 146 = 0
    16'b10000111_10010011 : OUT <= 0;  //135 / 147 = 0
    16'b10000111_10010100 : OUT <= 0;  //135 / 148 = 0
    16'b10000111_10010101 : OUT <= 0;  //135 / 149 = 0
    16'b10000111_10010110 : OUT <= 0;  //135 / 150 = 0
    16'b10000111_10010111 : OUT <= 0;  //135 / 151 = 0
    16'b10000111_10011000 : OUT <= 0;  //135 / 152 = 0
    16'b10000111_10011001 : OUT <= 0;  //135 / 153 = 0
    16'b10000111_10011010 : OUT <= 0;  //135 / 154 = 0
    16'b10000111_10011011 : OUT <= 0;  //135 / 155 = 0
    16'b10000111_10011100 : OUT <= 0;  //135 / 156 = 0
    16'b10000111_10011101 : OUT <= 0;  //135 / 157 = 0
    16'b10000111_10011110 : OUT <= 0;  //135 / 158 = 0
    16'b10000111_10011111 : OUT <= 0;  //135 / 159 = 0
    16'b10000111_10100000 : OUT <= 0;  //135 / 160 = 0
    16'b10000111_10100001 : OUT <= 0;  //135 / 161 = 0
    16'b10000111_10100010 : OUT <= 0;  //135 / 162 = 0
    16'b10000111_10100011 : OUT <= 0;  //135 / 163 = 0
    16'b10000111_10100100 : OUT <= 0;  //135 / 164 = 0
    16'b10000111_10100101 : OUT <= 0;  //135 / 165 = 0
    16'b10000111_10100110 : OUT <= 0;  //135 / 166 = 0
    16'b10000111_10100111 : OUT <= 0;  //135 / 167 = 0
    16'b10000111_10101000 : OUT <= 0;  //135 / 168 = 0
    16'b10000111_10101001 : OUT <= 0;  //135 / 169 = 0
    16'b10000111_10101010 : OUT <= 0;  //135 / 170 = 0
    16'b10000111_10101011 : OUT <= 0;  //135 / 171 = 0
    16'b10000111_10101100 : OUT <= 0;  //135 / 172 = 0
    16'b10000111_10101101 : OUT <= 0;  //135 / 173 = 0
    16'b10000111_10101110 : OUT <= 0;  //135 / 174 = 0
    16'b10000111_10101111 : OUT <= 0;  //135 / 175 = 0
    16'b10000111_10110000 : OUT <= 0;  //135 / 176 = 0
    16'b10000111_10110001 : OUT <= 0;  //135 / 177 = 0
    16'b10000111_10110010 : OUT <= 0;  //135 / 178 = 0
    16'b10000111_10110011 : OUT <= 0;  //135 / 179 = 0
    16'b10000111_10110100 : OUT <= 0;  //135 / 180 = 0
    16'b10000111_10110101 : OUT <= 0;  //135 / 181 = 0
    16'b10000111_10110110 : OUT <= 0;  //135 / 182 = 0
    16'b10000111_10110111 : OUT <= 0;  //135 / 183 = 0
    16'b10000111_10111000 : OUT <= 0;  //135 / 184 = 0
    16'b10000111_10111001 : OUT <= 0;  //135 / 185 = 0
    16'b10000111_10111010 : OUT <= 0;  //135 / 186 = 0
    16'b10000111_10111011 : OUT <= 0;  //135 / 187 = 0
    16'b10000111_10111100 : OUT <= 0;  //135 / 188 = 0
    16'b10000111_10111101 : OUT <= 0;  //135 / 189 = 0
    16'b10000111_10111110 : OUT <= 0;  //135 / 190 = 0
    16'b10000111_10111111 : OUT <= 0;  //135 / 191 = 0
    16'b10000111_11000000 : OUT <= 0;  //135 / 192 = 0
    16'b10000111_11000001 : OUT <= 0;  //135 / 193 = 0
    16'b10000111_11000010 : OUT <= 0;  //135 / 194 = 0
    16'b10000111_11000011 : OUT <= 0;  //135 / 195 = 0
    16'b10000111_11000100 : OUT <= 0;  //135 / 196 = 0
    16'b10000111_11000101 : OUT <= 0;  //135 / 197 = 0
    16'b10000111_11000110 : OUT <= 0;  //135 / 198 = 0
    16'b10000111_11000111 : OUT <= 0;  //135 / 199 = 0
    16'b10000111_11001000 : OUT <= 0;  //135 / 200 = 0
    16'b10000111_11001001 : OUT <= 0;  //135 / 201 = 0
    16'b10000111_11001010 : OUT <= 0;  //135 / 202 = 0
    16'b10000111_11001011 : OUT <= 0;  //135 / 203 = 0
    16'b10000111_11001100 : OUT <= 0;  //135 / 204 = 0
    16'b10000111_11001101 : OUT <= 0;  //135 / 205 = 0
    16'b10000111_11001110 : OUT <= 0;  //135 / 206 = 0
    16'b10000111_11001111 : OUT <= 0;  //135 / 207 = 0
    16'b10000111_11010000 : OUT <= 0;  //135 / 208 = 0
    16'b10000111_11010001 : OUT <= 0;  //135 / 209 = 0
    16'b10000111_11010010 : OUT <= 0;  //135 / 210 = 0
    16'b10000111_11010011 : OUT <= 0;  //135 / 211 = 0
    16'b10000111_11010100 : OUT <= 0;  //135 / 212 = 0
    16'b10000111_11010101 : OUT <= 0;  //135 / 213 = 0
    16'b10000111_11010110 : OUT <= 0;  //135 / 214 = 0
    16'b10000111_11010111 : OUT <= 0;  //135 / 215 = 0
    16'b10000111_11011000 : OUT <= 0;  //135 / 216 = 0
    16'b10000111_11011001 : OUT <= 0;  //135 / 217 = 0
    16'b10000111_11011010 : OUT <= 0;  //135 / 218 = 0
    16'b10000111_11011011 : OUT <= 0;  //135 / 219 = 0
    16'b10000111_11011100 : OUT <= 0;  //135 / 220 = 0
    16'b10000111_11011101 : OUT <= 0;  //135 / 221 = 0
    16'b10000111_11011110 : OUT <= 0;  //135 / 222 = 0
    16'b10000111_11011111 : OUT <= 0;  //135 / 223 = 0
    16'b10000111_11100000 : OUT <= 0;  //135 / 224 = 0
    16'b10000111_11100001 : OUT <= 0;  //135 / 225 = 0
    16'b10000111_11100010 : OUT <= 0;  //135 / 226 = 0
    16'b10000111_11100011 : OUT <= 0;  //135 / 227 = 0
    16'b10000111_11100100 : OUT <= 0;  //135 / 228 = 0
    16'b10000111_11100101 : OUT <= 0;  //135 / 229 = 0
    16'b10000111_11100110 : OUT <= 0;  //135 / 230 = 0
    16'b10000111_11100111 : OUT <= 0;  //135 / 231 = 0
    16'b10000111_11101000 : OUT <= 0;  //135 / 232 = 0
    16'b10000111_11101001 : OUT <= 0;  //135 / 233 = 0
    16'b10000111_11101010 : OUT <= 0;  //135 / 234 = 0
    16'b10000111_11101011 : OUT <= 0;  //135 / 235 = 0
    16'b10000111_11101100 : OUT <= 0;  //135 / 236 = 0
    16'b10000111_11101101 : OUT <= 0;  //135 / 237 = 0
    16'b10000111_11101110 : OUT <= 0;  //135 / 238 = 0
    16'b10000111_11101111 : OUT <= 0;  //135 / 239 = 0
    16'b10000111_11110000 : OUT <= 0;  //135 / 240 = 0
    16'b10000111_11110001 : OUT <= 0;  //135 / 241 = 0
    16'b10000111_11110010 : OUT <= 0;  //135 / 242 = 0
    16'b10000111_11110011 : OUT <= 0;  //135 / 243 = 0
    16'b10000111_11110100 : OUT <= 0;  //135 / 244 = 0
    16'b10000111_11110101 : OUT <= 0;  //135 / 245 = 0
    16'b10000111_11110110 : OUT <= 0;  //135 / 246 = 0
    16'b10000111_11110111 : OUT <= 0;  //135 / 247 = 0
    16'b10000111_11111000 : OUT <= 0;  //135 / 248 = 0
    16'b10000111_11111001 : OUT <= 0;  //135 / 249 = 0
    16'b10000111_11111010 : OUT <= 0;  //135 / 250 = 0
    16'b10000111_11111011 : OUT <= 0;  //135 / 251 = 0
    16'b10000111_11111100 : OUT <= 0;  //135 / 252 = 0
    16'b10000111_11111101 : OUT <= 0;  //135 / 253 = 0
    16'b10000111_11111110 : OUT <= 0;  //135 / 254 = 0
    16'b10000111_11111111 : OUT <= 0;  //135 / 255 = 0
    16'b10001000_00000000 : OUT <= 0;  //136 / 0 = 0
    16'b10001000_00000001 : OUT <= 136;  //136 / 1 = 136
    16'b10001000_00000010 : OUT <= 68;  //136 / 2 = 68
    16'b10001000_00000011 : OUT <= 45;  //136 / 3 = 45
    16'b10001000_00000100 : OUT <= 34;  //136 / 4 = 34
    16'b10001000_00000101 : OUT <= 27;  //136 / 5 = 27
    16'b10001000_00000110 : OUT <= 22;  //136 / 6 = 22
    16'b10001000_00000111 : OUT <= 19;  //136 / 7 = 19
    16'b10001000_00001000 : OUT <= 17;  //136 / 8 = 17
    16'b10001000_00001001 : OUT <= 15;  //136 / 9 = 15
    16'b10001000_00001010 : OUT <= 13;  //136 / 10 = 13
    16'b10001000_00001011 : OUT <= 12;  //136 / 11 = 12
    16'b10001000_00001100 : OUT <= 11;  //136 / 12 = 11
    16'b10001000_00001101 : OUT <= 10;  //136 / 13 = 10
    16'b10001000_00001110 : OUT <= 9;  //136 / 14 = 9
    16'b10001000_00001111 : OUT <= 9;  //136 / 15 = 9
    16'b10001000_00010000 : OUT <= 8;  //136 / 16 = 8
    16'b10001000_00010001 : OUT <= 8;  //136 / 17 = 8
    16'b10001000_00010010 : OUT <= 7;  //136 / 18 = 7
    16'b10001000_00010011 : OUT <= 7;  //136 / 19 = 7
    16'b10001000_00010100 : OUT <= 6;  //136 / 20 = 6
    16'b10001000_00010101 : OUT <= 6;  //136 / 21 = 6
    16'b10001000_00010110 : OUT <= 6;  //136 / 22 = 6
    16'b10001000_00010111 : OUT <= 5;  //136 / 23 = 5
    16'b10001000_00011000 : OUT <= 5;  //136 / 24 = 5
    16'b10001000_00011001 : OUT <= 5;  //136 / 25 = 5
    16'b10001000_00011010 : OUT <= 5;  //136 / 26 = 5
    16'b10001000_00011011 : OUT <= 5;  //136 / 27 = 5
    16'b10001000_00011100 : OUT <= 4;  //136 / 28 = 4
    16'b10001000_00011101 : OUT <= 4;  //136 / 29 = 4
    16'b10001000_00011110 : OUT <= 4;  //136 / 30 = 4
    16'b10001000_00011111 : OUT <= 4;  //136 / 31 = 4
    16'b10001000_00100000 : OUT <= 4;  //136 / 32 = 4
    16'b10001000_00100001 : OUT <= 4;  //136 / 33 = 4
    16'b10001000_00100010 : OUT <= 4;  //136 / 34 = 4
    16'b10001000_00100011 : OUT <= 3;  //136 / 35 = 3
    16'b10001000_00100100 : OUT <= 3;  //136 / 36 = 3
    16'b10001000_00100101 : OUT <= 3;  //136 / 37 = 3
    16'b10001000_00100110 : OUT <= 3;  //136 / 38 = 3
    16'b10001000_00100111 : OUT <= 3;  //136 / 39 = 3
    16'b10001000_00101000 : OUT <= 3;  //136 / 40 = 3
    16'b10001000_00101001 : OUT <= 3;  //136 / 41 = 3
    16'b10001000_00101010 : OUT <= 3;  //136 / 42 = 3
    16'b10001000_00101011 : OUT <= 3;  //136 / 43 = 3
    16'b10001000_00101100 : OUT <= 3;  //136 / 44 = 3
    16'b10001000_00101101 : OUT <= 3;  //136 / 45 = 3
    16'b10001000_00101110 : OUT <= 2;  //136 / 46 = 2
    16'b10001000_00101111 : OUT <= 2;  //136 / 47 = 2
    16'b10001000_00110000 : OUT <= 2;  //136 / 48 = 2
    16'b10001000_00110001 : OUT <= 2;  //136 / 49 = 2
    16'b10001000_00110010 : OUT <= 2;  //136 / 50 = 2
    16'b10001000_00110011 : OUT <= 2;  //136 / 51 = 2
    16'b10001000_00110100 : OUT <= 2;  //136 / 52 = 2
    16'b10001000_00110101 : OUT <= 2;  //136 / 53 = 2
    16'b10001000_00110110 : OUT <= 2;  //136 / 54 = 2
    16'b10001000_00110111 : OUT <= 2;  //136 / 55 = 2
    16'b10001000_00111000 : OUT <= 2;  //136 / 56 = 2
    16'b10001000_00111001 : OUT <= 2;  //136 / 57 = 2
    16'b10001000_00111010 : OUT <= 2;  //136 / 58 = 2
    16'b10001000_00111011 : OUT <= 2;  //136 / 59 = 2
    16'b10001000_00111100 : OUT <= 2;  //136 / 60 = 2
    16'b10001000_00111101 : OUT <= 2;  //136 / 61 = 2
    16'b10001000_00111110 : OUT <= 2;  //136 / 62 = 2
    16'b10001000_00111111 : OUT <= 2;  //136 / 63 = 2
    16'b10001000_01000000 : OUT <= 2;  //136 / 64 = 2
    16'b10001000_01000001 : OUT <= 2;  //136 / 65 = 2
    16'b10001000_01000010 : OUT <= 2;  //136 / 66 = 2
    16'b10001000_01000011 : OUT <= 2;  //136 / 67 = 2
    16'b10001000_01000100 : OUT <= 2;  //136 / 68 = 2
    16'b10001000_01000101 : OUT <= 1;  //136 / 69 = 1
    16'b10001000_01000110 : OUT <= 1;  //136 / 70 = 1
    16'b10001000_01000111 : OUT <= 1;  //136 / 71 = 1
    16'b10001000_01001000 : OUT <= 1;  //136 / 72 = 1
    16'b10001000_01001001 : OUT <= 1;  //136 / 73 = 1
    16'b10001000_01001010 : OUT <= 1;  //136 / 74 = 1
    16'b10001000_01001011 : OUT <= 1;  //136 / 75 = 1
    16'b10001000_01001100 : OUT <= 1;  //136 / 76 = 1
    16'b10001000_01001101 : OUT <= 1;  //136 / 77 = 1
    16'b10001000_01001110 : OUT <= 1;  //136 / 78 = 1
    16'b10001000_01001111 : OUT <= 1;  //136 / 79 = 1
    16'b10001000_01010000 : OUT <= 1;  //136 / 80 = 1
    16'b10001000_01010001 : OUT <= 1;  //136 / 81 = 1
    16'b10001000_01010010 : OUT <= 1;  //136 / 82 = 1
    16'b10001000_01010011 : OUT <= 1;  //136 / 83 = 1
    16'b10001000_01010100 : OUT <= 1;  //136 / 84 = 1
    16'b10001000_01010101 : OUT <= 1;  //136 / 85 = 1
    16'b10001000_01010110 : OUT <= 1;  //136 / 86 = 1
    16'b10001000_01010111 : OUT <= 1;  //136 / 87 = 1
    16'b10001000_01011000 : OUT <= 1;  //136 / 88 = 1
    16'b10001000_01011001 : OUT <= 1;  //136 / 89 = 1
    16'b10001000_01011010 : OUT <= 1;  //136 / 90 = 1
    16'b10001000_01011011 : OUT <= 1;  //136 / 91 = 1
    16'b10001000_01011100 : OUT <= 1;  //136 / 92 = 1
    16'b10001000_01011101 : OUT <= 1;  //136 / 93 = 1
    16'b10001000_01011110 : OUT <= 1;  //136 / 94 = 1
    16'b10001000_01011111 : OUT <= 1;  //136 / 95 = 1
    16'b10001000_01100000 : OUT <= 1;  //136 / 96 = 1
    16'b10001000_01100001 : OUT <= 1;  //136 / 97 = 1
    16'b10001000_01100010 : OUT <= 1;  //136 / 98 = 1
    16'b10001000_01100011 : OUT <= 1;  //136 / 99 = 1
    16'b10001000_01100100 : OUT <= 1;  //136 / 100 = 1
    16'b10001000_01100101 : OUT <= 1;  //136 / 101 = 1
    16'b10001000_01100110 : OUT <= 1;  //136 / 102 = 1
    16'b10001000_01100111 : OUT <= 1;  //136 / 103 = 1
    16'b10001000_01101000 : OUT <= 1;  //136 / 104 = 1
    16'b10001000_01101001 : OUT <= 1;  //136 / 105 = 1
    16'b10001000_01101010 : OUT <= 1;  //136 / 106 = 1
    16'b10001000_01101011 : OUT <= 1;  //136 / 107 = 1
    16'b10001000_01101100 : OUT <= 1;  //136 / 108 = 1
    16'b10001000_01101101 : OUT <= 1;  //136 / 109 = 1
    16'b10001000_01101110 : OUT <= 1;  //136 / 110 = 1
    16'b10001000_01101111 : OUT <= 1;  //136 / 111 = 1
    16'b10001000_01110000 : OUT <= 1;  //136 / 112 = 1
    16'b10001000_01110001 : OUT <= 1;  //136 / 113 = 1
    16'b10001000_01110010 : OUT <= 1;  //136 / 114 = 1
    16'b10001000_01110011 : OUT <= 1;  //136 / 115 = 1
    16'b10001000_01110100 : OUT <= 1;  //136 / 116 = 1
    16'b10001000_01110101 : OUT <= 1;  //136 / 117 = 1
    16'b10001000_01110110 : OUT <= 1;  //136 / 118 = 1
    16'b10001000_01110111 : OUT <= 1;  //136 / 119 = 1
    16'b10001000_01111000 : OUT <= 1;  //136 / 120 = 1
    16'b10001000_01111001 : OUT <= 1;  //136 / 121 = 1
    16'b10001000_01111010 : OUT <= 1;  //136 / 122 = 1
    16'b10001000_01111011 : OUT <= 1;  //136 / 123 = 1
    16'b10001000_01111100 : OUT <= 1;  //136 / 124 = 1
    16'b10001000_01111101 : OUT <= 1;  //136 / 125 = 1
    16'b10001000_01111110 : OUT <= 1;  //136 / 126 = 1
    16'b10001000_01111111 : OUT <= 1;  //136 / 127 = 1
    16'b10001000_10000000 : OUT <= 1;  //136 / 128 = 1
    16'b10001000_10000001 : OUT <= 1;  //136 / 129 = 1
    16'b10001000_10000010 : OUT <= 1;  //136 / 130 = 1
    16'b10001000_10000011 : OUT <= 1;  //136 / 131 = 1
    16'b10001000_10000100 : OUT <= 1;  //136 / 132 = 1
    16'b10001000_10000101 : OUT <= 1;  //136 / 133 = 1
    16'b10001000_10000110 : OUT <= 1;  //136 / 134 = 1
    16'b10001000_10000111 : OUT <= 1;  //136 / 135 = 1
    16'b10001000_10001000 : OUT <= 1;  //136 / 136 = 1
    16'b10001000_10001001 : OUT <= 0;  //136 / 137 = 0
    16'b10001000_10001010 : OUT <= 0;  //136 / 138 = 0
    16'b10001000_10001011 : OUT <= 0;  //136 / 139 = 0
    16'b10001000_10001100 : OUT <= 0;  //136 / 140 = 0
    16'b10001000_10001101 : OUT <= 0;  //136 / 141 = 0
    16'b10001000_10001110 : OUT <= 0;  //136 / 142 = 0
    16'b10001000_10001111 : OUT <= 0;  //136 / 143 = 0
    16'b10001000_10010000 : OUT <= 0;  //136 / 144 = 0
    16'b10001000_10010001 : OUT <= 0;  //136 / 145 = 0
    16'b10001000_10010010 : OUT <= 0;  //136 / 146 = 0
    16'b10001000_10010011 : OUT <= 0;  //136 / 147 = 0
    16'b10001000_10010100 : OUT <= 0;  //136 / 148 = 0
    16'b10001000_10010101 : OUT <= 0;  //136 / 149 = 0
    16'b10001000_10010110 : OUT <= 0;  //136 / 150 = 0
    16'b10001000_10010111 : OUT <= 0;  //136 / 151 = 0
    16'b10001000_10011000 : OUT <= 0;  //136 / 152 = 0
    16'b10001000_10011001 : OUT <= 0;  //136 / 153 = 0
    16'b10001000_10011010 : OUT <= 0;  //136 / 154 = 0
    16'b10001000_10011011 : OUT <= 0;  //136 / 155 = 0
    16'b10001000_10011100 : OUT <= 0;  //136 / 156 = 0
    16'b10001000_10011101 : OUT <= 0;  //136 / 157 = 0
    16'b10001000_10011110 : OUT <= 0;  //136 / 158 = 0
    16'b10001000_10011111 : OUT <= 0;  //136 / 159 = 0
    16'b10001000_10100000 : OUT <= 0;  //136 / 160 = 0
    16'b10001000_10100001 : OUT <= 0;  //136 / 161 = 0
    16'b10001000_10100010 : OUT <= 0;  //136 / 162 = 0
    16'b10001000_10100011 : OUT <= 0;  //136 / 163 = 0
    16'b10001000_10100100 : OUT <= 0;  //136 / 164 = 0
    16'b10001000_10100101 : OUT <= 0;  //136 / 165 = 0
    16'b10001000_10100110 : OUT <= 0;  //136 / 166 = 0
    16'b10001000_10100111 : OUT <= 0;  //136 / 167 = 0
    16'b10001000_10101000 : OUT <= 0;  //136 / 168 = 0
    16'b10001000_10101001 : OUT <= 0;  //136 / 169 = 0
    16'b10001000_10101010 : OUT <= 0;  //136 / 170 = 0
    16'b10001000_10101011 : OUT <= 0;  //136 / 171 = 0
    16'b10001000_10101100 : OUT <= 0;  //136 / 172 = 0
    16'b10001000_10101101 : OUT <= 0;  //136 / 173 = 0
    16'b10001000_10101110 : OUT <= 0;  //136 / 174 = 0
    16'b10001000_10101111 : OUT <= 0;  //136 / 175 = 0
    16'b10001000_10110000 : OUT <= 0;  //136 / 176 = 0
    16'b10001000_10110001 : OUT <= 0;  //136 / 177 = 0
    16'b10001000_10110010 : OUT <= 0;  //136 / 178 = 0
    16'b10001000_10110011 : OUT <= 0;  //136 / 179 = 0
    16'b10001000_10110100 : OUT <= 0;  //136 / 180 = 0
    16'b10001000_10110101 : OUT <= 0;  //136 / 181 = 0
    16'b10001000_10110110 : OUT <= 0;  //136 / 182 = 0
    16'b10001000_10110111 : OUT <= 0;  //136 / 183 = 0
    16'b10001000_10111000 : OUT <= 0;  //136 / 184 = 0
    16'b10001000_10111001 : OUT <= 0;  //136 / 185 = 0
    16'b10001000_10111010 : OUT <= 0;  //136 / 186 = 0
    16'b10001000_10111011 : OUT <= 0;  //136 / 187 = 0
    16'b10001000_10111100 : OUT <= 0;  //136 / 188 = 0
    16'b10001000_10111101 : OUT <= 0;  //136 / 189 = 0
    16'b10001000_10111110 : OUT <= 0;  //136 / 190 = 0
    16'b10001000_10111111 : OUT <= 0;  //136 / 191 = 0
    16'b10001000_11000000 : OUT <= 0;  //136 / 192 = 0
    16'b10001000_11000001 : OUT <= 0;  //136 / 193 = 0
    16'b10001000_11000010 : OUT <= 0;  //136 / 194 = 0
    16'b10001000_11000011 : OUT <= 0;  //136 / 195 = 0
    16'b10001000_11000100 : OUT <= 0;  //136 / 196 = 0
    16'b10001000_11000101 : OUT <= 0;  //136 / 197 = 0
    16'b10001000_11000110 : OUT <= 0;  //136 / 198 = 0
    16'b10001000_11000111 : OUT <= 0;  //136 / 199 = 0
    16'b10001000_11001000 : OUT <= 0;  //136 / 200 = 0
    16'b10001000_11001001 : OUT <= 0;  //136 / 201 = 0
    16'b10001000_11001010 : OUT <= 0;  //136 / 202 = 0
    16'b10001000_11001011 : OUT <= 0;  //136 / 203 = 0
    16'b10001000_11001100 : OUT <= 0;  //136 / 204 = 0
    16'b10001000_11001101 : OUT <= 0;  //136 / 205 = 0
    16'b10001000_11001110 : OUT <= 0;  //136 / 206 = 0
    16'b10001000_11001111 : OUT <= 0;  //136 / 207 = 0
    16'b10001000_11010000 : OUT <= 0;  //136 / 208 = 0
    16'b10001000_11010001 : OUT <= 0;  //136 / 209 = 0
    16'b10001000_11010010 : OUT <= 0;  //136 / 210 = 0
    16'b10001000_11010011 : OUT <= 0;  //136 / 211 = 0
    16'b10001000_11010100 : OUT <= 0;  //136 / 212 = 0
    16'b10001000_11010101 : OUT <= 0;  //136 / 213 = 0
    16'b10001000_11010110 : OUT <= 0;  //136 / 214 = 0
    16'b10001000_11010111 : OUT <= 0;  //136 / 215 = 0
    16'b10001000_11011000 : OUT <= 0;  //136 / 216 = 0
    16'b10001000_11011001 : OUT <= 0;  //136 / 217 = 0
    16'b10001000_11011010 : OUT <= 0;  //136 / 218 = 0
    16'b10001000_11011011 : OUT <= 0;  //136 / 219 = 0
    16'b10001000_11011100 : OUT <= 0;  //136 / 220 = 0
    16'b10001000_11011101 : OUT <= 0;  //136 / 221 = 0
    16'b10001000_11011110 : OUT <= 0;  //136 / 222 = 0
    16'b10001000_11011111 : OUT <= 0;  //136 / 223 = 0
    16'b10001000_11100000 : OUT <= 0;  //136 / 224 = 0
    16'b10001000_11100001 : OUT <= 0;  //136 / 225 = 0
    16'b10001000_11100010 : OUT <= 0;  //136 / 226 = 0
    16'b10001000_11100011 : OUT <= 0;  //136 / 227 = 0
    16'b10001000_11100100 : OUT <= 0;  //136 / 228 = 0
    16'b10001000_11100101 : OUT <= 0;  //136 / 229 = 0
    16'b10001000_11100110 : OUT <= 0;  //136 / 230 = 0
    16'b10001000_11100111 : OUT <= 0;  //136 / 231 = 0
    16'b10001000_11101000 : OUT <= 0;  //136 / 232 = 0
    16'b10001000_11101001 : OUT <= 0;  //136 / 233 = 0
    16'b10001000_11101010 : OUT <= 0;  //136 / 234 = 0
    16'b10001000_11101011 : OUT <= 0;  //136 / 235 = 0
    16'b10001000_11101100 : OUT <= 0;  //136 / 236 = 0
    16'b10001000_11101101 : OUT <= 0;  //136 / 237 = 0
    16'b10001000_11101110 : OUT <= 0;  //136 / 238 = 0
    16'b10001000_11101111 : OUT <= 0;  //136 / 239 = 0
    16'b10001000_11110000 : OUT <= 0;  //136 / 240 = 0
    16'b10001000_11110001 : OUT <= 0;  //136 / 241 = 0
    16'b10001000_11110010 : OUT <= 0;  //136 / 242 = 0
    16'b10001000_11110011 : OUT <= 0;  //136 / 243 = 0
    16'b10001000_11110100 : OUT <= 0;  //136 / 244 = 0
    16'b10001000_11110101 : OUT <= 0;  //136 / 245 = 0
    16'b10001000_11110110 : OUT <= 0;  //136 / 246 = 0
    16'b10001000_11110111 : OUT <= 0;  //136 / 247 = 0
    16'b10001000_11111000 : OUT <= 0;  //136 / 248 = 0
    16'b10001000_11111001 : OUT <= 0;  //136 / 249 = 0
    16'b10001000_11111010 : OUT <= 0;  //136 / 250 = 0
    16'b10001000_11111011 : OUT <= 0;  //136 / 251 = 0
    16'b10001000_11111100 : OUT <= 0;  //136 / 252 = 0
    16'b10001000_11111101 : OUT <= 0;  //136 / 253 = 0
    16'b10001000_11111110 : OUT <= 0;  //136 / 254 = 0
    16'b10001000_11111111 : OUT <= 0;  //136 / 255 = 0
    16'b10001001_00000000 : OUT <= 0;  //137 / 0 = 0
    16'b10001001_00000001 : OUT <= 137;  //137 / 1 = 137
    16'b10001001_00000010 : OUT <= 68;  //137 / 2 = 68
    16'b10001001_00000011 : OUT <= 45;  //137 / 3 = 45
    16'b10001001_00000100 : OUT <= 34;  //137 / 4 = 34
    16'b10001001_00000101 : OUT <= 27;  //137 / 5 = 27
    16'b10001001_00000110 : OUT <= 22;  //137 / 6 = 22
    16'b10001001_00000111 : OUT <= 19;  //137 / 7 = 19
    16'b10001001_00001000 : OUT <= 17;  //137 / 8 = 17
    16'b10001001_00001001 : OUT <= 15;  //137 / 9 = 15
    16'b10001001_00001010 : OUT <= 13;  //137 / 10 = 13
    16'b10001001_00001011 : OUT <= 12;  //137 / 11 = 12
    16'b10001001_00001100 : OUT <= 11;  //137 / 12 = 11
    16'b10001001_00001101 : OUT <= 10;  //137 / 13 = 10
    16'b10001001_00001110 : OUT <= 9;  //137 / 14 = 9
    16'b10001001_00001111 : OUT <= 9;  //137 / 15 = 9
    16'b10001001_00010000 : OUT <= 8;  //137 / 16 = 8
    16'b10001001_00010001 : OUT <= 8;  //137 / 17 = 8
    16'b10001001_00010010 : OUT <= 7;  //137 / 18 = 7
    16'b10001001_00010011 : OUT <= 7;  //137 / 19 = 7
    16'b10001001_00010100 : OUT <= 6;  //137 / 20 = 6
    16'b10001001_00010101 : OUT <= 6;  //137 / 21 = 6
    16'b10001001_00010110 : OUT <= 6;  //137 / 22 = 6
    16'b10001001_00010111 : OUT <= 5;  //137 / 23 = 5
    16'b10001001_00011000 : OUT <= 5;  //137 / 24 = 5
    16'b10001001_00011001 : OUT <= 5;  //137 / 25 = 5
    16'b10001001_00011010 : OUT <= 5;  //137 / 26 = 5
    16'b10001001_00011011 : OUT <= 5;  //137 / 27 = 5
    16'b10001001_00011100 : OUT <= 4;  //137 / 28 = 4
    16'b10001001_00011101 : OUT <= 4;  //137 / 29 = 4
    16'b10001001_00011110 : OUT <= 4;  //137 / 30 = 4
    16'b10001001_00011111 : OUT <= 4;  //137 / 31 = 4
    16'b10001001_00100000 : OUT <= 4;  //137 / 32 = 4
    16'b10001001_00100001 : OUT <= 4;  //137 / 33 = 4
    16'b10001001_00100010 : OUT <= 4;  //137 / 34 = 4
    16'b10001001_00100011 : OUT <= 3;  //137 / 35 = 3
    16'b10001001_00100100 : OUT <= 3;  //137 / 36 = 3
    16'b10001001_00100101 : OUT <= 3;  //137 / 37 = 3
    16'b10001001_00100110 : OUT <= 3;  //137 / 38 = 3
    16'b10001001_00100111 : OUT <= 3;  //137 / 39 = 3
    16'b10001001_00101000 : OUT <= 3;  //137 / 40 = 3
    16'b10001001_00101001 : OUT <= 3;  //137 / 41 = 3
    16'b10001001_00101010 : OUT <= 3;  //137 / 42 = 3
    16'b10001001_00101011 : OUT <= 3;  //137 / 43 = 3
    16'b10001001_00101100 : OUT <= 3;  //137 / 44 = 3
    16'b10001001_00101101 : OUT <= 3;  //137 / 45 = 3
    16'b10001001_00101110 : OUT <= 2;  //137 / 46 = 2
    16'b10001001_00101111 : OUT <= 2;  //137 / 47 = 2
    16'b10001001_00110000 : OUT <= 2;  //137 / 48 = 2
    16'b10001001_00110001 : OUT <= 2;  //137 / 49 = 2
    16'b10001001_00110010 : OUT <= 2;  //137 / 50 = 2
    16'b10001001_00110011 : OUT <= 2;  //137 / 51 = 2
    16'b10001001_00110100 : OUT <= 2;  //137 / 52 = 2
    16'b10001001_00110101 : OUT <= 2;  //137 / 53 = 2
    16'b10001001_00110110 : OUT <= 2;  //137 / 54 = 2
    16'b10001001_00110111 : OUT <= 2;  //137 / 55 = 2
    16'b10001001_00111000 : OUT <= 2;  //137 / 56 = 2
    16'b10001001_00111001 : OUT <= 2;  //137 / 57 = 2
    16'b10001001_00111010 : OUT <= 2;  //137 / 58 = 2
    16'b10001001_00111011 : OUT <= 2;  //137 / 59 = 2
    16'b10001001_00111100 : OUT <= 2;  //137 / 60 = 2
    16'b10001001_00111101 : OUT <= 2;  //137 / 61 = 2
    16'b10001001_00111110 : OUT <= 2;  //137 / 62 = 2
    16'b10001001_00111111 : OUT <= 2;  //137 / 63 = 2
    16'b10001001_01000000 : OUT <= 2;  //137 / 64 = 2
    16'b10001001_01000001 : OUT <= 2;  //137 / 65 = 2
    16'b10001001_01000010 : OUT <= 2;  //137 / 66 = 2
    16'b10001001_01000011 : OUT <= 2;  //137 / 67 = 2
    16'b10001001_01000100 : OUT <= 2;  //137 / 68 = 2
    16'b10001001_01000101 : OUT <= 1;  //137 / 69 = 1
    16'b10001001_01000110 : OUT <= 1;  //137 / 70 = 1
    16'b10001001_01000111 : OUT <= 1;  //137 / 71 = 1
    16'b10001001_01001000 : OUT <= 1;  //137 / 72 = 1
    16'b10001001_01001001 : OUT <= 1;  //137 / 73 = 1
    16'b10001001_01001010 : OUT <= 1;  //137 / 74 = 1
    16'b10001001_01001011 : OUT <= 1;  //137 / 75 = 1
    16'b10001001_01001100 : OUT <= 1;  //137 / 76 = 1
    16'b10001001_01001101 : OUT <= 1;  //137 / 77 = 1
    16'b10001001_01001110 : OUT <= 1;  //137 / 78 = 1
    16'b10001001_01001111 : OUT <= 1;  //137 / 79 = 1
    16'b10001001_01010000 : OUT <= 1;  //137 / 80 = 1
    16'b10001001_01010001 : OUT <= 1;  //137 / 81 = 1
    16'b10001001_01010010 : OUT <= 1;  //137 / 82 = 1
    16'b10001001_01010011 : OUT <= 1;  //137 / 83 = 1
    16'b10001001_01010100 : OUT <= 1;  //137 / 84 = 1
    16'b10001001_01010101 : OUT <= 1;  //137 / 85 = 1
    16'b10001001_01010110 : OUT <= 1;  //137 / 86 = 1
    16'b10001001_01010111 : OUT <= 1;  //137 / 87 = 1
    16'b10001001_01011000 : OUT <= 1;  //137 / 88 = 1
    16'b10001001_01011001 : OUT <= 1;  //137 / 89 = 1
    16'b10001001_01011010 : OUT <= 1;  //137 / 90 = 1
    16'b10001001_01011011 : OUT <= 1;  //137 / 91 = 1
    16'b10001001_01011100 : OUT <= 1;  //137 / 92 = 1
    16'b10001001_01011101 : OUT <= 1;  //137 / 93 = 1
    16'b10001001_01011110 : OUT <= 1;  //137 / 94 = 1
    16'b10001001_01011111 : OUT <= 1;  //137 / 95 = 1
    16'b10001001_01100000 : OUT <= 1;  //137 / 96 = 1
    16'b10001001_01100001 : OUT <= 1;  //137 / 97 = 1
    16'b10001001_01100010 : OUT <= 1;  //137 / 98 = 1
    16'b10001001_01100011 : OUT <= 1;  //137 / 99 = 1
    16'b10001001_01100100 : OUT <= 1;  //137 / 100 = 1
    16'b10001001_01100101 : OUT <= 1;  //137 / 101 = 1
    16'b10001001_01100110 : OUT <= 1;  //137 / 102 = 1
    16'b10001001_01100111 : OUT <= 1;  //137 / 103 = 1
    16'b10001001_01101000 : OUT <= 1;  //137 / 104 = 1
    16'b10001001_01101001 : OUT <= 1;  //137 / 105 = 1
    16'b10001001_01101010 : OUT <= 1;  //137 / 106 = 1
    16'b10001001_01101011 : OUT <= 1;  //137 / 107 = 1
    16'b10001001_01101100 : OUT <= 1;  //137 / 108 = 1
    16'b10001001_01101101 : OUT <= 1;  //137 / 109 = 1
    16'b10001001_01101110 : OUT <= 1;  //137 / 110 = 1
    16'b10001001_01101111 : OUT <= 1;  //137 / 111 = 1
    16'b10001001_01110000 : OUT <= 1;  //137 / 112 = 1
    16'b10001001_01110001 : OUT <= 1;  //137 / 113 = 1
    16'b10001001_01110010 : OUT <= 1;  //137 / 114 = 1
    16'b10001001_01110011 : OUT <= 1;  //137 / 115 = 1
    16'b10001001_01110100 : OUT <= 1;  //137 / 116 = 1
    16'b10001001_01110101 : OUT <= 1;  //137 / 117 = 1
    16'b10001001_01110110 : OUT <= 1;  //137 / 118 = 1
    16'b10001001_01110111 : OUT <= 1;  //137 / 119 = 1
    16'b10001001_01111000 : OUT <= 1;  //137 / 120 = 1
    16'b10001001_01111001 : OUT <= 1;  //137 / 121 = 1
    16'b10001001_01111010 : OUT <= 1;  //137 / 122 = 1
    16'b10001001_01111011 : OUT <= 1;  //137 / 123 = 1
    16'b10001001_01111100 : OUT <= 1;  //137 / 124 = 1
    16'b10001001_01111101 : OUT <= 1;  //137 / 125 = 1
    16'b10001001_01111110 : OUT <= 1;  //137 / 126 = 1
    16'b10001001_01111111 : OUT <= 1;  //137 / 127 = 1
    16'b10001001_10000000 : OUT <= 1;  //137 / 128 = 1
    16'b10001001_10000001 : OUT <= 1;  //137 / 129 = 1
    16'b10001001_10000010 : OUT <= 1;  //137 / 130 = 1
    16'b10001001_10000011 : OUT <= 1;  //137 / 131 = 1
    16'b10001001_10000100 : OUT <= 1;  //137 / 132 = 1
    16'b10001001_10000101 : OUT <= 1;  //137 / 133 = 1
    16'b10001001_10000110 : OUT <= 1;  //137 / 134 = 1
    16'b10001001_10000111 : OUT <= 1;  //137 / 135 = 1
    16'b10001001_10001000 : OUT <= 1;  //137 / 136 = 1
    16'b10001001_10001001 : OUT <= 1;  //137 / 137 = 1
    16'b10001001_10001010 : OUT <= 0;  //137 / 138 = 0
    16'b10001001_10001011 : OUT <= 0;  //137 / 139 = 0
    16'b10001001_10001100 : OUT <= 0;  //137 / 140 = 0
    16'b10001001_10001101 : OUT <= 0;  //137 / 141 = 0
    16'b10001001_10001110 : OUT <= 0;  //137 / 142 = 0
    16'b10001001_10001111 : OUT <= 0;  //137 / 143 = 0
    16'b10001001_10010000 : OUT <= 0;  //137 / 144 = 0
    16'b10001001_10010001 : OUT <= 0;  //137 / 145 = 0
    16'b10001001_10010010 : OUT <= 0;  //137 / 146 = 0
    16'b10001001_10010011 : OUT <= 0;  //137 / 147 = 0
    16'b10001001_10010100 : OUT <= 0;  //137 / 148 = 0
    16'b10001001_10010101 : OUT <= 0;  //137 / 149 = 0
    16'b10001001_10010110 : OUT <= 0;  //137 / 150 = 0
    16'b10001001_10010111 : OUT <= 0;  //137 / 151 = 0
    16'b10001001_10011000 : OUT <= 0;  //137 / 152 = 0
    16'b10001001_10011001 : OUT <= 0;  //137 / 153 = 0
    16'b10001001_10011010 : OUT <= 0;  //137 / 154 = 0
    16'b10001001_10011011 : OUT <= 0;  //137 / 155 = 0
    16'b10001001_10011100 : OUT <= 0;  //137 / 156 = 0
    16'b10001001_10011101 : OUT <= 0;  //137 / 157 = 0
    16'b10001001_10011110 : OUT <= 0;  //137 / 158 = 0
    16'b10001001_10011111 : OUT <= 0;  //137 / 159 = 0
    16'b10001001_10100000 : OUT <= 0;  //137 / 160 = 0
    16'b10001001_10100001 : OUT <= 0;  //137 / 161 = 0
    16'b10001001_10100010 : OUT <= 0;  //137 / 162 = 0
    16'b10001001_10100011 : OUT <= 0;  //137 / 163 = 0
    16'b10001001_10100100 : OUT <= 0;  //137 / 164 = 0
    16'b10001001_10100101 : OUT <= 0;  //137 / 165 = 0
    16'b10001001_10100110 : OUT <= 0;  //137 / 166 = 0
    16'b10001001_10100111 : OUT <= 0;  //137 / 167 = 0
    16'b10001001_10101000 : OUT <= 0;  //137 / 168 = 0
    16'b10001001_10101001 : OUT <= 0;  //137 / 169 = 0
    16'b10001001_10101010 : OUT <= 0;  //137 / 170 = 0
    16'b10001001_10101011 : OUT <= 0;  //137 / 171 = 0
    16'b10001001_10101100 : OUT <= 0;  //137 / 172 = 0
    16'b10001001_10101101 : OUT <= 0;  //137 / 173 = 0
    16'b10001001_10101110 : OUT <= 0;  //137 / 174 = 0
    16'b10001001_10101111 : OUT <= 0;  //137 / 175 = 0
    16'b10001001_10110000 : OUT <= 0;  //137 / 176 = 0
    16'b10001001_10110001 : OUT <= 0;  //137 / 177 = 0
    16'b10001001_10110010 : OUT <= 0;  //137 / 178 = 0
    16'b10001001_10110011 : OUT <= 0;  //137 / 179 = 0
    16'b10001001_10110100 : OUT <= 0;  //137 / 180 = 0
    16'b10001001_10110101 : OUT <= 0;  //137 / 181 = 0
    16'b10001001_10110110 : OUT <= 0;  //137 / 182 = 0
    16'b10001001_10110111 : OUT <= 0;  //137 / 183 = 0
    16'b10001001_10111000 : OUT <= 0;  //137 / 184 = 0
    16'b10001001_10111001 : OUT <= 0;  //137 / 185 = 0
    16'b10001001_10111010 : OUT <= 0;  //137 / 186 = 0
    16'b10001001_10111011 : OUT <= 0;  //137 / 187 = 0
    16'b10001001_10111100 : OUT <= 0;  //137 / 188 = 0
    16'b10001001_10111101 : OUT <= 0;  //137 / 189 = 0
    16'b10001001_10111110 : OUT <= 0;  //137 / 190 = 0
    16'b10001001_10111111 : OUT <= 0;  //137 / 191 = 0
    16'b10001001_11000000 : OUT <= 0;  //137 / 192 = 0
    16'b10001001_11000001 : OUT <= 0;  //137 / 193 = 0
    16'b10001001_11000010 : OUT <= 0;  //137 / 194 = 0
    16'b10001001_11000011 : OUT <= 0;  //137 / 195 = 0
    16'b10001001_11000100 : OUT <= 0;  //137 / 196 = 0
    16'b10001001_11000101 : OUT <= 0;  //137 / 197 = 0
    16'b10001001_11000110 : OUT <= 0;  //137 / 198 = 0
    16'b10001001_11000111 : OUT <= 0;  //137 / 199 = 0
    16'b10001001_11001000 : OUT <= 0;  //137 / 200 = 0
    16'b10001001_11001001 : OUT <= 0;  //137 / 201 = 0
    16'b10001001_11001010 : OUT <= 0;  //137 / 202 = 0
    16'b10001001_11001011 : OUT <= 0;  //137 / 203 = 0
    16'b10001001_11001100 : OUT <= 0;  //137 / 204 = 0
    16'b10001001_11001101 : OUT <= 0;  //137 / 205 = 0
    16'b10001001_11001110 : OUT <= 0;  //137 / 206 = 0
    16'b10001001_11001111 : OUT <= 0;  //137 / 207 = 0
    16'b10001001_11010000 : OUT <= 0;  //137 / 208 = 0
    16'b10001001_11010001 : OUT <= 0;  //137 / 209 = 0
    16'b10001001_11010010 : OUT <= 0;  //137 / 210 = 0
    16'b10001001_11010011 : OUT <= 0;  //137 / 211 = 0
    16'b10001001_11010100 : OUT <= 0;  //137 / 212 = 0
    16'b10001001_11010101 : OUT <= 0;  //137 / 213 = 0
    16'b10001001_11010110 : OUT <= 0;  //137 / 214 = 0
    16'b10001001_11010111 : OUT <= 0;  //137 / 215 = 0
    16'b10001001_11011000 : OUT <= 0;  //137 / 216 = 0
    16'b10001001_11011001 : OUT <= 0;  //137 / 217 = 0
    16'b10001001_11011010 : OUT <= 0;  //137 / 218 = 0
    16'b10001001_11011011 : OUT <= 0;  //137 / 219 = 0
    16'b10001001_11011100 : OUT <= 0;  //137 / 220 = 0
    16'b10001001_11011101 : OUT <= 0;  //137 / 221 = 0
    16'b10001001_11011110 : OUT <= 0;  //137 / 222 = 0
    16'b10001001_11011111 : OUT <= 0;  //137 / 223 = 0
    16'b10001001_11100000 : OUT <= 0;  //137 / 224 = 0
    16'b10001001_11100001 : OUT <= 0;  //137 / 225 = 0
    16'b10001001_11100010 : OUT <= 0;  //137 / 226 = 0
    16'b10001001_11100011 : OUT <= 0;  //137 / 227 = 0
    16'b10001001_11100100 : OUT <= 0;  //137 / 228 = 0
    16'b10001001_11100101 : OUT <= 0;  //137 / 229 = 0
    16'b10001001_11100110 : OUT <= 0;  //137 / 230 = 0
    16'b10001001_11100111 : OUT <= 0;  //137 / 231 = 0
    16'b10001001_11101000 : OUT <= 0;  //137 / 232 = 0
    16'b10001001_11101001 : OUT <= 0;  //137 / 233 = 0
    16'b10001001_11101010 : OUT <= 0;  //137 / 234 = 0
    16'b10001001_11101011 : OUT <= 0;  //137 / 235 = 0
    16'b10001001_11101100 : OUT <= 0;  //137 / 236 = 0
    16'b10001001_11101101 : OUT <= 0;  //137 / 237 = 0
    16'b10001001_11101110 : OUT <= 0;  //137 / 238 = 0
    16'b10001001_11101111 : OUT <= 0;  //137 / 239 = 0
    16'b10001001_11110000 : OUT <= 0;  //137 / 240 = 0
    16'b10001001_11110001 : OUT <= 0;  //137 / 241 = 0
    16'b10001001_11110010 : OUT <= 0;  //137 / 242 = 0
    16'b10001001_11110011 : OUT <= 0;  //137 / 243 = 0
    16'b10001001_11110100 : OUT <= 0;  //137 / 244 = 0
    16'b10001001_11110101 : OUT <= 0;  //137 / 245 = 0
    16'b10001001_11110110 : OUT <= 0;  //137 / 246 = 0
    16'b10001001_11110111 : OUT <= 0;  //137 / 247 = 0
    16'b10001001_11111000 : OUT <= 0;  //137 / 248 = 0
    16'b10001001_11111001 : OUT <= 0;  //137 / 249 = 0
    16'b10001001_11111010 : OUT <= 0;  //137 / 250 = 0
    16'b10001001_11111011 : OUT <= 0;  //137 / 251 = 0
    16'b10001001_11111100 : OUT <= 0;  //137 / 252 = 0
    16'b10001001_11111101 : OUT <= 0;  //137 / 253 = 0
    16'b10001001_11111110 : OUT <= 0;  //137 / 254 = 0
    16'b10001001_11111111 : OUT <= 0;  //137 / 255 = 0
    16'b10001010_00000000 : OUT <= 0;  //138 / 0 = 0
    16'b10001010_00000001 : OUT <= 138;  //138 / 1 = 138
    16'b10001010_00000010 : OUT <= 69;  //138 / 2 = 69
    16'b10001010_00000011 : OUT <= 46;  //138 / 3 = 46
    16'b10001010_00000100 : OUT <= 34;  //138 / 4 = 34
    16'b10001010_00000101 : OUT <= 27;  //138 / 5 = 27
    16'b10001010_00000110 : OUT <= 23;  //138 / 6 = 23
    16'b10001010_00000111 : OUT <= 19;  //138 / 7 = 19
    16'b10001010_00001000 : OUT <= 17;  //138 / 8 = 17
    16'b10001010_00001001 : OUT <= 15;  //138 / 9 = 15
    16'b10001010_00001010 : OUT <= 13;  //138 / 10 = 13
    16'b10001010_00001011 : OUT <= 12;  //138 / 11 = 12
    16'b10001010_00001100 : OUT <= 11;  //138 / 12 = 11
    16'b10001010_00001101 : OUT <= 10;  //138 / 13 = 10
    16'b10001010_00001110 : OUT <= 9;  //138 / 14 = 9
    16'b10001010_00001111 : OUT <= 9;  //138 / 15 = 9
    16'b10001010_00010000 : OUT <= 8;  //138 / 16 = 8
    16'b10001010_00010001 : OUT <= 8;  //138 / 17 = 8
    16'b10001010_00010010 : OUT <= 7;  //138 / 18 = 7
    16'b10001010_00010011 : OUT <= 7;  //138 / 19 = 7
    16'b10001010_00010100 : OUT <= 6;  //138 / 20 = 6
    16'b10001010_00010101 : OUT <= 6;  //138 / 21 = 6
    16'b10001010_00010110 : OUT <= 6;  //138 / 22 = 6
    16'b10001010_00010111 : OUT <= 6;  //138 / 23 = 6
    16'b10001010_00011000 : OUT <= 5;  //138 / 24 = 5
    16'b10001010_00011001 : OUT <= 5;  //138 / 25 = 5
    16'b10001010_00011010 : OUT <= 5;  //138 / 26 = 5
    16'b10001010_00011011 : OUT <= 5;  //138 / 27 = 5
    16'b10001010_00011100 : OUT <= 4;  //138 / 28 = 4
    16'b10001010_00011101 : OUT <= 4;  //138 / 29 = 4
    16'b10001010_00011110 : OUT <= 4;  //138 / 30 = 4
    16'b10001010_00011111 : OUT <= 4;  //138 / 31 = 4
    16'b10001010_00100000 : OUT <= 4;  //138 / 32 = 4
    16'b10001010_00100001 : OUT <= 4;  //138 / 33 = 4
    16'b10001010_00100010 : OUT <= 4;  //138 / 34 = 4
    16'b10001010_00100011 : OUT <= 3;  //138 / 35 = 3
    16'b10001010_00100100 : OUT <= 3;  //138 / 36 = 3
    16'b10001010_00100101 : OUT <= 3;  //138 / 37 = 3
    16'b10001010_00100110 : OUT <= 3;  //138 / 38 = 3
    16'b10001010_00100111 : OUT <= 3;  //138 / 39 = 3
    16'b10001010_00101000 : OUT <= 3;  //138 / 40 = 3
    16'b10001010_00101001 : OUT <= 3;  //138 / 41 = 3
    16'b10001010_00101010 : OUT <= 3;  //138 / 42 = 3
    16'b10001010_00101011 : OUT <= 3;  //138 / 43 = 3
    16'b10001010_00101100 : OUT <= 3;  //138 / 44 = 3
    16'b10001010_00101101 : OUT <= 3;  //138 / 45 = 3
    16'b10001010_00101110 : OUT <= 3;  //138 / 46 = 3
    16'b10001010_00101111 : OUT <= 2;  //138 / 47 = 2
    16'b10001010_00110000 : OUT <= 2;  //138 / 48 = 2
    16'b10001010_00110001 : OUT <= 2;  //138 / 49 = 2
    16'b10001010_00110010 : OUT <= 2;  //138 / 50 = 2
    16'b10001010_00110011 : OUT <= 2;  //138 / 51 = 2
    16'b10001010_00110100 : OUT <= 2;  //138 / 52 = 2
    16'b10001010_00110101 : OUT <= 2;  //138 / 53 = 2
    16'b10001010_00110110 : OUT <= 2;  //138 / 54 = 2
    16'b10001010_00110111 : OUT <= 2;  //138 / 55 = 2
    16'b10001010_00111000 : OUT <= 2;  //138 / 56 = 2
    16'b10001010_00111001 : OUT <= 2;  //138 / 57 = 2
    16'b10001010_00111010 : OUT <= 2;  //138 / 58 = 2
    16'b10001010_00111011 : OUT <= 2;  //138 / 59 = 2
    16'b10001010_00111100 : OUT <= 2;  //138 / 60 = 2
    16'b10001010_00111101 : OUT <= 2;  //138 / 61 = 2
    16'b10001010_00111110 : OUT <= 2;  //138 / 62 = 2
    16'b10001010_00111111 : OUT <= 2;  //138 / 63 = 2
    16'b10001010_01000000 : OUT <= 2;  //138 / 64 = 2
    16'b10001010_01000001 : OUT <= 2;  //138 / 65 = 2
    16'b10001010_01000010 : OUT <= 2;  //138 / 66 = 2
    16'b10001010_01000011 : OUT <= 2;  //138 / 67 = 2
    16'b10001010_01000100 : OUT <= 2;  //138 / 68 = 2
    16'b10001010_01000101 : OUT <= 2;  //138 / 69 = 2
    16'b10001010_01000110 : OUT <= 1;  //138 / 70 = 1
    16'b10001010_01000111 : OUT <= 1;  //138 / 71 = 1
    16'b10001010_01001000 : OUT <= 1;  //138 / 72 = 1
    16'b10001010_01001001 : OUT <= 1;  //138 / 73 = 1
    16'b10001010_01001010 : OUT <= 1;  //138 / 74 = 1
    16'b10001010_01001011 : OUT <= 1;  //138 / 75 = 1
    16'b10001010_01001100 : OUT <= 1;  //138 / 76 = 1
    16'b10001010_01001101 : OUT <= 1;  //138 / 77 = 1
    16'b10001010_01001110 : OUT <= 1;  //138 / 78 = 1
    16'b10001010_01001111 : OUT <= 1;  //138 / 79 = 1
    16'b10001010_01010000 : OUT <= 1;  //138 / 80 = 1
    16'b10001010_01010001 : OUT <= 1;  //138 / 81 = 1
    16'b10001010_01010010 : OUT <= 1;  //138 / 82 = 1
    16'b10001010_01010011 : OUT <= 1;  //138 / 83 = 1
    16'b10001010_01010100 : OUT <= 1;  //138 / 84 = 1
    16'b10001010_01010101 : OUT <= 1;  //138 / 85 = 1
    16'b10001010_01010110 : OUT <= 1;  //138 / 86 = 1
    16'b10001010_01010111 : OUT <= 1;  //138 / 87 = 1
    16'b10001010_01011000 : OUT <= 1;  //138 / 88 = 1
    16'b10001010_01011001 : OUT <= 1;  //138 / 89 = 1
    16'b10001010_01011010 : OUT <= 1;  //138 / 90 = 1
    16'b10001010_01011011 : OUT <= 1;  //138 / 91 = 1
    16'b10001010_01011100 : OUT <= 1;  //138 / 92 = 1
    16'b10001010_01011101 : OUT <= 1;  //138 / 93 = 1
    16'b10001010_01011110 : OUT <= 1;  //138 / 94 = 1
    16'b10001010_01011111 : OUT <= 1;  //138 / 95 = 1
    16'b10001010_01100000 : OUT <= 1;  //138 / 96 = 1
    16'b10001010_01100001 : OUT <= 1;  //138 / 97 = 1
    16'b10001010_01100010 : OUT <= 1;  //138 / 98 = 1
    16'b10001010_01100011 : OUT <= 1;  //138 / 99 = 1
    16'b10001010_01100100 : OUT <= 1;  //138 / 100 = 1
    16'b10001010_01100101 : OUT <= 1;  //138 / 101 = 1
    16'b10001010_01100110 : OUT <= 1;  //138 / 102 = 1
    16'b10001010_01100111 : OUT <= 1;  //138 / 103 = 1
    16'b10001010_01101000 : OUT <= 1;  //138 / 104 = 1
    16'b10001010_01101001 : OUT <= 1;  //138 / 105 = 1
    16'b10001010_01101010 : OUT <= 1;  //138 / 106 = 1
    16'b10001010_01101011 : OUT <= 1;  //138 / 107 = 1
    16'b10001010_01101100 : OUT <= 1;  //138 / 108 = 1
    16'b10001010_01101101 : OUT <= 1;  //138 / 109 = 1
    16'b10001010_01101110 : OUT <= 1;  //138 / 110 = 1
    16'b10001010_01101111 : OUT <= 1;  //138 / 111 = 1
    16'b10001010_01110000 : OUT <= 1;  //138 / 112 = 1
    16'b10001010_01110001 : OUT <= 1;  //138 / 113 = 1
    16'b10001010_01110010 : OUT <= 1;  //138 / 114 = 1
    16'b10001010_01110011 : OUT <= 1;  //138 / 115 = 1
    16'b10001010_01110100 : OUT <= 1;  //138 / 116 = 1
    16'b10001010_01110101 : OUT <= 1;  //138 / 117 = 1
    16'b10001010_01110110 : OUT <= 1;  //138 / 118 = 1
    16'b10001010_01110111 : OUT <= 1;  //138 / 119 = 1
    16'b10001010_01111000 : OUT <= 1;  //138 / 120 = 1
    16'b10001010_01111001 : OUT <= 1;  //138 / 121 = 1
    16'b10001010_01111010 : OUT <= 1;  //138 / 122 = 1
    16'b10001010_01111011 : OUT <= 1;  //138 / 123 = 1
    16'b10001010_01111100 : OUT <= 1;  //138 / 124 = 1
    16'b10001010_01111101 : OUT <= 1;  //138 / 125 = 1
    16'b10001010_01111110 : OUT <= 1;  //138 / 126 = 1
    16'b10001010_01111111 : OUT <= 1;  //138 / 127 = 1
    16'b10001010_10000000 : OUT <= 1;  //138 / 128 = 1
    16'b10001010_10000001 : OUT <= 1;  //138 / 129 = 1
    16'b10001010_10000010 : OUT <= 1;  //138 / 130 = 1
    16'b10001010_10000011 : OUT <= 1;  //138 / 131 = 1
    16'b10001010_10000100 : OUT <= 1;  //138 / 132 = 1
    16'b10001010_10000101 : OUT <= 1;  //138 / 133 = 1
    16'b10001010_10000110 : OUT <= 1;  //138 / 134 = 1
    16'b10001010_10000111 : OUT <= 1;  //138 / 135 = 1
    16'b10001010_10001000 : OUT <= 1;  //138 / 136 = 1
    16'b10001010_10001001 : OUT <= 1;  //138 / 137 = 1
    16'b10001010_10001010 : OUT <= 1;  //138 / 138 = 1
    16'b10001010_10001011 : OUT <= 0;  //138 / 139 = 0
    16'b10001010_10001100 : OUT <= 0;  //138 / 140 = 0
    16'b10001010_10001101 : OUT <= 0;  //138 / 141 = 0
    16'b10001010_10001110 : OUT <= 0;  //138 / 142 = 0
    16'b10001010_10001111 : OUT <= 0;  //138 / 143 = 0
    16'b10001010_10010000 : OUT <= 0;  //138 / 144 = 0
    16'b10001010_10010001 : OUT <= 0;  //138 / 145 = 0
    16'b10001010_10010010 : OUT <= 0;  //138 / 146 = 0
    16'b10001010_10010011 : OUT <= 0;  //138 / 147 = 0
    16'b10001010_10010100 : OUT <= 0;  //138 / 148 = 0
    16'b10001010_10010101 : OUT <= 0;  //138 / 149 = 0
    16'b10001010_10010110 : OUT <= 0;  //138 / 150 = 0
    16'b10001010_10010111 : OUT <= 0;  //138 / 151 = 0
    16'b10001010_10011000 : OUT <= 0;  //138 / 152 = 0
    16'b10001010_10011001 : OUT <= 0;  //138 / 153 = 0
    16'b10001010_10011010 : OUT <= 0;  //138 / 154 = 0
    16'b10001010_10011011 : OUT <= 0;  //138 / 155 = 0
    16'b10001010_10011100 : OUT <= 0;  //138 / 156 = 0
    16'b10001010_10011101 : OUT <= 0;  //138 / 157 = 0
    16'b10001010_10011110 : OUT <= 0;  //138 / 158 = 0
    16'b10001010_10011111 : OUT <= 0;  //138 / 159 = 0
    16'b10001010_10100000 : OUT <= 0;  //138 / 160 = 0
    16'b10001010_10100001 : OUT <= 0;  //138 / 161 = 0
    16'b10001010_10100010 : OUT <= 0;  //138 / 162 = 0
    16'b10001010_10100011 : OUT <= 0;  //138 / 163 = 0
    16'b10001010_10100100 : OUT <= 0;  //138 / 164 = 0
    16'b10001010_10100101 : OUT <= 0;  //138 / 165 = 0
    16'b10001010_10100110 : OUT <= 0;  //138 / 166 = 0
    16'b10001010_10100111 : OUT <= 0;  //138 / 167 = 0
    16'b10001010_10101000 : OUT <= 0;  //138 / 168 = 0
    16'b10001010_10101001 : OUT <= 0;  //138 / 169 = 0
    16'b10001010_10101010 : OUT <= 0;  //138 / 170 = 0
    16'b10001010_10101011 : OUT <= 0;  //138 / 171 = 0
    16'b10001010_10101100 : OUT <= 0;  //138 / 172 = 0
    16'b10001010_10101101 : OUT <= 0;  //138 / 173 = 0
    16'b10001010_10101110 : OUT <= 0;  //138 / 174 = 0
    16'b10001010_10101111 : OUT <= 0;  //138 / 175 = 0
    16'b10001010_10110000 : OUT <= 0;  //138 / 176 = 0
    16'b10001010_10110001 : OUT <= 0;  //138 / 177 = 0
    16'b10001010_10110010 : OUT <= 0;  //138 / 178 = 0
    16'b10001010_10110011 : OUT <= 0;  //138 / 179 = 0
    16'b10001010_10110100 : OUT <= 0;  //138 / 180 = 0
    16'b10001010_10110101 : OUT <= 0;  //138 / 181 = 0
    16'b10001010_10110110 : OUT <= 0;  //138 / 182 = 0
    16'b10001010_10110111 : OUT <= 0;  //138 / 183 = 0
    16'b10001010_10111000 : OUT <= 0;  //138 / 184 = 0
    16'b10001010_10111001 : OUT <= 0;  //138 / 185 = 0
    16'b10001010_10111010 : OUT <= 0;  //138 / 186 = 0
    16'b10001010_10111011 : OUT <= 0;  //138 / 187 = 0
    16'b10001010_10111100 : OUT <= 0;  //138 / 188 = 0
    16'b10001010_10111101 : OUT <= 0;  //138 / 189 = 0
    16'b10001010_10111110 : OUT <= 0;  //138 / 190 = 0
    16'b10001010_10111111 : OUT <= 0;  //138 / 191 = 0
    16'b10001010_11000000 : OUT <= 0;  //138 / 192 = 0
    16'b10001010_11000001 : OUT <= 0;  //138 / 193 = 0
    16'b10001010_11000010 : OUT <= 0;  //138 / 194 = 0
    16'b10001010_11000011 : OUT <= 0;  //138 / 195 = 0
    16'b10001010_11000100 : OUT <= 0;  //138 / 196 = 0
    16'b10001010_11000101 : OUT <= 0;  //138 / 197 = 0
    16'b10001010_11000110 : OUT <= 0;  //138 / 198 = 0
    16'b10001010_11000111 : OUT <= 0;  //138 / 199 = 0
    16'b10001010_11001000 : OUT <= 0;  //138 / 200 = 0
    16'b10001010_11001001 : OUT <= 0;  //138 / 201 = 0
    16'b10001010_11001010 : OUT <= 0;  //138 / 202 = 0
    16'b10001010_11001011 : OUT <= 0;  //138 / 203 = 0
    16'b10001010_11001100 : OUT <= 0;  //138 / 204 = 0
    16'b10001010_11001101 : OUT <= 0;  //138 / 205 = 0
    16'b10001010_11001110 : OUT <= 0;  //138 / 206 = 0
    16'b10001010_11001111 : OUT <= 0;  //138 / 207 = 0
    16'b10001010_11010000 : OUT <= 0;  //138 / 208 = 0
    16'b10001010_11010001 : OUT <= 0;  //138 / 209 = 0
    16'b10001010_11010010 : OUT <= 0;  //138 / 210 = 0
    16'b10001010_11010011 : OUT <= 0;  //138 / 211 = 0
    16'b10001010_11010100 : OUT <= 0;  //138 / 212 = 0
    16'b10001010_11010101 : OUT <= 0;  //138 / 213 = 0
    16'b10001010_11010110 : OUT <= 0;  //138 / 214 = 0
    16'b10001010_11010111 : OUT <= 0;  //138 / 215 = 0
    16'b10001010_11011000 : OUT <= 0;  //138 / 216 = 0
    16'b10001010_11011001 : OUT <= 0;  //138 / 217 = 0
    16'b10001010_11011010 : OUT <= 0;  //138 / 218 = 0
    16'b10001010_11011011 : OUT <= 0;  //138 / 219 = 0
    16'b10001010_11011100 : OUT <= 0;  //138 / 220 = 0
    16'b10001010_11011101 : OUT <= 0;  //138 / 221 = 0
    16'b10001010_11011110 : OUT <= 0;  //138 / 222 = 0
    16'b10001010_11011111 : OUT <= 0;  //138 / 223 = 0
    16'b10001010_11100000 : OUT <= 0;  //138 / 224 = 0
    16'b10001010_11100001 : OUT <= 0;  //138 / 225 = 0
    16'b10001010_11100010 : OUT <= 0;  //138 / 226 = 0
    16'b10001010_11100011 : OUT <= 0;  //138 / 227 = 0
    16'b10001010_11100100 : OUT <= 0;  //138 / 228 = 0
    16'b10001010_11100101 : OUT <= 0;  //138 / 229 = 0
    16'b10001010_11100110 : OUT <= 0;  //138 / 230 = 0
    16'b10001010_11100111 : OUT <= 0;  //138 / 231 = 0
    16'b10001010_11101000 : OUT <= 0;  //138 / 232 = 0
    16'b10001010_11101001 : OUT <= 0;  //138 / 233 = 0
    16'b10001010_11101010 : OUT <= 0;  //138 / 234 = 0
    16'b10001010_11101011 : OUT <= 0;  //138 / 235 = 0
    16'b10001010_11101100 : OUT <= 0;  //138 / 236 = 0
    16'b10001010_11101101 : OUT <= 0;  //138 / 237 = 0
    16'b10001010_11101110 : OUT <= 0;  //138 / 238 = 0
    16'b10001010_11101111 : OUT <= 0;  //138 / 239 = 0
    16'b10001010_11110000 : OUT <= 0;  //138 / 240 = 0
    16'b10001010_11110001 : OUT <= 0;  //138 / 241 = 0
    16'b10001010_11110010 : OUT <= 0;  //138 / 242 = 0
    16'b10001010_11110011 : OUT <= 0;  //138 / 243 = 0
    16'b10001010_11110100 : OUT <= 0;  //138 / 244 = 0
    16'b10001010_11110101 : OUT <= 0;  //138 / 245 = 0
    16'b10001010_11110110 : OUT <= 0;  //138 / 246 = 0
    16'b10001010_11110111 : OUT <= 0;  //138 / 247 = 0
    16'b10001010_11111000 : OUT <= 0;  //138 / 248 = 0
    16'b10001010_11111001 : OUT <= 0;  //138 / 249 = 0
    16'b10001010_11111010 : OUT <= 0;  //138 / 250 = 0
    16'b10001010_11111011 : OUT <= 0;  //138 / 251 = 0
    16'b10001010_11111100 : OUT <= 0;  //138 / 252 = 0
    16'b10001010_11111101 : OUT <= 0;  //138 / 253 = 0
    16'b10001010_11111110 : OUT <= 0;  //138 / 254 = 0
    16'b10001010_11111111 : OUT <= 0;  //138 / 255 = 0
    16'b10001011_00000000 : OUT <= 0;  //139 / 0 = 0
    16'b10001011_00000001 : OUT <= 139;  //139 / 1 = 139
    16'b10001011_00000010 : OUT <= 69;  //139 / 2 = 69
    16'b10001011_00000011 : OUT <= 46;  //139 / 3 = 46
    16'b10001011_00000100 : OUT <= 34;  //139 / 4 = 34
    16'b10001011_00000101 : OUT <= 27;  //139 / 5 = 27
    16'b10001011_00000110 : OUT <= 23;  //139 / 6 = 23
    16'b10001011_00000111 : OUT <= 19;  //139 / 7 = 19
    16'b10001011_00001000 : OUT <= 17;  //139 / 8 = 17
    16'b10001011_00001001 : OUT <= 15;  //139 / 9 = 15
    16'b10001011_00001010 : OUT <= 13;  //139 / 10 = 13
    16'b10001011_00001011 : OUT <= 12;  //139 / 11 = 12
    16'b10001011_00001100 : OUT <= 11;  //139 / 12 = 11
    16'b10001011_00001101 : OUT <= 10;  //139 / 13 = 10
    16'b10001011_00001110 : OUT <= 9;  //139 / 14 = 9
    16'b10001011_00001111 : OUT <= 9;  //139 / 15 = 9
    16'b10001011_00010000 : OUT <= 8;  //139 / 16 = 8
    16'b10001011_00010001 : OUT <= 8;  //139 / 17 = 8
    16'b10001011_00010010 : OUT <= 7;  //139 / 18 = 7
    16'b10001011_00010011 : OUT <= 7;  //139 / 19 = 7
    16'b10001011_00010100 : OUT <= 6;  //139 / 20 = 6
    16'b10001011_00010101 : OUT <= 6;  //139 / 21 = 6
    16'b10001011_00010110 : OUT <= 6;  //139 / 22 = 6
    16'b10001011_00010111 : OUT <= 6;  //139 / 23 = 6
    16'b10001011_00011000 : OUT <= 5;  //139 / 24 = 5
    16'b10001011_00011001 : OUT <= 5;  //139 / 25 = 5
    16'b10001011_00011010 : OUT <= 5;  //139 / 26 = 5
    16'b10001011_00011011 : OUT <= 5;  //139 / 27 = 5
    16'b10001011_00011100 : OUT <= 4;  //139 / 28 = 4
    16'b10001011_00011101 : OUT <= 4;  //139 / 29 = 4
    16'b10001011_00011110 : OUT <= 4;  //139 / 30 = 4
    16'b10001011_00011111 : OUT <= 4;  //139 / 31 = 4
    16'b10001011_00100000 : OUT <= 4;  //139 / 32 = 4
    16'b10001011_00100001 : OUT <= 4;  //139 / 33 = 4
    16'b10001011_00100010 : OUT <= 4;  //139 / 34 = 4
    16'b10001011_00100011 : OUT <= 3;  //139 / 35 = 3
    16'b10001011_00100100 : OUT <= 3;  //139 / 36 = 3
    16'b10001011_00100101 : OUT <= 3;  //139 / 37 = 3
    16'b10001011_00100110 : OUT <= 3;  //139 / 38 = 3
    16'b10001011_00100111 : OUT <= 3;  //139 / 39 = 3
    16'b10001011_00101000 : OUT <= 3;  //139 / 40 = 3
    16'b10001011_00101001 : OUT <= 3;  //139 / 41 = 3
    16'b10001011_00101010 : OUT <= 3;  //139 / 42 = 3
    16'b10001011_00101011 : OUT <= 3;  //139 / 43 = 3
    16'b10001011_00101100 : OUT <= 3;  //139 / 44 = 3
    16'b10001011_00101101 : OUT <= 3;  //139 / 45 = 3
    16'b10001011_00101110 : OUT <= 3;  //139 / 46 = 3
    16'b10001011_00101111 : OUT <= 2;  //139 / 47 = 2
    16'b10001011_00110000 : OUT <= 2;  //139 / 48 = 2
    16'b10001011_00110001 : OUT <= 2;  //139 / 49 = 2
    16'b10001011_00110010 : OUT <= 2;  //139 / 50 = 2
    16'b10001011_00110011 : OUT <= 2;  //139 / 51 = 2
    16'b10001011_00110100 : OUT <= 2;  //139 / 52 = 2
    16'b10001011_00110101 : OUT <= 2;  //139 / 53 = 2
    16'b10001011_00110110 : OUT <= 2;  //139 / 54 = 2
    16'b10001011_00110111 : OUT <= 2;  //139 / 55 = 2
    16'b10001011_00111000 : OUT <= 2;  //139 / 56 = 2
    16'b10001011_00111001 : OUT <= 2;  //139 / 57 = 2
    16'b10001011_00111010 : OUT <= 2;  //139 / 58 = 2
    16'b10001011_00111011 : OUT <= 2;  //139 / 59 = 2
    16'b10001011_00111100 : OUT <= 2;  //139 / 60 = 2
    16'b10001011_00111101 : OUT <= 2;  //139 / 61 = 2
    16'b10001011_00111110 : OUT <= 2;  //139 / 62 = 2
    16'b10001011_00111111 : OUT <= 2;  //139 / 63 = 2
    16'b10001011_01000000 : OUT <= 2;  //139 / 64 = 2
    16'b10001011_01000001 : OUT <= 2;  //139 / 65 = 2
    16'b10001011_01000010 : OUT <= 2;  //139 / 66 = 2
    16'b10001011_01000011 : OUT <= 2;  //139 / 67 = 2
    16'b10001011_01000100 : OUT <= 2;  //139 / 68 = 2
    16'b10001011_01000101 : OUT <= 2;  //139 / 69 = 2
    16'b10001011_01000110 : OUT <= 1;  //139 / 70 = 1
    16'b10001011_01000111 : OUT <= 1;  //139 / 71 = 1
    16'b10001011_01001000 : OUT <= 1;  //139 / 72 = 1
    16'b10001011_01001001 : OUT <= 1;  //139 / 73 = 1
    16'b10001011_01001010 : OUT <= 1;  //139 / 74 = 1
    16'b10001011_01001011 : OUT <= 1;  //139 / 75 = 1
    16'b10001011_01001100 : OUT <= 1;  //139 / 76 = 1
    16'b10001011_01001101 : OUT <= 1;  //139 / 77 = 1
    16'b10001011_01001110 : OUT <= 1;  //139 / 78 = 1
    16'b10001011_01001111 : OUT <= 1;  //139 / 79 = 1
    16'b10001011_01010000 : OUT <= 1;  //139 / 80 = 1
    16'b10001011_01010001 : OUT <= 1;  //139 / 81 = 1
    16'b10001011_01010010 : OUT <= 1;  //139 / 82 = 1
    16'b10001011_01010011 : OUT <= 1;  //139 / 83 = 1
    16'b10001011_01010100 : OUT <= 1;  //139 / 84 = 1
    16'b10001011_01010101 : OUT <= 1;  //139 / 85 = 1
    16'b10001011_01010110 : OUT <= 1;  //139 / 86 = 1
    16'b10001011_01010111 : OUT <= 1;  //139 / 87 = 1
    16'b10001011_01011000 : OUT <= 1;  //139 / 88 = 1
    16'b10001011_01011001 : OUT <= 1;  //139 / 89 = 1
    16'b10001011_01011010 : OUT <= 1;  //139 / 90 = 1
    16'b10001011_01011011 : OUT <= 1;  //139 / 91 = 1
    16'b10001011_01011100 : OUT <= 1;  //139 / 92 = 1
    16'b10001011_01011101 : OUT <= 1;  //139 / 93 = 1
    16'b10001011_01011110 : OUT <= 1;  //139 / 94 = 1
    16'b10001011_01011111 : OUT <= 1;  //139 / 95 = 1
    16'b10001011_01100000 : OUT <= 1;  //139 / 96 = 1
    16'b10001011_01100001 : OUT <= 1;  //139 / 97 = 1
    16'b10001011_01100010 : OUT <= 1;  //139 / 98 = 1
    16'b10001011_01100011 : OUT <= 1;  //139 / 99 = 1
    16'b10001011_01100100 : OUT <= 1;  //139 / 100 = 1
    16'b10001011_01100101 : OUT <= 1;  //139 / 101 = 1
    16'b10001011_01100110 : OUT <= 1;  //139 / 102 = 1
    16'b10001011_01100111 : OUT <= 1;  //139 / 103 = 1
    16'b10001011_01101000 : OUT <= 1;  //139 / 104 = 1
    16'b10001011_01101001 : OUT <= 1;  //139 / 105 = 1
    16'b10001011_01101010 : OUT <= 1;  //139 / 106 = 1
    16'b10001011_01101011 : OUT <= 1;  //139 / 107 = 1
    16'b10001011_01101100 : OUT <= 1;  //139 / 108 = 1
    16'b10001011_01101101 : OUT <= 1;  //139 / 109 = 1
    16'b10001011_01101110 : OUT <= 1;  //139 / 110 = 1
    16'b10001011_01101111 : OUT <= 1;  //139 / 111 = 1
    16'b10001011_01110000 : OUT <= 1;  //139 / 112 = 1
    16'b10001011_01110001 : OUT <= 1;  //139 / 113 = 1
    16'b10001011_01110010 : OUT <= 1;  //139 / 114 = 1
    16'b10001011_01110011 : OUT <= 1;  //139 / 115 = 1
    16'b10001011_01110100 : OUT <= 1;  //139 / 116 = 1
    16'b10001011_01110101 : OUT <= 1;  //139 / 117 = 1
    16'b10001011_01110110 : OUT <= 1;  //139 / 118 = 1
    16'b10001011_01110111 : OUT <= 1;  //139 / 119 = 1
    16'b10001011_01111000 : OUT <= 1;  //139 / 120 = 1
    16'b10001011_01111001 : OUT <= 1;  //139 / 121 = 1
    16'b10001011_01111010 : OUT <= 1;  //139 / 122 = 1
    16'b10001011_01111011 : OUT <= 1;  //139 / 123 = 1
    16'b10001011_01111100 : OUT <= 1;  //139 / 124 = 1
    16'b10001011_01111101 : OUT <= 1;  //139 / 125 = 1
    16'b10001011_01111110 : OUT <= 1;  //139 / 126 = 1
    16'b10001011_01111111 : OUT <= 1;  //139 / 127 = 1
    16'b10001011_10000000 : OUT <= 1;  //139 / 128 = 1
    16'b10001011_10000001 : OUT <= 1;  //139 / 129 = 1
    16'b10001011_10000010 : OUT <= 1;  //139 / 130 = 1
    16'b10001011_10000011 : OUT <= 1;  //139 / 131 = 1
    16'b10001011_10000100 : OUT <= 1;  //139 / 132 = 1
    16'b10001011_10000101 : OUT <= 1;  //139 / 133 = 1
    16'b10001011_10000110 : OUT <= 1;  //139 / 134 = 1
    16'b10001011_10000111 : OUT <= 1;  //139 / 135 = 1
    16'b10001011_10001000 : OUT <= 1;  //139 / 136 = 1
    16'b10001011_10001001 : OUT <= 1;  //139 / 137 = 1
    16'b10001011_10001010 : OUT <= 1;  //139 / 138 = 1
    16'b10001011_10001011 : OUT <= 1;  //139 / 139 = 1
    16'b10001011_10001100 : OUT <= 0;  //139 / 140 = 0
    16'b10001011_10001101 : OUT <= 0;  //139 / 141 = 0
    16'b10001011_10001110 : OUT <= 0;  //139 / 142 = 0
    16'b10001011_10001111 : OUT <= 0;  //139 / 143 = 0
    16'b10001011_10010000 : OUT <= 0;  //139 / 144 = 0
    16'b10001011_10010001 : OUT <= 0;  //139 / 145 = 0
    16'b10001011_10010010 : OUT <= 0;  //139 / 146 = 0
    16'b10001011_10010011 : OUT <= 0;  //139 / 147 = 0
    16'b10001011_10010100 : OUT <= 0;  //139 / 148 = 0
    16'b10001011_10010101 : OUT <= 0;  //139 / 149 = 0
    16'b10001011_10010110 : OUT <= 0;  //139 / 150 = 0
    16'b10001011_10010111 : OUT <= 0;  //139 / 151 = 0
    16'b10001011_10011000 : OUT <= 0;  //139 / 152 = 0
    16'b10001011_10011001 : OUT <= 0;  //139 / 153 = 0
    16'b10001011_10011010 : OUT <= 0;  //139 / 154 = 0
    16'b10001011_10011011 : OUT <= 0;  //139 / 155 = 0
    16'b10001011_10011100 : OUT <= 0;  //139 / 156 = 0
    16'b10001011_10011101 : OUT <= 0;  //139 / 157 = 0
    16'b10001011_10011110 : OUT <= 0;  //139 / 158 = 0
    16'b10001011_10011111 : OUT <= 0;  //139 / 159 = 0
    16'b10001011_10100000 : OUT <= 0;  //139 / 160 = 0
    16'b10001011_10100001 : OUT <= 0;  //139 / 161 = 0
    16'b10001011_10100010 : OUT <= 0;  //139 / 162 = 0
    16'b10001011_10100011 : OUT <= 0;  //139 / 163 = 0
    16'b10001011_10100100 : OUT <= 0;  //139 / 164 = 0
    16'b10001011_10100101 : OUT <= 0;  //139 / 165 = 0
    16'b10001011_10100110 : OUT <= 0;  //139 / 166 = 0
    16'b10001011_10100111 : OUT <= 0;  //139 / 167 = 0
    16'b10001011_10101000 : OUT <= 0;  //139 / 168 = 0
    16'b10001011_10101001 : OUT <= 0;  //139 / 169 = 0
    16'b10001011_10101010 : OUT <= 0;  //139 / 170 = 0
    16'b10001011_10101011 : OUT <= 0;  //139 / 171 = 0
    16'b10001011_10101100 : OUT <= 0;  //139 / 172 = 0
    16'b10001011_10101101 : OUT <= 0;  //139 / 173 = 0
    16'b10001011_10101110 : OUT <= 0;  //139 / 174 = 0
    16'b10001011_10101111 : OUT <= 0;  //139 / 175 = 0
    16'b10001011_10110000 : OUT <= 0;  //139 / 176 = 0
    16'b10001011_10110001 : OUT <= 0;  //139 / 177 = 0
    16'b10001011_10110010 : OUT <= 0;  //139 / 178 = 0
    16'b10001011_10110011 : OUT <= 0;  //139 / 179 = 0
    16'b10001011_10110100 : OUT <= 0;  //139 / 180 = 0
    16'b10001011_10110101 : OUT <= 0;  //139 / 181 = 0
    16'b10001011_10110110 : OUT <= 0;  //139 / 182 = 0
    16'b10001011_10110111 : OUT <= 0;  //139 / 183 = 0
    16'b10001011_10111000 : OUT <= 0;  //139 / 184 = 0
    16'b10001011_10111001 : OUT <= 0;  //139 / 185 = 0
    16'b10001011_10111010 : OUT <= 0;  //139 / 186 = 0
    16'b10001011_10111011 : OUT <= 0;  //139 / 187 = 0
    16'b10001011_10111100 : OUT <= 0;  //139 / 188 = 0
    16'b10001011_10111101 : OUT <= 0;  //139 / 189 = 0
    16'b10001011_10111110 : OUT <= 0;  //139 / 190 = 0
    16'b10001011_10111111 : OUT <= 0;  //139 / 191 = 0
    16'b10001011_11000000 : OUT <= 0;  //139 / 192 = 0
    16'b10001011_11000001 : OUT <= 0;  //139 / 193 = 0
    16'b10001011_11000010 : OUT <= 0;  //139 / 194 = 0
    16'b10001011_11000011 : OUT <= 0;  //139 / 195 = 0
    16'b10001011_11000100 : OUT <= 0;  //139 / 196 = 0
    16'b10001011_11000101 : OUT <= 0;  //139 / 197 = 0
    16'b10001011_11000110 : OUT <= 0;  //139 / 198 = 0
    16'b10001011_11000111 : OUT <= 0;  //139 / 199 = 0
    16'b10001011_11001000 : OUT <= 0;  //139 / 200 = 0
    16'b10001011_11001001 : OUT <= 0;  //139 / 201 = 0
    16'b10001011_11001010 : OUT <= 0;  //139 / 202 = 0
    16'b10001011_11001011 : OUT <= 0;  //139 / 203 = 0
    16'b10001011_11001100 : OUT <= 0;  //139 / 204 = 0
    16'b10001011_11001101 : OUT <= 0;  //139 / 205 = 0
    16'b10001011_11001110 : OUT <= 0;  //139 / 206 = 0
    16'b10001011_11001111 : OUT <= 0;  //139 / 207 = 0
    16'b10001011_11010000 : OUT <= 0;  //139 / 208 = 0
    16'b10001011_11010001 : OUT <= 0;  //139 / 209 = 0
    16'b10001011_11010010 : OUT <= 0;  //139 / 210 = 0
    16'b10001011_11010011 : OUT <= 0;  //139 / 211 = 0
    16'b10001011_11010100 : OUT <= 0;  //139 / 212 = 0
    16'b10001011_11010101 : OUT <= 0;  //139 / 213 = 0
    16'b10001011_11010110 : OUT <= 0;  //139 / 214 = 0
    16'b10001011_11010111 : OUT <= 0;  //139 / 215 = 0
    16'b10001011_11011000 : OUT <= 0;  //139 / 216 = 0
    16'b10001011_11011001 : OUT <= 0;  //139 / 217 = 0
    16'b10001011_11011010 : OUT <= 0;  //139 / 218 = 0
    16'b10001011_11011011 : OUT <= 0;  //139 / 219 = 0
    16'b10001011_11011100 : OUT <= 0;  //139 / 220 = 0
    16'b10001011_11011101 : OUT <= 0;  //139 / 221 = 0
    16'b10001011_11011110 : OUT <= 0;  //139 / 222 = 0
    16'b10001011_11011111 : OUT <= 0;  //139 / 223 = 0
    16'b10001011_11100000 : OUT <= 0;  //139 / 224 = 0
    16'b10001011_11100001 : OUT <= 0;  //139 / 225 = 0
    16'b10001011_11100010 : OUT <= 0;  //139 / 226 = 0
    16'b10001011_11100011 : OUT <= 0;  //139 / 227 = 0
    16'b10001011_11100100 : OUT <= 0;  //139 / 228 = 0
    16'b10001011_11100101 : OUT <= 0;  //139 / 229 = 0
    16'b10001011_11100110 : OUT <= 0;  //139 / 230 = 0
    16'b10001011_11100111 : OUT <= 0;  //139 / 231 = 0
    16'b10001011_11101000 : OUT <= 0;  //139 / 232 = 0
    16'b10001011_11101001 : OUT <= 0;  //139 / 233 = 0
    16'b10001011_11101010 : OUT <= 0;  //139 / 234 = 0
    16'b10001011_11101011 : OUT <= 0;  //139 / 235 = 0
    16'b10001011_11101100 : OUT <= 0;  //139 / 236 = 0
    16'b10001011_11101101 : OUT <= 0;  //139 / 237 = 0
    16'b10001011_11101110 : OUT <= 0;  //139 / 238 = 0
    16'b10001011_11101111 : OUT <= 0;  //139 / 239 = 0
    16'b10001011_11110000 : OUT <= 0;  //139 / 240 = 0
    16'b10001011_11110001 : OUT <= 0;  //139 / 241 = 0
    16'b10001011_11110010 : OUT <= 0;  //139 / 242 = 0
    16'b10001011_11110011 : OUT <= 0;  //139 / 243 = 0
    16'b10001011_11110100 : OUT <= 0;  //139 / 244 = 0
    16'b10001011_11110101 : OUT <= 0;  //139 / 245 = 0
    16'b10001011_11110110 : OUT <= 0;  //139 / 246 = 0
    16'b10001011_11110111 : OUT <= 0;  //139 / 247 = 0
    16'b10001011_11111000 : OUT <= 0;  //139 / 248 = 0
    16'b10001011_11111001 : OUT <= 0;  //139 / 249 = 0
    16'b10001011_11111010 : OUT <= 0;  //139 / 250 = 0
    16'b10001011_11111011 : OUT <= 0;  //139 / 251 = 0
    16'b10001011_11111100 : OUT <= 0;  //139 / 252 = 0
    16'b10001011_11111101 : OUT <= 0;  //139 / 253 = 0
    16'b10001011_11111110 : OUT <= 0;  //139 / 254 = 0
    16'b10001011_11111111 : OUT <= 0;  //139 / 255 = 0
    16'b10001100_00000000 : OUT <= 0;  //140 / 0 = 0
    16'b10001100_00000001 : OUT <= 140;  //140 / 1 = 140
    16'b10001100_00000010 : OUT <= 70;  //140 / 2 = 70
    16'b10001100_00000011 : OUT <= 46;  //140 / 3 = 46
    16'b10001100_00000100 : OUT <= 35;  //140 / 4 = 35
    16'b10001100_00000101 : OUT <= 28;  //140 / 5 = 28
    16'b10001100_00000110 : OUT <= 23;  //140 / 6 = 23
    16'b10001100_00000111 : OUT <= 20;  //140 / 7 = 20
    16'b10001100_00001000 : OUT <= 17;  //140 / 8 = 17
    16'b10001100_00001001 : OUT <= 15;  //140 / 9 = 15
    16'b10001100_00001010 : OUT <= 14;  //140 / 10 = 14
    16'b10001100_00001011 : OUT <= 12;  //140 / 11 = 12
    16'b10001100_00001100 : OUT <= 11;  //140 / 12 = 11
    16'b10001100_00001101 : OUT <= 10;  //140 / 13 = 10
    16'b10001100_00001110 : OUT <= 10;  //140 / 14 = 10
    16'b10001100_00001111 : OUT <= 9;  //140 / 15 = 9
    16'b10001100_00010000 : OUT <= 8;  //140 / 16 = 8
    16'b10001100_00010001 : OUT <= 8;  //140 / 17 = 8
    16'b10001100_00010010 : OUT <= 7;  //140 / 18 = 7
    16'b10001100_00010011 : OUT <= 7;  //140 / 19 = 7
    16'b10001100_00010100 : OUT <= 7;  //140 / 20 = 7
    16'b10001100_00010101 : OUT <= 6;  //140 / 21 = 6
    16'b10001100_00010110 : OUT <= 6;  //140 / 22 = 6
    16'b10001100_00010111 : OUT <= 6;  //140 / 23 = 6
    16'b10001100_00011000 : OUT <= 5;  //140 / 24 = 5
    16'b10001100_00011001 : OUT <= 5;  //140 / 25 = 5
    16'b10001100_00011010 : OUT <= 5;  //140 / 26 = 5
    16'b10001100_00011011 : OUT <= 5;  //140 / 27 = 5
    16'b10001100_00011100 : OUT <= 5;  //140 / 28 = 5
    16'b10001100_00011101 : OUT <= 4;  //140 / 29 = 4
    16'b10001100_00011110 : OUT <= 4;  //140 / 30 = 4
    16'b10001100_00011111 : OUT <= 4;  //140 / 31 = 4
    16'b10001100_00100000 : OUT <= 4;  //140 / 32 = 4
    16'b10001100_00100001 : OUT <= 4;  //140 / 33 = 4
    16'b10001100_00100010 : OUT <= 4;  //140 / 34 = 4
    16'b10001100_00100011 : OUT <= 4;  //140 / 35 = 4
    16'b10001100_00100100 : OUT <= 3;  //140 / 36 = 3
    16'b10001100_00100101 : OUT <= 3;  //140 / 37 = 3
    16'b10001100_00100110 : OUT <= 3;  //140 / 38 = 3
    16'b10001100_00100111 : OUT <= 3;  //140 / 39 = 3
    16'b10001100_00101000 : OUT <= 3;  //140 / 40 = 3
    16'b10001100_00101001 : OUT <= 3;  //140 / 41 = 3
    16'b10001100_00101010 : OUT <= 3;  //140 / 42 = 3
    16'b10001100_00101011 : OUT <= 3;  //140 / 43 = 3
    16'b10001100_00101100 : OUT <= 3;  //140 / 44 = 3
    16'b10001100_00101101 : OUT <= 3;  //140 / 45 = 3
    16'b10001100_00101110 : OUT <= 3;  //140 / 46 = 3
    16'b10001100_00101111 : OUT <= 2;  //140 / 47 = 2
    16'b10001100_00110000 : OUT <= 2;  //140 / 48 = 2
    16'b10001100_00110001 : OUT <= 2;  //140 / 49 = 2
    16'b10001100_00110010 : OUT <= 2;  //140 / 50 = 2
    16'b10001100_00110011 : OUT <= 2;  //140 / 51 = 2
    16'b10001100_00110100 : OUT <= 2;  //140 / 52 = 2
    16'b10001100_00110101 : OUT <= 2;  //140 / 53 = 2
    16'b10001100_00110110 : OUT <= 2;  //140 / 54 = 2
    16'b10001100_00110111 : OUT <= 2;  //140 / 55 = 2
    16'b10001100_00111000 : OUT <= 2;  //140 / 56 = 2
    16'b10001100_00111001 : OUT <= 2;  //140 / 57 = 2
    16'b10001100_00111010 : OUT <= 2;  //140 / 58 = 2
    16'b10001100_00111011 : OUT <= 2;  //140 / 59 = 2
    16'b10001100_00111100 : OUT <= 2;  //140 / 60 = 2
    16'b10001100_00111101 : OUT <= 2;  //140 / 61 = 2
    16'b10001100_00111110 : OUT <= 2;  //140 / 62 = 2
    16'b10001100_00111111 : OUT <= 2;  //140 / 63 = 2
    16'b10001100_01000000 : OUT <= 2;  //140 / 64 = 2
    16'b10001100_01000001 : OUT <= 2;  //140 / 65 = 2
    16'b10001100_01000010 : OUT <= 2;  //140 / 66 = 2
    16'b10001100_01000011 : OUT <= 2;  //140 / 67 = 2
    16'b10001100_01000100 : OUT <= 2;  //140 / 68 = 2
    16'b10001100_01000101 : OUT <= 2;  //140 / 69 = 2
    16'b10001100_01000110 : OUT <= 2;  //140 / 70 = 2
    16'b10001100_01000111 : OUT <= 1;  //140 / 71 = 1
    16'b10001100_01001000 : OUT <= 1;  //140 / 72 = 1
    16'b10001100_01001001 : OUT <= 1;  //140 / 73 = 1
    16'b10001100_01001010 : OUT <= 1;  //140 / 74 = 1
    16'b10001100_01001011 : OUT <= 1;  //140 / 75 = 1
    16'b10001100_01001100 : OUT <= 1;  //140 / 76 = 1
    16'b10001100_01001101 : OUT <= 1;  //140 / 77 = 1
    16'b10001100_01001110 : OUT <= 1;  //140 / 78 = 1
    16'b10001100_01001111 : OUT <= 1;  //140 / 79 = 1
    16'b10001100_01010000 : OUT <= 1;  //140 / 80 = 1
    16'b10001100_01010001 : OUT <= 1;  //140 / 81 = 1
    16'b10001100_01010010 : OUT <= 1;  //140 / 82 = 1
    16'b10001100_01010011 : OUT <= 1;  //140 / 83 = 1
    16'b10001100_01010100 : OUT <= 1;  //140 / 84 = 1
    16'b10001100_01010101 : OUT <= 1;  //140 / 85 = 1
    16'b10001100_01010110 : OUT <= 1;  //140 / 86 = 1
    16'b10001100_01010111 : OUT <= 1;  //140 / 87 = 1
    16'b10001100_01011000 : OUT <= 1;  //140 / 88 = 1
    16'b10001100_01011001 : OUT <= 1;  //140 / 89 = 1
    16'b10001100_01011010 : OUT <= 1;  //140 / 90 = 1
    16'b10001100_01011011 : OUT <= 1;  //140 / 91 = 1
    16'b10001100_01011100 : OUT <= 1;  //140 / 92 = 1
    16'b10001100_01011101 : OUT <= 1;  //140 / 93 = 1
    16'b10001100_01011110 : OUT <= 1;  //140 / 94 = 1
    16'b10001100_01011111 : OUT <= 1;  //140 / 95 = 1
    16'b10001100_01100000 : OUT <= 1;  //140 / 96 = 1
    16'b10001100_01100001 : OUT <= 1;  //140 / 97 = 1
    16'b10001100_01100010 : OUT <= 1;  //140 / 98 = 1
    16'b10001100_01100011 : OUT <= 1;  //140 / 99 = 1
    16'b10001100_01100100 : OUT <= 1;  //140 / 100 = 1
    16'b10001100_01100101 : OUT <= 1;  //140 / 101 = 1
    16'b10001100_01100110 : OUT <= 1;  //140 / 102 = 1
    16'b10001100_01100111 : OUT <= 1;  //140 / 103 = 1
    16'b10001100_01101000 : OUT <= 1;  //140 / 104 = 1
    16'b10001100_01101001 : OUT <= 1;  //140 / 105 = 1
    16'b10001100_01101010 : OUT <= 1;  //140 / 106 = 1
    16'b10001100_01101011 : OUT <= 1;  //140 / 107 = 1
    16'b10001100_01101100 : OUT <= 1;  //140 / 108 = 1
    16'b10001100_01101101 : OUT <= 1;  //140 / 109 = 1
    16'b10001100_01101110 : OUT <= 1;  //140 / 110 = 1
    16'b10001100_01101111 : OUT <= 1;  //140 / 111 = 1
    16'b10001100_01110000 : OUT <= 1;  //140 / 112 = 1
    16'b10001100_01110001 : OUT <= 1;  //140 / 113 = 1
    16'b10001100_01110010 : OUT <= 1;  //140 / 114 = 1
    16'b10001100_01110011 : OUT <= 1;  //140 / 115 = 1
    16'b10001100_01110100 : OUT <= 1;  //140 / 116 = 1
    16'b10001100_01110101 : OUT <= 1;  //140 / 117 = 1
    16'b10001100_01110110 : OUT <= 1;  //140 / 118 = 1
    16'b10001100_01110111 : OUT <= 1;  //140 / 119 = 1
    16'b10001100_01111000 : OUT <= 1;  //140 / 120 = 1
    16'b10001100_01111001 : OUT <= 1;  //140 / 121 = 1
    16'b10001100_01111010 : OUT <= 1;  //140 / 122 = 1
    16'b10001100_01111011 : OUT <= 1;  //140 / 123 = 1
    16'b10001100_01111100 : OUT <= 1;  //140 / 124 = 1
    16'b10001100_01111101 : OUT <= 1;  //140 / 125 = 1
    16'b10001100_01111110 : OUT <= 1;  //140 / 126 = 1
    16'b10001100_01111111 : OUT <= 1;  //140 / 127 = 1
    16'b10001100_10000000 : OUT <= 1;  //140 / 128 = 1
    16'b10001100_10000001 : OUT <= 1;  //140 / 129 = 1
    16'b10001100_10000010 : OUT <= 1;  //140 / 130 = 1
    16'b10001100_10000011 : OUT <= 1;  //140 / 131 = 1
    16'b10001100_10000100 : OUT <= 1;  //140 / 132 = 1
    16'b10001100_10000101 : OUT <= 1;  //140 / 133 = 1
    16'b10001100_10000110 : OUT <= 1;  //140 / 134 = 1
    16'b10001100_10000111 : OUT <= 1;  //140 / 135 = 1
    16'b10001100_10001000 : OUT <= 1;  //140 / 136 = 1
    16'b10001100_10001001 : OUT <= 1;  //140 / 137 = 1
    16'b10001100_10001010 : OUT <= 1;  //140 / 138 = 1
    16'b10001100_10001011 : OUT <= 1;  //140 / 139 = 1
    16'b10001100_10001100 : OUT <= 1;  //140 / 140 = 1
    16'b10001100_10001101 : OUT <= 0;  //140 / 141 = 0
    16'b10001100_10001110 : OUT <= 0;  //140 / 142 = 0
    16'b10001100_10001111 : OUT <= 0;  //140 / 143 = 0
    16'b10001100_10010000 : OUT <= 0;  //140 / 144 = 0
    16'b10001100_10010001 : OUT <= 0;  //140 / 145 = 0
    16'b10001100_10010010 : OUT <= 0;  //140 / 146 = 0
    16'b10001100_10010011 : OUT <= 0;  //140 / 147 = 0
    16'b10001100_10010100 : OUT <= 0;  //140 / 148 = 0
    16'b10001100_10010101 : OUT <= 0;  //140 / 149 = 0
    16'b10001100_10010110 : OUT <= 0;  //140 / 150 = 0
    16'b10001100_10010111 : OUT <= 0;  //140 / 151 = 0
    16'b10001100_10011000 : OUT <= 0;  //140 / 152 = 0
    16'b10001100_10011001 : OUT <= 0;  //140 / 153 = 0
    16'b10001100_10011010 : OUT <= 0;  //140 / 154 = 0
    16'b10001100_10011011 : OUT <= 0;  //140 / 155 = 0
    16'b10001100_10011100 : OUT <= 0;  //140 / 156 = 0
    16'b10001100_10011101 : OUT <= 0;  //140 / 157 = 0
    16'b10001100_10011110 : OUT <= 0;  //140 / 158 = 0
    16'b10001100_10011111 : OUT <= 0;  //140 / 159 = 0
    16'b10001100_10100000 : OUT <= 0;  //140 / 160 = 0
    16'b10001100_10100001 : OUT <= 0;  //140 / 161 = 0
    16'b10001100_10100010 : OUT <= 0;  //140 / 162 = 0
    16'b10001100_10100011 : OUT <= 0;  //140 / 163 = 0
    16'b10001100_10100100 : OUT <= 0;  //140 / 164 = 0
    16'b10001100_10100101 : OUT <= 0;  //140 / 165 = 0
    16'b10001100_10100110 : OUT <= 0;  //140 / 166 = 0
    16'b10001100_10100111 : OUT <= 0;  //140 / 167 = 0
    16'b10001100_10101000 : OUT <= 0;  //140 / 168 = 0
    16'b10001100_10101001 : OUT <= 0;  //140 / 169 = 0
    16'b10001100_10101010 : OUT <= 0;  //140 / 170 = 0
    16'b10001100_10101011 : OUT <= 0;  //140 / 171 = 0
    16'b10001100_10101100 : OUT <= 0;  //140 / 172 = 0
    16'b10001100_10101101 : OUT <= 0;  //140 / 173 = 0
    16'b10001100_10101110 : OUT <= 0;  //140 / 174 = 0
    16'b10001100_10101111 : OUT <= 0;  //140 / 175 = 0
    16'b10001100_10110000 : OUT <= 0;  //140 / 176 = 0
    16'b10001100_10110001 : OUT <= 0;  //140 / 177 = 0
    16'b10001100_10110010 : OUT <= 0;  //140 / 178 = 0
    16'b10001100_10110011 : OUT <= 0;  //140 / 179 = 0
    16'b10001100_10110100 : OUT <= 0;  //140 / 180 = 0
    16'b10001100_10110101 : OUT <= 0;  //140 / 181 = 0
    16'b10001100_10110110 : OUT <= 0;  //140 / 182 = 0
    16'b10001100_10110111 : OUT <= 0;  //140 / 183 = 0
    16'b10001100_10111000 : OUT <= 0;  //140 / 184 = 0
    16'b10001100_10111001 : OUT <= 0;  //140 / 185 = 0
    16'b10001100_10111010 : OUT <= 0;  //140 / 186 = 0
    16'b10001100_10111011 : OUT <= 0;  //140 / 187 = 0
    16'b10001100_10111100 : OUT <= 0;  //140 / 188 = 0
    16'b10001100_10111101 : OUT <= 0;  //140 / 189 = 0
    16'b10001100_10111110 : OUT <= 0;  //140 / 190 = 0
    16'b10001100_10111111 : OUT <= 0;  //140 / 191 = 0
    16'b10001100_11000000 : OUT <= 0;  //140 / 192 = 0
    16'b10001100_11000001 : OUT <= 0;  //140 / 193 = 0
    16'b10001100_11000010 : OUT <= 0;  //140 / 194 = 0
    16'b10001100_11000011 : OUT <= 0;  //140 / 195 = 0
    16'b10001100_11000100 : OUT <= 0;  //140 / 196 = 0
    16'b10001100_11000101 : OUT <= 0;  //140 / 197 = 0
    16'b10001100_11000110 : OUT <= 0;  //140 / 198 = 0
    16'b10001100_11000111 : OUT <= 0;  //140 / 199 = 0
    16'b10001100_11001000 : OUT <= 0;  //140 / 200 = 0
    16'b10001100_11001001 : OUT <= 0;  //140 / 201 = 0
    16'b10001100_11001010 : OUT <= 0;  //140 / 202 = 0
    16'b10001100_11001011 : OUT <= 0;  //140 / 203 = 0
    16'b10001100_11001100 : OUT <= 0;  //140 / 204 = 0
    16'b10001100_11001101 : OUT <= 0;  //140 / 205 = 0
    16'b10001100_11001110 : OUT <= 0;  //140 / 206 = 0
    16'b10001100_11001111 : OUT <= 0;  //140 / 207 = 0
    16'b10001100_11010000 : OUT <= 0;  //140 / 208 = 0
    16'b10001100_11010001 : OUT <= 0;  //140 / 209 = 0
    16'b10001100_11010010 : OUT <= 0;  //140 / 210 = 0
    16'b10001100_11010011 : OUT <= 0;  //140 / 211 = 0
    16'b10001100_11010100 : OUT <= 0;  //140 / 212 = 0
    16'b10001100_11010101 : OUT <= 0;  //140 / 213 = 0
    16'b10001100_11010110 : OUT <= 0;  //140 / 214 = 0
    16'b10001100_11010111 : OUT <= 0;  //140 / 215 = 0
    16'b10001100_11011000 : OUT <= 0;  //140 / 216 = 0
    16'b10001100_11011001 : OUT <= 0;  //140 / 217 = 0
    16'b10001100_11011010 : OUT <= 0;  //140 / 218 = 0
    16'b10001100_11011011 : OUT <= 0;  //140 / 219 = 0
    16'b10001100_11011100 : OUT <= 0;  //140 / 220 = 0
    16'b10001100_11011101 : OUT <= 0;  //140 / 221 = 0
    16'b10001100_11011110 : OUT <= 0;  //140 / 222 = 0
    16'b10001100_11011111 : OUT <= 0;  //140 / 223 = 0
    16'b10001100_11100000 : OUT <= 0;  //140 / 224 = 0
    16'b10001100_11100001 : OUT <= 0;  //140 / 225 = 0
    16'b10001100_11100010 : OUT <= 0;  //140 / 226 = 0
    16'b10001100_11100011 : OUT <= 0;  //140 / 227 = 0
    16'b10001100_11100100 : OUT <= 0;  //140 / 228 = 0
    16'b10001100_11100101 : OUT <= 0;  //140 / 229 = 0
    16'b10001100_11100110 : OUT <= 0;  //140 / 230 = 0
    16'b10001100_11100111 : OUT <= 0;  //140 / 231 = 0
    16'b10001100_11101000 : OUT <= 0;  //140 / 232 = 0
    16'b10001100_11101001 : OUT <= 0;  //140 / 233 = 0
    16'b10001100_11101010 : OUT <= 0;  //140 / 234 = 0
    16'b10001100_11101011 : OUT <= 0;  //140 / 235 = 0
    16'b10001100_11101100 : OUT <= 0;  //140 / 236 = 0
    16'b10001100_11101101 : OUT <= 0;  //140 / 237 = 0
    16'b10001100_11101110 : OUT <= 0;  //140 / 238 = 0
    16'b10001100_11101111 : OUT <= 0;  //140 / 239 = 0
    16'b10001100_11110000 : OUT <= 0;  //140 / 240 = 0
    16'b10001100_11110001 : OUT <= 0;  //140 / 241 = 0
    16'b10001100_11110010 : OUT <= 0;  //140 / 242 = 0
    16'b10001100_11110011 : OUT <= 0;  //140 / 243 = 0
    16'b10001100_11110100 : OUT <= 0;  //140 / 244 = 0
    16'b10001100_11110101 : OUT <= 0;  //140 / 245 = 0
    16'b10001100_11110110 : OUT <= 0;  //140 / 246 = 0
    16'b10001100_11110111 : OUT <= 0;  //140 / 247 = 0
    16'b10001100_11111000 : OUT <= 0;  //140 / 248 = 0
    16'b10001100_11111001 : OUT <= 0;  //140 / 249 = 0
    16'b10001100_11111010 : OUT <= 0;  //140 / 250 = 0
    16'b10001100_11111011 : OUT <= 0;  //140 / 251 = 0
    16'b10001100_11111100 : OUT <= 0;  //140 / 252 = 0
    16'b10001100_11111101 : OUT <= 0;  //140 / 253 = 0
    16'b10001100_11111110 : OUT <= 0;  //140 / 254 = 0
    16'b10001100_11111111 : OUT <= 0;  //140 / 255 = 0
    16'b10001101_00000000 : OUT <= 0;  //141 / 0 = 0
    16'b10001101_00000001 : OUT <= 141;  //141 / 1 = 141
    16'b10001101_00000010 : OUT <= 70;  //141 / 2 = 70
    16'b10001101_00000011 : OUT <= 47;  //141 / 3 = 47
    16'b10001101_00000100 : OUT <= 35;  //141 / 4 = 35
    16'b10001101_00000101 : OUT <= 28;  //141 / 5 = 28
    16'b10001101_00000110 : OUT <= 23;  //141 / 6 = 23
    16'b10001101_00000111 : OUT <= 20;  //141 / 7 = 20
    16'b10001101_00001000 : OUT <= 17;  //141 / 8 = 17
    16'b10001101_00001001 : OUT <= 15;  //141 / 9 = 15
    16'b10001101_00001010 : OUT <= 14;  //141 / 10 = 14
    16'b10001101_00001011 : OUT <= 12;  //141 / 11 = 12
    16'b10001101_00001100 : OUT <= 11;  //141 / 12 = 11
    16'b10001101_00001101 : OUT <= 10;  //141 / 13 = 10
    16'b10001101_00001110 : OUT <= 10;  //141 / 14 = 10
    16'b10001101_00001111 : OUT <= 9;  //141 / 15 = 9
    16'b10001101_00010000 : OUT <= 8;  //141 / 16 = 8
    16'b10001101_00010001 : OUT <= 8;  //141 / 17 = 8
    16'b10001101_00010010 : OUT <= 7;  //141 / 18 = 7
    16'b10001101_00010011 : OUT <= 7;  //141 / 19 = 7
    16'b10001101_00010100 : OUT <= 7;  //141 / 20 = 7
    16'b10001101_00010101 : OUT <= 6;  //141 / 21 = 6
    16'b10001101_00010110 : OUT <= 6;  //141 / 22 = 6
    16'b10001101_00010111 : OUT <= 6;  //141 / 23 = 6
    16'b10001101_00011000 : OUT <= 5;  //141 / 24 = 5
    16'b10001101_00011001 : OUT <= 5;  //141 / 25 = 5
    16'b10001101_00011010 : OUT <= 5;  //141 / 26 = 5
    16'b10001101_00011011 : OUT <= 5;  //141 / 27 = 5
    16'b10001101_00011100 : OUT <= 5;  //141 / 28 = 5
    16'b10001101_00011101 : OUT <= 4;  //141 / 29 = 4
    16'b10001101_00011110 : OUT <= 4;  //141 / 30 = 4
    16'b10001101_00011111 : OUT <= 4;  //141 / 31 = 4
    16'b10001101_00100000 : OUT <= 4;  //141 / 32 = 4
    16'b10001101_00100001 : OUT <= 4;  //141 / 33 = 4
    16'b10001101_00100010 : OUT <= 4;  //141 / 34 = 4
    16'b10001101_00100011 : OUT <= 4;  //141 / 35 = 4
    16'b10001101_00100100 : OUT <= 3;  //141 / 36 = 3
    16'b10001101_00100101 : OUT <= 3;  //141 / 37 = 3
    16'b10001101_00100110 : OUT <= 3;  //141 / 38 = 3
    16'b10001101_00100111 : OUT <= 3;  //141 / 39 = 3
    16'b10001101_00101000 : OUT <= 3;  //141 / 40 = 3
    16'b10001101_00101001 : OUT <= 3;  //141 / 41 = 3
    16'b10001101_00101010 : OUT <= 3;  //141 / 42 = 3
    16'b10001101_00101011 : OUT <= 3;  //141 / 43 = 3
    16'b10001101_00101100 : OUT <= 3;  //141 / 44 = 3
    16'b10001101_00101101 : OUT <= 3;  //141 / 45 = 3
    16'b10001101_00101110 : OUT <= 3;  //141 / 46 = 3
    16'b10001101_00101111 : OUT <= 3;  //141 / 47 = 3
    16'b10001101_00110000 : OUT <= 2;  //141 / 48 = 2
    16'b10001101_00110001 : OUT <= 2;  //141 / 49 = 2
    16'b10001101_00110010 : OUT <= 2;  //141 / 50 = 2
    16'b10001101_00110011 : OUT <= 2;  //141 / 51 = 2
    16'b10001101_00110100 : OUT <= 2;  //141 / 52 = 2
    16'b10001101_00110101 : OUT <= 2;  //141 / 53 = 2
    16'b10001101_00110110 : OUT <= 2;  //141 / 54 = 2
    16'b10001101_00110111 : OUT <= 2;  //141 / 55 = 2
    16'b10001101_00111000 : OUT <= 2;  //141 / 56 = 2
    16'b10001101_00111001 : OUT <= 2;  //141 / 57 = 2
    16'b10001101_00111010 : OUT <= 2;  //141 / 58 = 2
    16'b10001101_00111011 : OUT <= 2;  //141 / 59 = 2
    16'b10001101_00111100 : OUT <= 2;  //141 / 60 = 2
    16'b10001101_00111101 : OUT <= 2;  //141 / 61 = 2
    16'b10001101_00111110 : OUT <= 2;  //141 / 62 = 2
    16'b10001101_00111111 : OUT <= 2;  //141 / 63 = 2
    16'b10001101_01000000 : OUT <= 2;  //141 / 64 = 2
    16'b10001101_01000001 : OUT <= 2;  //141 / 65 = 2
    16'b10001101_01000010 : OUT <= 2;  //141 / 66 = 2
    16'b10001101_01000011 : OUT <= 2;  //141 / 67 = 2
    16'b10001101_01000100 : OUT <= 2;  //141 / 68 = 2
    16'b10001101_01000101 : OUT <= 2;  //141 / 69 = 2
    16'b10001101_01000110 : OUT <= 2;  //141 / 70 = 2
    16'b10001101_01000111 : OUT <= 1;  //141 / 71 = 1
    16'b10001101_01001000 : OUT <= 1;  //141 / 72 = 1
    16'b10001101_01001001 : OUT <= 1;  //141 / 73 = 1
    16'b10001101_01001010 : OUT <= 1;  //141 / 74 = 1
    16'b10001101_01001011 : OUT <= 1;  //141 / 75 = 1
    16'b10001101_01001100 : OUT <= 1;  //141 / 76 = 1
    16'b10001101_01001101 : OUT <= 1;  //141 / 77 = 1
    16'b10001101_01001110 : OUT <= 1;  //141 / 78 = 1
    16'b10001101_01001111 : OUT <= 1;  //141 / 79 = 1
    16'b10001101_01010000 : OUT <= 1;  //141 / 80 = 1
    16'b10001101_01010001 : OUT <= 1;  //141 / 81 = 1
    16'b10001101_01010010 : OUT <= 1;  //141 / 82 = 1
    16'b10001101_01010011 : OUT <= 1;  //141 / 83 = 1
    16'b10001101_01010100 : OUT <= 1;  //141 / 84 = 1
    16'b10001101_01010101 : OUT <= 1;  //141 / 85 = 1
    16'b10001101_01010110 : OUT <= 1;  //141 / 86 = 1
    16'b10001101_01010111 : OUT <= 1;  //141 / 87 = 1
    16'b10001101_01011000 : OUT <= 1;  //141 / 88 = 1
    16'b10001101_01011001 : OUT <= 1;  //141 / 89 = 1
    16'b10001101_01011010 : OUT <= 1;  //141 / 90 = 1
    16'b10001101_01011011 : OUT <= 1;  //141 / 91 = 1
    16'b10001101_01011100 : OUT <= 1;  //141 / 92 = 1
    16'b10001101_01011101 : OUT <= 1;  //141 / 93 = 1
    16'b10001101_01011110 : OUT <= 1;  //141 / 94 = 1
    16'b10001101_01011111 : OUT <= 1;  //141 / 95 = 1
    16'b10001101_01100000 : OUT <= 1;  //141 / 96 = 1
    16'b10001101_01100001 : OUT <= 1;  //141 / 97 = 1
    16'b10001101_01100010 : OUT <= 1;  //141 / 98 = 1
    16'b10001101_01100011 : OUT <= 1;  //141 / 99 = 1
    16'b10001101_01100100 : OUT <= 1;  //141 / 100 = 1
    16'b10001101_01100101 : OUT <= 1;  //141 / 101 = 1
    16'b10001101_01100110 : OUT <= 1;  //141 / 102 = 1
    16'b10001101_01100111 : OUT <= 1;  //141 / 103 = 1
    16'b10001101_01101000 : OUT <= 1;  //141 / 104 = 1
    16'b10001101_01101001 : OUT <= 1;  //141 / 105 = 1
    16'b10001101_01101010 : OUT <= 1;  //141 / 106 = 1
    16'b10001101_01101011 : OUT <= 1;  //141 / 107 = 1
    16'b10001101_01101100 : OUT <= 1;  //141 / 108 = 1
    16'b10001101_01101101 : OUT <= 1;  //141 / 109 = 1
    16'b10001101_01101110 : OUT <= 1;  //141 / 110 = 1
    16'b10001101_01101111 : OUT <= 1;  //141 / 111 = 1
    16'b10001101_01110000 : OUT <= 1;  //141 / 112 = 1
    16'b10001101_01110001 : OUT <= 1;  //141 / 113 = 1
    16'b10001101_01110010 : OUT <= 1;  //141 / 114 = 1
    16'b10001101_01110011 : OUT <= 1;  //141 / 115 = 1
    16'b10001101_01110100 : OUT <= 1;  //141 / 116 = 1
    16'b10001101_01110101 : OUT <= 1;  //141 / 117 = 1
    16'b10001101_01110110 : OUT <= 1;  //141 / 118 = 1
    16'b10001101_01110111 : OUT <= 1;  //141 / 119 = 1
    16'b10001101_01111000 : OUT <= 1;  //141 / 120 = 1
    16'b10001101_01111001 : OUT <= 1;  //141 / 121 = 1
    16'b10001101_01111010 : OUT <= 1;  //141 / 122 = 1
    16'b10001101_01111011 : OUT <= 1;  //141 / 123 = 1
    16'b10001101_01111100 : OUT <= 1;  //141 / 124 = 1
    16'b10001101_01111101 : OUT <= 1;  //141 / 125 = 1
    16'b10001101_01111110 : OUT <= 1;  //141 / 126 = 1
    16'b10001101_01111111 : OUT <= 1;  //141 / 127 = 1
    16'b10001101_10000000 : OUT <= 1;  //141 / 128 = 1
    16'b10001101_10000001 : OUT <= 1;  //141 / 129 = 1
    16'b10001101_10000010 : OUT <= 1;  //141 / 130 = 1
    16'b10001101_10000011 : OUT <= 1;  //141 / 131 = 1
    16'b10001101_10000100 : OUT <= 1;  //141 / 132 = 1
    16'b10001101_10000101 : OUT <= 1;  //141 / 133 = 1
    16'b10001101_10000110 : OUT <= 1;  //141 / 134 = 1
    16'b10001101_10000111 : OUT <= 1;  //141 / 135 = 1
    16'b10001101_10001000 : OUT <= 1;  //141 / 136 = 1
    16'b10001101_10001001 : OUT <= 1;  //141 / 137 = 1
    16'b10001101_10001010 : OUT <= 1;  //141 / 138 = 1
    16'b10001101_10001011 : OUT <= 1;  //141 / 139 = 1
    16'b10001101_10001100 : OUT <= 1;  //141 / 140 = 1
    16'b10001101_10001101 : OUT <= 1;  //141 / 141 = 1
    16'b10001101_10001110 : OUT <= 0;  //141 / 142 = 0
    16'b10001101_10001111 : OUT <= 0;  //141 / 143 = 0
    16'b10001101_10010000 : OUT <= 0;  //141 / 144 = 0
    16'b10001101_10010001 : OUT <= 0;  //141 / 145 = 0
    16'b10001101_10010010 : OUT <= 0;  //141 / 146 = 0
    16'b10001101_10010011 : OUT <= 0;  //141 / 147 = 0
    16'b10001101_10010100 : OUT <= 0;  //141 / 148 = 0
    16'b10001101_10010101 : OUT <= 0;  //141 / 149 = 0
    16'b10001101_10010110 : OUT <= 0;  //141 / 150 = 0
    16'b10001101_10010111 : OUT <= 0;  //141 / 151 = 0
    16'b10001101_10011000 : OUT <= 0;  //141 / 152 = 0
    16'b10001101_10011001 : OUT <= 0;  //141 / 153 = 0
    16'b10001101_10011010 : OUT <= 0;  //141 / 154 = 0
    16'b10001101_10011011 : OUT <= 0;  //141 / 155 = 0
    16'b10001101_10011100 : OUT <= 0;  //141 / 156 = 0
    16'b10001101_10011101 : OUT <= 0;  //141 / 157 = 0
    16'b10001101_10011110 : OUT <= 0;  //141 / 158 = 0
    16'b10001101_10011111 : OUT <= 0;  //141 / 159 = 0
    16'b10001101_10100000 : OUT <= 0;  //141 / 160 = 0
    16'b10001101_10100001 : OUT <= 0;  //141 / 161 = 0
    16'b10001101_10100010 : OUT <= 0;  //141 / 162 = 0
    16'b10001101_10100011 : OUT <= 0;  //141 / 163 = 0
    16'b10001101_10100100 : OUT <= 0;  //141 / 164 = 0
    16'b10001101_10100101 : OUT <= 0;  //141 / 165 = 0
    16'b10001101_10100110 : OUT <= 0;  //141 / 166 = 0
    16'b10001101_10100111 : OUT <= 0;  //141 / 167 = 0
    16'b10001101_10101000 : OUT <= 0;  //141 / 168 = 0
    16'b10001101_10101001 : OUT <= 0;  //141 / 169 = 0
    16'b10001101_10101010 : OUT <= 0;  //141 / 170 = 0
    16'b10001101_10101011 : OUT <= 0;  //141 / 171 = 0
    16'b10001101_10101100 : OUT <= 0;  //141 / 172 = 0
    16'b10001101_10101101 : OUT <= 0;  //141 / 173 = 0
    16'b10001101_10101110 : OUT <= 0;  //141 / 174 = 0
    16'b10001101_10101111 : OUT <= 0;  //141 / 175 = 0
    16'b10001101_10110000 : OUT <= 0;  //141 / 176 = 0
    16'b10001101_10110001 : OUT <= 0;  //141 / 177 = 0
    16'b10001101_10110010 : OUT <= 0;  //141 / 178 = 0
    16'b10001101_10110011 : OUT <= 0;  //141 / 179 = 0
    16'b10001101_10110100 : OUT <= 0;  //141 / 180 = 0
    16'b10001101_10110101 : OUT <= 0;  //141 / 181 = 0
    16'b10001101_10110110 : OUT <= 0;  //141 / 182 = 0
    16'b10001101_10110111 : OUT <= 0;  //141 / 183 = 0
    16'b10001101_10111000 : OUT <= 0;  //141 / 184 = 0
    16'b10001101_10111001 : OUT <= 0;  //141 / 185 = 0
    16'b10001101_10111010 : OUT <= 0;  //141 / 186 = 0
    16'b10001101_10111011 : OUT <= 0;  //141 / 187 = 0
    16'b10001101_10111100 : OUT <= 0;  //141 / 188 = 0
    16'b10001101_10111101 : OUT <= 0;  //141 / 189 = 0
    16'b10001101_10111110 : OUT <= 0;  //141 / 190 = 0
    16'b10001101_10111111 : OUT <= 0;  //141 / 191 = 0
    16'b10001101_11000000 : OUT <= 0;  //141 / 192 = 0
    16'b10001101_11000001 : OUT <= 0;  //141 / 193 = 0
    16'b10001101_11000010 : OUT <= 0;  //141 / 194 = 0
    16'b10001101_11000011 : OUT <= 0;  //141 / 195 = 0
    16'b10001101_11000100 : OUT <= 0;  //141 / 196 = 0
    16'b10001101_11000101 : OUT <= 0;  //141 / 197 = 0
    16'b10001101_11000110 : OUT <= 0;  //141 / 198 = 0
    16'b10001101_11000111 : OUT <= 0;  //141 / 199 = 0
    16'b10001101_11001000 : OUT <= 0;  //141 / 200 = 0
    16'b10001101_11001001 : OUT <= 0;  //141 / 201 = 0
    16'b10001101_11001010 : OUT <= 0;  //141 / 202 = 0
    16'b10001101_11001011 : OUT <= 0;  //141 / 203 = 0
    16'b10001101_11001100 : OUT <= 0;  //141 / 204 = 0
    16'b10001101_11001101 : OUT <= 0;  //141 / 205 = 0
    16'b10001101_11001110 : OUT <= 0;  //141 / 206 = 0
    16'b10001101_11001111 : OUT <= 0;  //141 / 207 = 0
    16'b10001101_11010000 : OUT <= 0;  //141 / 208 = 0
    16'b10001101_11010001 : OUT <= 0;  //141 / 209 = 0
    16'b10001101_11010010 : OUT <= 0;  //141 / 210 = 0
    16'b10001101_11010011 : OUT <= 0;  //141 / 211 = 0
    16'b10001101_11010100 : OUT <= 0;  //141 / 212 = 0
    16'b10001101_11010101 : OUT <= 0;  //141 / 213 = 0
    16'b10001101_11010110 : OUT <= 0;  //141 / 214 = 0
    16'b10001101_11010111 : OUT <= 0;  //141 / 215 = 0
    16'b10001101_11011000 : OUT <= 0;  //141 / 216 = 0
    16'b10001101_11011001 : OUT <= 0;  //141 / 217 = 0
    16'b10001101_11011010 : OUT <= 0;  //141 / 218 = 0
    16'b10001101_11011011 : OUT <= 0;  //141 / 219 = 0
    16'b10001101_11011100 : OUT <= 0;  //141 / 220 = 0
    16'b10001101_11011101 : OUT <= 0;  //141 / 221 = 0
    16'b10001101_11011110 : OUT <= 0;  //141 / 222 = 0
    16'b10001101_11011111 : OUT <= 0;  //141 / 223 = 0
    16'b10001101_11100000 : OUT <= 0;  //141 / 224 = 0
    16'b10001101_11100001 : OUT <= 0;  //141 / 225 = 0
    16'b10001101_11100010 : OUT <= 0;  //141 / 226 = 0
    16'b10001101_11100011 : OUT <= 0;  //141 / 227 = 0
    16'b10001101_11100100 : OUT <= 0;  //141 / 228 = 0
    16'b10001101_11100101 : OUT <= 0;  //141 / 229 = 0
    16'b10001101_11100110 : OUT <= 0;  //141 / 230 = 0
    16'b10001101_11100111 : OUT <= 0;  //141 / 231 = 0
    16'b10001101_11101000 : OUT <= 0;  //141 / 232 = 0
    16'b10001101_11101001 : OUT <= 0;  //141 / 233 = 0
    16'b10001101_11101010 : OUT <= 0;  //141 / 234 = 0
    16'b10001101_11101011 : OUT <= 0;  //141 / 235 = 0
    16'b10001101_11101100 : OUT <= 0;  //141 / 236 = 0
    16'b10001101_11101101 : OUT <= 0;  //141 / 237 = 0
    16'b10001101_11101110 : OUT <= 0;  //141 / 238 = 0
    16'b10001101_11101111 : OUT <= 0;  //141 / 239 = 0
    16'b10001101_11110000 : OUT <= 0;  //141 / 240 = 0
    16'b10001101_11110001 : OUT <= 0;  //141 / 241 = 0
    16'b10001101_11110010 : OUT <= 0;  //141 / 242 = 0
    16'b10001101_11110011 : OUT <= 0;  //141 / 243 = 0
    16'b10001101_11110100 : OUT <= 0;  //141 / 244 = 0
    16'b10001101_11110101 : OUT <= 0;  //141 / 245 = 0
    16'b10001101_11110110 : OUT <= 0;  //141 / 246 = 0
    16'b10001101_11110111 : OUT <= 0;  //141 / 247 = 0
    16'b10001101_11111000 : OUT <= 0;  //141 / 248 = 0
    16'b10001101_11111001 : OUT <= 0;  //141 / 249 = 0
    16'b10001101_11111010 : OUT <= 0;  //141 / 250 = 0
    16'b10001101_11111011 : OUT <= 0;  //141 / 251 = 0
    16'b10001101_11111100 : OUT <= 0;  //141 / 252 = 0
    16'b10001101_11111101 : OUT <= 0;  //141 / 253 = 0
    16'b10001101_11111110 : OUT <= 0;  //141 / 254 = 0
    16'b10001101_11111111 : OUT <= 0;  //141 / 255 = 0
    16'b10001110_00000000 : OUT <= 0;  //142 / 0 = 0
    16'b10001110_00000001 : OUT <= 142;  //142 / 1 = 142
    16'b10001110_00000010 : OUT <= 71;  //142 / 2 = 71
    16'b10001110_00000011 : OUT <= 47;  //142 / 3 = 47
    16'b10001110_00000100 : OUT <= 35;  //142 / 4 = 35
    16'b10001110_00000101 : OUT <= 28;  //142 / 5 = 28
    16'b10001110_00000110 : OUT <= 23;  //142 / 6 = 23
    16'b10001110_00000111 : OUT <= 20;  //142 / 7 = 20
    16'b10001110_00001000 : OUT <= 17;  //142 / 8 = 17
    16'b10001110_00001001 : OUT <= 15;  //142 / 9 = 15
    16'b10001110_00001010 : OUT <= 14;  //142 / 10 = 14
    16'b10001110_00001011 : OUT <= 12;  //142 / 11 = 12
    16'b10001110_00001100 : OUT <= 11;  //142 / 12 = 11
    16'b10001110_00001101 : OUT <= 10;  //142 / 13 = 10
    16'b10001110_00001110 : OUT <= 10;  //142 / 14 = 10
    16'b10001110_00001111 : OUT <= 9;  //142 / 15 = 9
    16'b10001110_00010000 : OUT <= 8;  //142 / 16 = 8
    16'b10001110_00010001 : OUT <= 8;  //142 / 17 = 8
    16'b10001110_00010010 : OUT <= 7;  //142 / 18 = 7
    16'b10001110_00010011 : OUT <= 7;  //142 / 19 = 7
    16'b10001110_00010100 : OUT <= 7;  //142 / 20 = 7
    16'b10001110_00010101 : OUT <= 6;  //142 / 21 = 6
    16'b10001110_00010110 : OUT <= 6;  //142 / 22 = 6
    16'b10001110_00010111 : OUT <= 6;  //142 / 23 = 6
    16'b10001110_00011000 : OUT <= 5;  //142 / 24 = 5
    16'b10001110_00011001 : OUT <= 5;  //142 / 25 = 5
    16'b10001110_00011010 : OUT <= 5;  //142 / 26 = 5
    16'b10001110_00011011 : OUT <= 5;  //142 / 27 = 5
    16'b10001110_00011100 : OUT <= 5;  //142 / 28 = 5
    16'b10001110_00011101 : OUT <= 4;  //142 / 29 = 4
    16'b10001110_00011110 : OUT <= 4;  //142 / 30 = 4
    16'b10001110_00011111 : OUT <= 4;  //142 / 31 = 4
    16'b10001110_00100000 : OUT <= 4;  //142 / 32 = 4
    16'b10001110_00100001 : OUT <= 4;  //142 / 33 = 4
    16'b10001110_00100010 : OUT <= 4;  //142 / 34 = 4
    16'b10001110_00100011 : OUT <= 4;  //142 / 35 = 4
    16'b10001110_00100100 : OUT <= 3;  //142 / 36 = 3
    16'b10001110_00100101 : OUT <= 3;  //142 / 37 = 3
    16'b10001110_00100110 : OUT <= 3;  //142 / 38 = 3
    16'b10001110_00100111 : OUT <= 3;  //142 / 39 = 3
    16'b10001110_00101000 : OUT <= 3;  //142 / 40 = 3
    16'b10001110_00101001 : OUT <= 3;  //142 / 41 = 3
    16'b10001110_00101010 : OUT <= 3;  //142 / 42 = 3
    16'b10001110_00101011 : OUT <= 3;  //142 / 43 = 3
    16'b10001110_00101100 : OUT <= 3;  //142 / 44 = 3
    16'b10001110_00101101 : OUT <= 3;  //142 / 45 = 3
    16'b10001110_00101110 : OUT <= 3;  //142 / 46 = 3
    16'b10001110_00101111 : OUT <= 3;  //142 / 47 = 3
    16'b10001110_00110000 : OUT <= 2;  //142 / 48 = 2
    16'b10001110_00110001 : OUT <= 2;  //142 / 49 = 2
    16'b10001110_00110010 : OUT <= 2;  //142 / 50 = 2
    16'b10001110_00110011 : OUT <= 2;  //142 / 51 = 2
    16'b10001110_00110100 : OUT <= 2;  //142 / 52 = 2
    16'b10001110_00110101 : OUT <= 2;  //142 / 53 = 2
    16'b10001110_00110110 : OUT <= 2;  //142 / 54 = 2
    16'b10001110_00110111 : OUT <= 2;  //142 / 55 = 2
    16'b10001110_00111000 : OUT <= 2;  //142 / 56 = 2
    16'b10001110_00111001 : OUT <= 2;  //142 / 57 = 2
    16'b10001110_00111010 : OUT <= 2;  //142 / 58 = 2
    16'b10001110_00111011 : OUT <= 2;  //142 / 59 = 2
    16'b10001110_00111100 : OUT <= 2;  //142 / 60 = 2
    16'b10001110_00111101 : OUT <= 2;  //142 / 61 = 2
    16'b10001110_00111110 : OUT <= 2;  //142 / 62 = 2
    16'b10001110_00111111 : OUT <= 2;  //142 / 63 = 2
    16'b10001110_01000000 : OUT <= 2;  //142 / 64 = 2
    16'b10001110_01000001 : OUT <= 2;  //142 / 65 = 2
    16'b10001110_01000010 : OUT <= 2;  //142 / 66 = 2
    16'b10001110_01000011 : OUT <= 2;  //142 / 67 = 2
    16'b10001110_01000100 : OUT <= 2;  //142 / 68 = 2
    16'b10001110_01000101 : OUT <= 2;  //142 / 69 = 2
    16'b10001110_01000110 : OUT <= 2;  //142 / 70 = 2
    16'b10001110_01000111 : OUT <= 2;  //142 / 71 = 2
    16'b10001110_01001000 : OUT <= 1;  //142 / 72 = 1
    16'b10001110_01001001 : OUT <= 1;  //142 / 73 = 1
    16'b10001110_01001010 : OUT <= 1;  //142 / 74 = 1
    16'b10001110_01001011 : OUT <= 1;  //142 / 75 = 1
    16'b10001110_01001100 : OUT <= 1;  //142 / 76 = 1
    16'b10001110_01001101 : OUT <= 1;  //142 / 77 = 1
    16'b10001110_01001110 : OUT <= 1;  //142 / 78 = 1
    16'b10001110_01001111 : OUT <= 1;  //142 / 79 = 1
    16'b10001110_01010000 : OUT <= 1;  //142 / 80 = 1
    16'b10001110_01010001 : OUT <= 1;  //142 / 81 = 1
    16'b10001110_01010010 : OUT <= 1;  //142 / 82 = 1
    16'b10001110_01010011 : OUT <= 1;  //142 / 83 = 1
    16'b10001110_01010100 : OUT <= 1;  //142 / 84 = 1
    16'b10001110_01010101 : OUT <= 1;  //142 / 85 = 1
    16'b10001110_01010110 : OUT <= 1;  //142 / 86 = 1
    16'b10001110_01010111 : OUT <= 1;  //142 / 87 = 1
    16'b10001110_01011000 : OUT <= 1;  //142 / 88 = 1
    16'b10001110_01011001 : OUT <= 1;  //142 / 89 = 1
    16'b10001110_01011010 : OUT <= 1;  //142 / 90 = 1
    16'b10001110_01011011 : OUT <= 1;  //142 / 91 = 1
    16'b10001110_01011100 : OUT <= 1;  //142 / 92 = 1
    16'b10001110_01011101 : OUT <= 1;  //142 / 93 = 1
    16'b10001110_01011110 : OUT <= 1;  //142 / 94 = 1
    16'b10001110_01011111 : OUT <= 1;  //142 / 95 = 1
    16'b10001110_01100000 : OUT <= 1;  //142 / 96 = 1
    16'b10001110_01100001 : OUT <= 1;  //142 / 97 = 1
    16'b10001110_01100010 : OUT <= 1;  //142 / 98 = 1
    16'b10001110_01100011 : OUT <= 1;  //142 / 99 = 1
    16'b10001110_01100100 : OUT <= 1;  //142 / 100 = 1
    16'b10001110_01100101 : OUT <= 1;  //142 / 101 = 1
    16'b10001110_01100110 : OUT <= 1;  //142 / 102 = 1
    16'b10001110_01100111 : OUT <= 1;  //142 / 103 = 1
    16'b10001110_01101000 : OUT <= 1;  //142 / 104 = 1
    16'b10001110_01101001 : OUT <= 1;  //142 / 105 = 1
    16'b10001110_01101010 : OUT <= 1;  //142 / 106 = 1
    16'b10001110_01101011 : OUT <= 1;  //142 / 107 = 1
    16'b10001110_01101100 : OUT <= 1;  //142 / 108 = 1
    16'b10001110_01101101 : OUT <= 1;  //142 / 109 = 1
    16'b10001110_01101110 : OUT <= 1;  //142 / 110 = 1
    16'b10001110_01101111 : OUT <= 1;  //142 / 111 = 1
    16'b10001110_01110000 : OUT <= 1;  //142 / 112 = 1
    16'b10001110_01110001 : OUT <= 1;  //142 / 113 = 1
    16'b10001110_01110010 : OUT <= 1;  //142 / 114 = 1
    16'b10001110_01110011 : OUT <= 1;  //142 / 115 = 1
    16'b10001110_01110100 : OUT <= 1;  //142 / 116 = 1
    16'b10001110_01110101 : OUT <= 1;  //142 / 117 = 1
    16'b10001110_01110110 : OUT <= 1;  //142 / 118 = 1
    16'b10001110_01110111 : OUT <= 1;  //142 / 119 = 1
    16'b10001110_01111000 : OUT <= 1;  //142 / 120 = 1
    16'b10001110_01111001 : OUT <= 1;  //142 / 121 = 1
    16'b10001110_01111010 : OUT <= 1;  //142 / 122 = 1
    16'b10001110_01111011 : OUT <= 1;  //142 / 123 = 1
    16'b10001110_01111100 : OUT <= 1;  //142 / 124 = 1
    16'b10001110_01111101 : OUT <= 1;  //142 / 125 = 1
    16'b10001110_01111110 : OUT <= 1;  //142 / 126 = 1
    16'b10001110_01111111 : OUT <= 1;  //142 / 127 = 1
    16'b10001110_10000000 : OUT <= 1;  //142 / 128 = 1
    16'b10001110_10000001 : OUT <= 1;  //142 / 129 = 1
    16'b10001110_10000010 : OUT <= 1;  //142 / 130 = 1
    16'b10001110_10000011 : OUT <= 1;  //142 / 131 = 1
    16'b10001110_10000100 : OUT <= 1;  //142 / 132 = 1
    16'b10001110_10000101 : OUT <= 1;  //142 / 133 = 1
    16'b10001110_10000110 : OUT <= 1;  //142 / 134 = 1
    16'b10001110_10000111 : OUT <= 1;  //142 / 135 = 1
    16'b10001110_10001000 : OUT <= 1;  //142 / 136 = 1
    16'b10001110_10001001 : OUT <= 1;  //142 / 137 = 1
    16'b10001110_10001010 : OUT <= 1;  //142 / 138 = 1
    16'b10001110_10001011 : OUT <= 1;  //142 / 139 = 1
    16'b10001110_10001100 : OUT <= 1;  //142 / 140 = 1
    16'b10001110_10001101 : OUT <= 1;  //142 / 141 = 1
    16'b10001110_10001110 : OUT <= 1;  //142 / 142 = 1
    16'b10001110_10001111 : OUT <= 0;  //142 / 143 = 0
    16'b10001110_10010000 : OUT <= 0;  //142 / 144 = 0
    16'b10001110_10010001 : OUT <= 0;  //142 / 145 = 0
    16'b10001110_10010010 : OUT <= 0;  //142 / 146 = 0
    16'b10001110_10010011 : OUT <= 0;  //142 / 147 = 0
    16'b10001110_10010100 : OUT <= 0;  //142 / 148 = 0
    16'b10001110_10010101 : OUT <= 0;  //142 / 149 = 0
    16'b10001110_10010110 : OUT <= 0;  //142 / 150 = 0
    16'b10001110_10010111 : OUT <= 0;  //142 / 151 = 0
    16'b10001110_10011000 : OUT <= 0;  //142 / 152 = 0
    16'b10001110_10011001 : OUT <= 0;  //142 / 153 = 0
    16'b10001110_10011010 : OUT <= 0;  //142 / 154 = 0
    16'b10001110_10011011 : OUT <= 0;  //142 / 155 = 0
    16'b10001110_10011100 : OUT <= 0;  //142 / 156 = 0
    16'b10001110_10011101 : OUT <= 0;  //142 / 157 = 0
    16'b10001110_10011110 : OUT <= 0;  //142 / 158 = 0
    16'b10001110_10011111 : OUT <= 0;  //142 / 159 = 0
    16'b10001110_10100000 : OUT <= 0;  //142 / 160 = 0
    16'b10001110_10100001 : OUT <= 0;  //142 / 161 = 0
    16'b10001110_10100010 : OUT <= 0;  //142 / 162 = 0
    16'b10001110_10100011 : OUT <= 0;  //142 / 163 = 0
    16'b10001110_10100100 : OUT <= 0;  //142 / 164 = 0
    16'b10001110_10100101 : OUT <= 0;  //142 / 165 = 0
    16'b10001110_10100110 : OUT <= 0;  //142 / 166 = 0
    16'b10001110_10100111 : OUT <= 0;  //142 / 167 = 0
    16'b10001110_10101000 : OUT <= 0;  //142 / 168 = 0
    16'b10001110_10101001 : OUT <= 0;  //142 / 169 = 0
    16'b10001110_10101010 : OUT <= 0;  //142 / 170 = 0
    16'b10001110_10101011 : OUT <= 0;  //142 / 171 = 0
    16'b10001110_10101100 : OUT <= 0;  //142 / 172 = 0
    16'b10001110_10101101 : OUT <= 0;  //142 / 173 = 0
    16'b10001110_10101110 : OUT <= 0;  //142 / 174 = 0
    16'b10001110_10101111 : OUT <= 0;  //142 / 175 = 0
    16'b10001110_10110000 : OUT <= 0;  //142 / 176 = 0
    16'b10001110_10110001 : OUT <= 0;  //142 / 177 = 0
    16'b10001110_10110010 : OUT <= 0;  //142 / 178 = 0
    16'b10001110_10110011 : OUT <= 0;  //142 / 179 = 0
    16'b10001110_10110100 : OUT <= 0;  //142 / 180 = 0
    16'b10001110_10110101 : OUT <= 0;  //142 / 181 = 0
    16'b10001110_10110110 : OUT <= 0;  //142 / 182 = 0
    16'b10001110_10110111 : OUT <= 0;  //142 / 183 = 0
    16'b10001110_10111000 : OUT <= 0;  //142 / 184 = 0
    16'b10001110_10111001 : OUT <= 0;  //142 / 185 = 0
    16'b10001110_10111010 : OUT <= 0;  //142 / 186 = 0
    16'b10001110_10111011 : OUT <= 0;  //142 / 187 = 0
    16'b10001110_10111100 : OUT <= 0;  //142 / 188 = 0
    16'b10001110_10111101 : OUT <= 0;  //142 / 189 = 0
    16'b10001110_10111110 : OUT <= 0;  //142 / 190 = 0
    16'b10001110_10111111 : OUT <= 0;  //142 / 191 = 0
    16'b10001110_11000000 : OUT <= 0;  //142 / 192 = 0
    16'b10001110_11000001 : OUT <= 0;  //142 / 193 = 0
    16'b10001110_11000010 : OUT <= 0;  //142 / 194 = 0
    16'b10001110_11000011 : OUT <= 0;  //142 / 195 = 0
    16'b10001110_11000100 : OUT <= 0;  //142 / 196 = 0
    16'b10001110_11000101 : OUT <= 0;  //142 / 197 = 0
    16'b10001110_11000110 : OUT <= 0;  //142 / 198 = 0
    16'b10001110_11000111 : OUT <= 0;  //142 / 199 = 0
    16'b10001110_11001000 : OUT <= 0;  //142 / 200 = 0
    16'b10001110_11001001 : OUT <= 0;  //142 / 201 = 0
    16'b10001110_11001010 : OUT <= 0;  //142 / 202 = 0
    16'b10001110_11001011 : OUT <= 0;  //142 / 203 = 0
    16'b10001110_11001100 : OUT <= 0;  //142 / 204 = 0
    16'b10001110_11001101 : OUT <= 0;  //142 / 205 = 0
    16'b10001110_11001110 : OUT <= 0;  //142 / 206 = 0
    16'b10001110_11001111 : OUT <= 0;  //142 / 207 = 0
    16'b10001110_11010000 : OUT <= 0;  //142 / 208 = 0
    16'b10001110_11010001 : OUT <= 0;  //142 / 209 = 0
    16'b10001110_11010010 : OUT <= 0;  //142 / 210 = 0
    16'b10001110_11010011 : OUT <= 0;  //142 / 211 = 0
    16'b10001110_11010100 : OUT <= 0;  //142 / 212 = 0
    16'b10001110_11010101 : OUT <= 0;  //142 / 213 = 0
    16'b10001110_11010110 : OUT <= 0;  //142 / 214 = 0
    16'b10001110_11010111 : OUT <= 0;  //142 / 215 = 0
    16'b10001110_11011000 : OUT <= 0;  //142 / 216 = 0
    16'b10001110_11011001 : OUT <= 0;  //142 / 217 = 0
    16'b10001110_11011010 : OUT <= 0;  //142 / 218 = 0
    16'b10001110_11011011 : OUT <= 0;  //142 / 219 = 0
    16'b10001110_11011100 : OUT <= 0;  //142 / 220 = 0
    16'b10001110_11011101 : OUT <= 0;  //142 / 221 = 0
    16'b10001110_11011110 : OUT <= 0;  //142 / 222 = 0
    16'b10001110_11011111 : OUT <= 0;  //142 / 223 = 0
    16'b10001110_11100000 : OUT <= 0;  //142 / 224 = 0
    16'b10001110_11100001 : OUT <= 0;  //142 / 225 = 0
    16'b10001110_11100010 : OUT <= 0;  //142 / 226 = 0
    16'b10001110_11100011 : OUT <= 0;  //142 / 227 = 0
    16'b10001110_11100100 : OUT <= 0;  //142 / 228 = 0
    16'b10001110_11100101 : OUT <= 0;  //142 / 229 = 0
    16'b10001110_11100110 : OUT <= 0;  //142 / 230 = 0
    16'b10001110_11100111 : OUT <= 0;  //142 / 231 = 0
    16'b10001110_11101000 : OUT <= 0;  //142 / 232 = 0
    16'b10001110_11101001 : OUT <= 0;  //142 / 233 = 0
    16'b10001110_11101010 : OUT <= 0;  //142 / 234 = 0
    16'b10001110_11101011 : OUT <= 0;  //142 / 235 = 0
    16'b10001110_11101100 : OUT <= 0;  //142 / 236 = 0
    16'b10001110_11101101 : OUT <= 0;  //142 / 237 = 0
    16'b10001110_11101110 : OUT <= 0;  //142 / 238 = 0
    16'b10001110_11101111 : OUT <= 0;  //142 / 239 = 0
    16'b10001110_11110000 : OUT <= 0;  //142 / 240 = 0
    16'b10001110_11110001 : OUT <= 0;  //142 / 241 = 0
    16'b10001110_11110010 : OUT <= 0;  //142 / 242 = 0
    16'b10001110_11110011 : OUT <= 0;  //142 / 243 = 0
    16'b10001110_11110100 : OUT <= 0;  //142 / 244 = 0
    16'b10001110_11110101 : OUT <= 0;  //142 / 245 = 0
    16'b10001110_11110110 : OUT <= 0;  //142 / 246 = 0
    16'b10001110_11110111 : OUT <= 0;  //142 / 247 = 0
    16'b10001110_11111000 : OUT <= 0;  //142 / 248 = 0
    16'b10001110_11111001 : OUT <= 0;  //142 / 249 = 0
    16'b10001110_11111010 : OUT <= 0;  //142 / 250 = 0
    16'b10001110_11111011 : OUT <= 0;  //142 / 251 = 0
    16'b10001110_11111100 : OUT <= 0;  //142 / 252 = 0
    16'b10001110_11111101 : OUT <= 0;  //142 / 253 = 0
    16'b10001110_11111110 : OUT <= 0;  //142 / 254 = 0
    16'b10001110_11111111 : OUT <= 0;  //142 / 255 = 0
    16'b10001111_00000000 : OUT <= 0;  //143 / 0 = 0
    16'b10001111_00000001 : OUT <= 143;  //143 / 1 = 143
    16'b10001111_00000010 : OUT <= 71;  //143 / 2 = 71
    16'b10001111_00000011 : OUT <= 47;  //143 / 3 = 47
    16'b10001111_00000100 : OUT <= 35;  //143 / 4 = 35
    16'b10001111_00000101 : OUT <= 28;  //143 / 5 = 28
    16'b10001111_00000110 : OUT <= 23;  //143 / 6 = 23
    16'b10001111_00000111 : OUT <= 20;  //143 / 7 = 20
    16'b10001111_00001000 : OUT <= 17;  //143 / 8 = 17
    16'b10001111_00001001 : OUT <= 15;  //143 / 9 = 15
    16'b10001111_00001010 : OUT <= 14;  //143 / 10 = 14
    16'b10001111_00001011 : OUT <= 13;  //143 / 11 = 13
    16'b10001111_00001100 : OUT <= 11;  //143 / 12 = 11
    16'b10001111_00001101 : OUT <= 11;  //143 / 13 = 11
    16'b10001111_00001110 : OUT <= 10;  //143 / 14 = 10
    16'b10001111_00001111 : OUT <= 9;  //143 / 15 = 9
    16'b10001111_00010000 : OUT <= 8;  //143 / 16 = 8
    16'b10001111_00010001 : OUT <= 8;  //143 / 17 = 8
    16'b10001111_00010010 : OUT <= 7;  //143 / 18 = 7
    16'b10001111_00010011 : OUT <= 7;  //143 / 19 = 7
    16'b10001111_00010100 : OUT <= 7;  //143 / 20 = 7
    16'b10001111_00010101 : OUT <= 6;  //143 / 21 = 6
    16'b10001111_00010110 : OUT <= 6;  //143 / 22 = 6
    16'b10001111_00010111 : OUT <= 6;  //143 / 23 = 6
    16'b10001111_00011000 : OUT <= 5;  //143 / 24 = 5
    16'b10001111_00011001 : OUT <= 5;  //143 / 25 = 5
    16'b10001111_00011010 : OUT <= 5;  //143 / 26 = 5
    16'b10001111_00011011 : OUT <= 5;  //143 / 27 = 5
    16'b10001111_00011100 : OUT <= 5;  //143 / 28 = 5
    16'b10001111_00011101 : OUT <= 4;  //143 / 29 = 4
    16'b10001111_00011110 : OUT <= 4;  //143 / 30 = 4
    16'b10001111_00011111 : OUT <= 4;  //143 / 31 = 4
    16'b10001111_00100000 : OUT <= 4;  //143 / 32 = 4
    16'b10001111_00100001 : OUT <= 4;  //143 / 33 = 4
    16'b10001111_00100010 : OUT <= 4;  //143 / 34 = 4
    16'b10001111_00100011 : OUT <= 4;  //143 / 35 = 4
    16'b10001111_00100100 : OUT <= 3;  //143 / 36 = 3
    16'b10001111_00100101 : OUT <= 3;  //143 / 37 = 3
    16'b10001111_00100110 : OUT <= 3;  //143 / 38 = 3
    16'b10001111_00100111 : OUT <= 3;  //143 / 39 = 3
    16'b10001111_00101000 : OUT <= 3;  //143 / 40 = 3
    16'b10001111_00101001 : OUT <= 3;  //143 / 41 = 3
    16'b10001111_00101010 : OUT <= 3;  //143 / 42 = 3
    16'b10001111_00101011 : OUT <= 3;  //143 / 43 = 3
    16'b10001111_00101100 : OUT <= 3;  //143 / 44 = 3
    16'b10001111_00101101 : OUT <= 3;  //143 / 45 = 3
    16'b10001111_00101110 : OUT <= 3;  //143 / 46 = 3
    16'b10001111_00101111 : OUT <= 3;  //143 / 47 = 3
    16'b10001111_00110000 : OUT <= 2;  //143 / 48 = 2
    16'b10001111_00110001 : OUT <= 2;  //143 / 49 = 2
    16'b10001111_00110010 : OUT <= 2;  //143 / 50 = 2
    16'b10001111_00110011 : OUT <= 2;  //143 / 51 = 2
    16'b10001111_00110100 : OUT <= 2;  //143 / 52 = 2
    16'b10001111_00110101 : OUT <= 2;  //143 / 53 = 2
    16'b10001111_00110110 : OUT <= 2;  //143 / 54 = 2
    16'b10001111_00110111 : OUT <= 2;  //143 / 55 = 2
    16'b10001111_00111000 : OUT <= 2;  //143 / 56 = 2
    16'b10001111_00111001 : OUT <= 2;  //143 / 57 = 2
    16'b10001111_00111010 : OUT <= 2;  //143 / 58 = 2
    16'b10001111_00111011 : OUT <= 2;  //143 / 59 = 2
    16'b10001111_00111100 : OUT <= 2;  //143 / 60 = 2
    16'b10001111_00111101 : OUT <= 2;  //143 / 61 = 2
    16'b10001111_00111110 : OUT <= 2;  //143 / 62 = 2
    16'b10001111_00111111 : OUT <= 2;  //143 / 63 = 2
    16'b10001111_01000000 : OUT <= 2;  //143 / 64 = 2
    16'b10001111_01000001 : OUT <= 2;  //143 / 65 = 2
    16'b10001111_01000010 : OUT <= 2;  //143 / 66 = 2
    16'b10001111_01000011 : OUT <= 2;  //143 / 67 = 2
    16'b10001111_01000100 : OUT <= 2;  //143 / 68 = 2
    16'b10001111_01000101 : OUT <= 2;  //143 / 69 = 2
    16'b10001111_01000110 : OUT <= 2;  //143 / 70 = 2
    16'b10001111_01000111 : OUT <= 2;  //143 / 71 = 2
    16'b10001111_01001000 : OUT <= 1;  //143 / 72 = 1
    16'b10001111_01001001 : OUT <= 1;  //143 / 73 = 1
    16'b10001111_01001010 : OUT <= 1;  //143 / 74 = 1
    16'b10001111_01001011 : OUT <= 1;  //143 / 75 = 1
    16'b10001111_01001100 : OUT <= 1;  //143 / 76 = 1
    16'b10001111_01001101 : OUT <= 1;  //143 / 77 = 1
    16'b10001111_01001110 : OUT <= 1;  //143 / 78 = 1
    16'b10001111_01001111 : OUT <= 1;  //143 / 79 = 1
    16'b10001111_01010000 : OUT <= 1;  //143 / 80 = 1
    16'b10001111_01010001 : OUT <= 1;  //143 / 81 = 1
    16'b10001111_01010010 : OUT <= 1;  //143 / 82 = 1
    16'b10001111_01010011 : OUT <= 1;  //143 / 83 = 1
    16'b10001111_01010100 : OUT <= 1;  //143 / 84 = 1
    16'b10001111_01010101 : OUT <= 1;  //143 / 85 = 1
    16'b10001111_01010110 : OUT <= 1;  //143 / 86 = 1
    16'b10001111_01010111 : OUT <= 1;  //143 / 87 = 1
    16'b10001111_01011000 : OUT <= 1;  //143 / 88 = 1
    16'b10001111_01011001 : OUT <= 1;  //143 / 89 = 1
    16'b10001111_01011010 : OUT <= 1;  //143 / 90 = 1
    16'b10001111_01011011 : OUT <= 1;  //143 / 91 = 1
    16'b10001111_01011100 : OUT <= 1;  //143 / 92 = 1
    16'b10001111_01011101 : OUT <= 1;  //143 / 93 = 1
    16'b10001111_01011110 : OUT <= 1;  //143 / 94 = 1
    16'b10001111_01011111 : OUT <= 1;  //143 / 95 = 1
    16'b10001111_01100000 : OUT <= 1;  //143 / 96 = 1
    16'b10001111_01100001 : OUT <= 1;  //143 / 97 = 1
    16'b10001111_01100010 : OUT <= 1;  //143 / 98 = 1
    16'b10001111_01100011 : OUT <= 1;  //143 / 99 = 1
    16'b10001111_01100100 : OUT <= 1;  //143 / 100 = 1
    16'b10001111_01100101 : OUT <= 1;  //143 / 101 = 1
    16'b10001111_01100110 : OUT <= 1;  //143 / 102 = 1
    16'b10001111_01100111 : OUT <= 1;  //143 / 103 = 1
    16'b10001111_01101000 : OUT <= 1;  //143 / 104 = 1
    16'b10001111_01101001 : OUT <= 1;  //143 / 105 = 1
    16'b10001111_01101010 : OUT <= 1;  //143 / 106 = 1
    16'b10001111_01101011 : OUT <= 1;  //143 / 107 = 1
    16'b10001111_01101100 : OUT <= 1;  //143 / 108 = 1
    16'b10001111_01101101 : OUT <= 1;  //143 / 109 = 1
    16'b10001111_01101110 : OUT <= 1;  //143 / 110 = 1
    16'b10001111_01101111 : OUT <= 1;  //143 / 111 = 1
    16'b10001111_01110000 : OUT <= 1;  //143 / 112 = 1
    16'b10001111_01110001 : OUT <= 1;  //143 / 113 = 1
    16'b10001111_01110010 : OUT <= 1;  //143 / 114 = 1
    16'b10001111_01110011 : OUT <= 1;  //143 / 115 = 1
    16'b10001111_01110100 : OUT <= 1;  //143 / 116 = 1
    16'b10001111_01110101 : OUT <= 1;  //143 / 117 = 1
    16'b10001111_01110110 : OUT <= 1;  //143 / 118 = 1
    16'b10001111_01110111 : OUT <= 1;  //143 / 119 = 1
    16'b10001111_01111000 : OUT <= 1;  //143 / 120 = 1
    16'b10001111_01111001 : OUT <= 1;  //143 / 121 = 1
    16'b10001111_01111010 : OUT <= 1;  //143 / 122 = 1
    16'b10001111_01111011 : OUT <= 1;  //143 / 123 = 1
    16'b10001111_01111100 : OUT <= 1;  //143 / 124 = 1
    16'b10001111_01111101 : OUT <= 1;  //143 / 125 = 1
    16'b10001111_01111110 : OUT <= 1;  //143 / 126 = 1
    16'b10001111_01111111 : OUT <= 1;  //143 / 127 = 1
    16'b10001111_10000000 : OUT <= 1;  //143 / 128 = 1
    16'b10001111_10000001 : OUT <= 1;  //143 / 129 = 1
    16'b10001111_10000010 : OUT <= 1;  //143 / 130 = 1
    16'b10001111_10000011 : OUT <= 1;  //143 / 131 = 1
    16'b10001111_10000100 : OUT <= 1;  //143 / 132 = 1
    16'b10001111_10000101 : OUT <= 1;  //143 / 133 = 1
    16'b10001111_10000110 : OUT <= 1;  //143 / 134 = 1
    16'b10001111_10000111 : OUT <= 1;  //143 / 135 = 1
    16'b10001111_10001000 : OUT <= 1;  //143 / 136 = 1
    16'b10001111_10001001 : OUT <= 1;  //143 / 137 = 1
    16'b10001111_10001010 : OUT <= 1;  //143 / 138 = 1
    16'b10001111_10001011 : OUT <= 1;  //143 / 139 = 1
    16'b10001111_10001100 : OUT <= 1;  //143 / 140 = 1
    16'b10001111_10001101 : OUT <= 1;  //143 / 141 = 1
    16'b10001111_10001110 : OUT <= 1;  //143 / 142 = 1
    16'b10001111_10001111 : OUT <= 1;  //143 / 143 = 1
    16'b10001111_10010000 : OUT <= 0;  //143 / 144 = 0
    16'b10001111_10010001 : OUT <= 0;  //143 / 145 = 0
    16'b10001111_10010010 : OUT <= 0;  //143 / 146 = 0
    16'b10001111_10010011 : OUT <= 0;  //143 / 147 = 0
    16'b10001111_10010100 : OUT <= 0;  //143 / 148 = 0
    16'b10001111_10010101 : OUT <= 0;  //143 / 149 = 0
    16'b10001111_10010110 : OUT <= 0;  //143 / 150 = 0
    16'b10001111_10010111 : OUT <= 0;  //143 / 151 = 0
    16'b10001111_10011000 : OUT <= 0;  //143 / 152 = 0
    16'b10001111_10011001 : OUT <= 0;  //143 / 153 = 0
    16'b10001111_10011010 : OUT <= 0;  //143 / 154 = 0
    16'b10001111_10011011 : OUT <= 0;  //143 / 155 = 0
    16'b10001111_10011100 : OUT <= 0;  //143 / 156 = 0
    16'b10001111_10011101 : OUT <= 0;  //143 / 157 = 0
    16'b10001111_10011110 : OUT <= 0;  //143 / 158 = 0
    16'b10001111_10011111 : OUT <= 0;  //143 / 159 = 0
    16'b10001111_10100000 : OUT <= 0;  //143 / 160 = 0
    16'b10001111_10100001 : OUT <= 0;  //143 / 161 = 0
    16'b10001111_10100010 : OUT <= 0;  //143 / 162 = 0
    16'b10001111_10100011 : OUT <= 0;  //143 / 163 = 0
    16'b10001111_10100100 : OUT <= 0;  //143 / 164 = 0
    16'b10001111_10100101 : OUT <= 0;  //143 / 165 = 0
    16'b10001111_10100110 : OUT <= 0;  //143 / 166 = 0
    16'b10001111_10100111 : OUT <= 0;  //143 / 167 = 0
    16'b10001111_10101000 : OUT <= 0;  //143 / 168 = 0
    16'b10001111_10101001 : OUT <= 0;  //143 / 169 = 0
    16'b10001111_10101010 : OUT <= 0;  //143 / 170 = 0
    16'b10001111_10101011 : OUT <= 0;  //143 / 171 = 0
    16'b10001111_10101100 : OUT <= 0;  //143 / 172 = 0
    16'b10001111_10101101 : OUT <= 0;  //143 / 173 = 0
    16'b10001111_10101110 : OUT <= 0;  //143 / 174 = 0
    16'b10001111_10101111 : OUT <= 0;  //143 / 175 = 0
    16'b10001111_10110000 : OUT <= 0;  //143 / 176 = 0
    16'b10001111_10110001 : OUT <= 0;  //143 / 177 = 0
    16'b10001111_10110010 : OUT <= 0;  //143 / 178 = 0
    16'b10001111_10110011 : OUT <= 0;  //143 / 179 = 0
    16'b10001111_10110100 : OUT <= 0;  //143 / 180 = 0
    16'b10001111_10110101 : OUT <= 0;  //143 / 181 = 0
    16'b10001111_10110110 : OUT <= 0;  //143 / 182 = 0
    16'b10001111_10110111 : OUT <= 0;  //143 / 183 = 0
    16'b10001111_10111000 : OUT <= 0;  //143 / 184 = 0
    16'b10001111_10111001 : OUT <= 0;  //143 / 185 = 0
    16'b10001111_10111010 : OUT <= 0;  //143 / 186 = 0
    16'b10001111_10111011 : OUT <= 0;  //143 / 187 = 0
    16'b10001111_10111100 : OUT <= 0;  //143 / 188 = 0
    16'b10001111_10111101 : OUT <= 0;  //143 / 189 = 0
    16'b10001111_10111110 : OUT <= 0;  //143 / 190 = 0
    16'b10001111_10111111 : OUT <= 0;  //143 / 191 = 0
    16'b10001111_11000000 : OUT <= 0;  //143 / 192 = 0
    16'b10001111_11000001 : OUT <= 0;  //143 / 193 = 0
    16'b10001111_11000010 : OUT <= 0;  //143 / 194 = 0
    16'b10001111_11000011 : OUT <= 0;  //143 / 195 = 0
    16'b10001111_11000100 : OUT <= 0;  //143 / 196 = 0
    16'b10001111_11000101 : OUT <= 0;  //143 / 197 = 0
    16'b10001111_11000110 : OUT <= 0;  //143 / 198 = 0
    16'b10001111_11000111 : OUT <= 0;  //143 / 199 = 0
    16'b10001111_11001000 : OUT <= 0;  //143 / 200 = 0
    16'b10001111_11001001 : OUT <= 0;  //143 / 201 = 0
    16'b10001111_11001010 : OUT <= 0;  //143 / 202 = 0
    16'b10001111_11001011 : OUT <= 0;  //143 / 203 = 0
    16'b10001111_11001100 : OUT <= 0;  //143 / 204 = 0
    16'b10001111_11001101 : OUT <= 0;  //143 / 205 = 0
    16'b10001111_11001110 : OUT <= 0;  //143 / 206 = 0
    16'b10001111_11001111 : OUT <= 0;  //143 / 207 = 0
    16'b10001111_11010000 : OUT <= 0;  //143 / 208 = 0
    16'b10001111_11010001 : OUT <= 0;  //143 / 209 = 0
    16'b10001111_11010010 : OUT <= 0;  //143 / 210 = 0
    16'b10001111_11010011 : OUT <= 0;  //143 / 211 = 0
    16'b10001111_11010100 : OUT <= 0;  //143 / 212 = 0
    16'b10001111_11010101 : OUT <= 0;  //143 / 213 = 0
    16'b10001111_11010110 : OUT <= 0;  //143 / 214 = 0
    16'b10001111_11010111 : OUT <= 0;  //143 / 215 = 0
    16'b10001111_11011000 : OUT <= 0;  //143 / 216 = 0
    16'b10001111_11011001 : OUT <= 0;  //143 / 217 = 0
    16'b10001111_11011010 : OUT <= 0;  //143 / 218 = 0
    16'b10001111_11011011 : OUT <= 0;  //143 / 219 = 0
    16'b10001111_11011100 : OUT <= 0;  //143 / 220 = 0
    16'b10001111_11011101 : OUT <= 0;  //143 / 221 = 0
    16'b10001111_11011110 : OUT <= 0;  //143 / 222 = 0
    16'b10001111_11011111 : OUT <= 0;  //143 / 223 = 0
    16'b10001111_11100000 : OUT <= 0;  //143 / 224 = 0
    16'b10001111_11100001 : OUT <= 0;  //143 / 225 = 0
    16'b10001111_11100010 : OUT <= 0;  //143 / 226 = 0
    16'b10001111_11100011 : OUT <= 0;  //143 / 227 = 0
    16'b10001111_11100100 : OUT <= 0;  //143 / 228 = 0
    16'b10001111_11100101 : OUT <= 0;  //143 / 229 = 0
    16'b10001111_11100110 : OUT <= 0;  //143 / 230 = 0
    16'b10001111_11100111 : OUT <= 0;  //143 / 231 = 0
    16'b10001111_11101000 : OUT <= 0;  //143 / 232 = 0
    16'b10001111_11101001 : OUT <= 0;  //143 / 233 = 0
    16'b10001111_11101010 : OUT <= 0;  //143 / 234 = 0
    16'b10001111_11101011 : OUT <= 0;  //143 / 235 = 0
    16'b10001111_11101100 : OUT <= 0;  //143 / 236 = 0
    16'b10001111_11101101 : OUT <= 0;  //143 / 237 = 0
    16'b10001111_11101110 : OUT <= 0;  //143 / 238 = 0
    16'b10001111_11101111 : OUT <= 0;  //143 / 239 = 0
    16'b10001111_11110000 : OUT <= 0;  //143 / 240 = 0
    16'b10001111_11110001 : OUT <= 0;  //143 / 241 = 0
    16'b10001111_11110010 : OUT <= 0;  //143 / 242 = 0
    16'b10001111_11110011 : OUT <= 0;  //143 / 243 = 0
    16'b10001111_11110100 : OUT <= 0;  //143 / 244 = 0
    16'b10001111_11110101 : OUT <= 0;  //143 / 245 = 0
    16'b10001111_11110110 : OUT <= 0;  //143 / 246 = 0
    16'b10001111_11110111 : OUT <= 0;  //143 / 247 = 0
    16'b10001111_11111000 : OUT <= 0;  //143 / 248 = 0
    16'b10001111_11111001 : OUT <= 0;  //143 / 249 = 0
    16'b10001111_11111010 : OUT <= 0;  //143 / 250 = 0
    16'b10001111_11111011 : OUT <= 0;  //143 / 251 = 0
    16'b10001111_11111100 : OUT <= 0;  //143 / 252 = 0
    16'b10001111_11111101 : OUT <= 0;  //143 / 253 = 0
    16'b10001111_11111110 : OUT <= 0;  //143 / 254 = 0
    16'b10001111_11111111 : OUT <= 0;  //143 / 255 = 0
    16'b10010000_00000000 : OUT <= 0;  //144 / 0 = 0
    16'b10010000_00000001 : OUT <= 144;  //144 / 1 = 144
    16'b10010000_00000010 : OUT <= 72;  //144 / 2 = 72
    16'b10010000_00000011 : OUT <= 48;  //144 / 3 = 48
    16'b10010000_00000100 : OUT <= 36;  //144 / 4 = 36
    16'b10010000_00000101 : OUT <= 28;  //144 / 5 = 28
    16'b10010000_00000110 : OUT <= 24;  //144 / 6 = 24
    16'b10010000_00000111 : OUT <= 20;  //144 / 7 = 20
    16'b10010000_00001000 : OUT <= 18;  //144 / 8 = 18
    16'b10010000_00001001 : OUT <= 16;  //144 / 9 = 16
    16'b10010000_00001010 : OUT <= 14;  //144 / 10 = 14
    16'b10010000_00001011 : OUT <= 13;  //144 / 11 = 13
    16'b10010000_00001100 : OUT <= 12;  //144 / 12 = 12
    16'b10010000_00001101 : OUT <= 11;  //144 / 13 = 11
    16'b10010000_00001110 : OUT <= 10;  //144 / 14 = 10
    16'b10010000_00001111 : OUT <= 9;  //144 / 15 = 9
    16'b10010000_00010000 : OUT <= 9;  //144 / 16 = 9
    16'b10010000_00010001 : OUT <= 8;  //144 / 17 = 8
    16'b10010000_00010010 : OUT <= 8;  //144 / 18 = 8
    16'b10010000_00010011 : OUT <= 7;  //144 / 19 = 7
    16'b10010000_00010100 : OUT <= 7;  //144 / 20 = 7
    16'b10010000_00010101 : OUT <= 6;  //144 / 21 = 6
    16'b10010000_00010110 : OUT <= 6;  //144 / 22 = 6
    16'b10010000_00010111 : OUT <= 6;  //144 / 23 = 6
    16'b10010000_00011000 : OUT <= 6;  //144 / 24 = 6
    16'b10010000_00011001 : OUT <= 5;  //144 / 25 = 5
    16'b10010000_00011010 : OUT <= 5;  //144 / 26 = 5
    16'b10010000_00011011 : OUT <= 5;  //144 / 27 = 5
    16'b10010000_00011100 : OUT <= 5;  //144 / 28 = 5
    16'b10010000_00011101 : OUT <= 4;  //144 / 29 = 4
    16'b10010000_00011110 : OUT <= 4;  //144 / 30 = 4
    16'b10010000_00011111 : OUT <= 4;  //144 / 31 = 4
    16'b10010000_00100000 : OUT <= 4;  //144 / 32 = 4
    16'b10010000_00100001 : OUT <= 4;  //144 / 33 = 4
    16'b10010000_00100010 : OUT <= 4;  //144 / 34 = 4
    16'b10010000_00100011 : OUT <= 4;  //144 / 35 = 4
    16'b10010000_00100100 : OUT <= 4;  //144 / 36 = 4
    16'b10010000_00100101 : OUT <= 3;  //144 / 37 = 3
    16'b10010000_00100110 : OUT <= 3;  //144 / 38 = 3
    16'b10010000_00100111 : OUT <= 3;  //144 / 39 = 3
    16'b10010000_00101000 : OUT <= 3;  //144 / 40 = 3
    16'b10010000_00101001 : OUT <= 3;  //144 / 41 = 3
    16'b10010000_00101010 : OUT <= 3;  //144 / 42 = 3
    16'b10010000_00101011 : OUT <= 3;  //144 / 43 = 3
    16'b10010000_00101100 : OUT <= 3;  //144 / 44 = 3
    16'b10010000_00101101 : OUT <= 3;  //144 / 45 = 3
    16'b10010000_00101110 : OUT <= 3;  //144 / 46 = 3
    16'b10010000_00101111 : OUT <= 3;  //144 / 47 = 3
    16'b10010000_00110000 : OUT <= 3;  //144 / 48 = 3
    16'b10010000_00110001 : OUT <= 2;  //144 / 49 = 2
    16'b10010000_00110010 : OUT <= 2;  //144 / 50 = 2
    16'b10010000_00110011 : OUT <= 2;  //144 / 51 = 2
    16'b10010000_00110100 : OUT <= 2;  //144 / 52 = 2
    16'b10010000_00110101 : OUT <= 2;  //144 / 53 = 2
    16'b10010000_00110110 : OUT <= 2;  //144 / 54 = 2
    16'b10010000_00110111 : OUT <= 2;  //144 / 55 = 2
    16'b10010000_00111000 : OUT <= 2;  //144 / 56 = 2
    16'b10010000_00111001 : OUT <= 2;  //144 / 57 = 2
    16'b10010000_00111010 : OUT <= 2;  //144 / 58 = 2
    16'b10010000_00111011 : OUT <= 2;  //144 / 59 = 2
    16'b10010000_00111100 : OUT <= 2;  //144 / 60 = 2
    16'b10010000_00111101 : OUT <= 2;  //144 / 61 = 2
    16'b10010000_00111110 : OUT <= 2;  //144 / 62 = 2
    16'b10010000_00111111 : OUT <= 2;  //144 / 63 = 2
    16'b10010000_01000000 : OUT <= 2;  //144 / 64 = 2
    16'b10010000_01000001 : OUT <= 2;  //144 / 65 = 2
    16'b10010000_01000010 : OUT <= 2;  //144 / 66 = 2
    16'b10010000_01000011 : OUT <= 2;  //144 / 67 = 2
    16'b10010000_01000100 : OUT <= 2;  //144 / 68 = 2
    16'b10010000_01000101 : OUT <= 2;  //144 / 69 = 2
    16'b10010000_01000110 : OUT <= 2;  //144 / 70 = 2
    16'b10010000_01000111 : OUT <= 2;  //144 / 71 = 2
    16'b10010000_01001000 : OUT <= 2;  //144 / 72 = 2
    16'b10010000_01001001 : OUT <= 1;  //144 / 73 = 1
    16'b10010000_01001010 : OUT <= 1;  //144 / 74 = 1
    16'b10010000_01001011 : OUT <= 1;  //144 / 75 = 1
    16'b10010000_01001100 : OUT <= 1;  //144 / 76 = 1
    16'b10010000_01001101 : OUT <= 1;  //144 / 77 = 1
    16'b10010000_01001110 : OUT <= 1;  //144 / 78 = 1
    16'b10010000_01001111 : OUT <= 1;  //144 / 79 = 1
    16'b10010000_01010000 : OUT <= 1;  //144 / 80 = 1
    16'b10010000_01010001 : OUT <= 1;  //144 / 81 = 1
    16'b10010000_01010010 : OUT <= 1;  //144 / 82 = 1
    16'b10010000_01010011 : OUT <= 1;  //144 / 83 = 1
    16'b10010000_01010100 : OUT <= 1;  //144 / 84 = 1
    16'b10010000_01010101 : OUT <= 1;  //144 / 85 = 1
    16'b10010000_01010110 : OUT <= 1;  //144 / 86 = 1
    16'b10010000_01010111 : OUT <= 1;  //144 / 87 = 1
    16'b10010000_01011000 : OUT <= 1;  //144 / 88 = 1
    16'b10010000_01011001 : OUT <= 1;  //144 / 89 = 1
    16'b10010000_01011010 : OUT <= 1;  //144 / 90 = 1
    16'b10010000_01011011 : OUT <= 1;  //144 / 91 = 1
    16'b10010000_01011100 : OUT <= 1;  //144 / 92 = 1
    16'b10010000_01011101 : OUT <= 1;  //144 / 93 = 1
    16'b10010000_01011110 : OUT <= 1;  //144 / 94 = 1
    16'b10010000_01011111 : OUT <= 1;  //144 / 95 = 1
    16'b10010000_01100000 : OUT <= 1;  //144 / 96 = 1
    16'b10010000_01100001 : OUT <= 1;  //144 / 97 = 1
    16'b10010000_01100010 : OUT <= 1;  //144 / 98 = 1
    16'b10010000_01100011 : OUT <= 1;  //144 / 99 = 1
    16'b10010000_01100100 : OUT <= 1;  //144 / 100 = 1
    16'b10010000_01100101 : OUT <= 1;  //144 / 101 = 1
    16'b10010000_01100110 : OUT <= 1;  //144 / 102 = 1
    16'b10010000_01100111 : OUT <= 1;  //144 / 103 = 1
    16'b10010000_01101000 : OUT <= 1;  //144 / 104 = 1
    16'b10010000_01101001 : OUT <= 1;  //144 / 105 = 1
    16'b10010000_01101010 : OUT <= 1;  //144 / 106 = 1
    16'b10010000_01101011 : OUT <= 1;  //144 / 107 = 1
    16'b10010000_01101100 : OUT <= 1;  //144 / 108 = 1
    16'b10010000_01101101 : OUT <= 1;  //144 / 109 = 1
    16'b10010000_01101110 : OUT <= 1;  //144 / 110 = 1
    16'b10010000_01101111 : OUT <= 1;  //144 / 111 = 1
    16'b10010000_01110000 : OUT <= 1;  //144 / 112 = 1
    16'b10010000_01110001 : OUT <= 1;  //144 / 113 = 1
    16'b10010000_01110010 : OUT <= 1;  //144 / 114 = 1
    16'b10010000_01110011 : OUT <= 1;  //144 / 115 = 1
    16'b10010000_01110100 : OUT <= 1;  //144 / 116 = 1
    16'b10010000_01110101 : OUT <= 1;  //144 / 117 = 1
    16'b10010000_01110110 : OUT <= 1;  //144 / 118 = 1
    16'b10010000_01110111 : OUT <= 1;  //144 / 119 = 1
    16'b10010000_01111000 : OUT <= 1;  //144 / 120 = 1
    16'b10010000_01111001 : OUT <= 1;  //144 / 121 = 1
    16'b10010000_01111010 : OUT <= 1;  //144 / 122 = 1
    16'b10010000_01111011 : OUT <= 1;  //144 / 123 = 1
    16'b10010000_01111100 : OUT <= 1;  //144 / 124 = 1
    16'b10010000_01111101 : OUT <= 1;  //144 / 125 = 1
    16'b10010000_01111110 : OUT <= 1;  //144 / 126 = 1
    16'b10010000_01111111 : OUT <= 1;  //144 / 127 = 1
    16'b10010000_10000000 : OUT <= 1;  //144 / 128 = 1
    16'b10010000_10000001 : OUT <= 1;  //144 / 129 = 1
    16'b10010000_10000010 : OUT <= 1;  //144 / 130 = 1
    16'b10010000_10000011 : OUT <= 1;  //144 / 131 = 1
    16'b10010000_10000100 : OUT <= 1;  //144 / 132 = 1
    16'b10010000_10000101 : OUT <= 1;  //144 / 133 = 1
    16'b10010000_10000110 : OUT <= 1;  //144 / 134 = 1
    16'b10010000_10000111 : OUT <= 1;  //144 / 135 = 1
    16'b10010000_10001000 : OUT <= 1;  //144 / 136 = 1
    16'b10010000_10001001 : OUT <= 1;  //144 / 137 = 1
    16'b10010000_10001010 : OUT <= 1;  //144 / 138 = 1
    16'b10010000_10001011 : OUT <= 1;  //144 / 139 = 1
    16'b10010000_10001100 : OUT <= 1;  //144 / 140 = 1
    16'b10010000_10001101 : OUT <= 1;  //144 / 141 = 1
    16'b10010000_10001110 : OUT <= 1;  //144 / 142 = 1
    16'b10010000_10001111 : OUT <= 1;  //144 / 143 = 1
    16'b10010000_10010000 : OUT <= 1;  //144 / 144 = 1
    16'b10010000_10010001 : OUT <= 0;  //144 / 145 = 0
    16'b10010000_10010010 : OUT <= 0;  //144 / 146 = 0
    16'b10010000_10010011 : OUT <= 0;  //144 / 147 = 0
    16'b10010000_10010100 : OUT <= 0;  //144 / 148 = 0
    16'b10010000_10010101 : OUT <= 0;  //144 / 149 = 0
    16'b10010000_10010110 : OUT <= 0;  //144 / 150 = 0
    16'b10010000_10010111 : OUT <= 0;  //144 / 151 = 0
    16'b10010000_10011000 : OUT <= 0;  //144 / 152 = 0
    16'b10010000_10011001 : OUT <= 0;  //144 / 153 = 0
    16'b10010000_10011010 : OUT <= 0;  //144 / 154 = 0
    16'b10010000_10011011 : OUT <= 0;  //144 / 155 = 0
    16'b10010000_10011100 : OUT <= 0;  //144 / 156 = 0
    16'b10010000_10011101 : OUT <= 0;  //144 / 157 = 0
    16'b10010000_10011110 : OUT <= 0;  //144 / 158 = 0
    16'b10010000_10011111 : OUT <= 0;  //144 / 159 = 0
    16'b10010000_10100000 : OUT <= 0;  //144 / 160 = 0
    16'b10010000_10100001 : OUT <= 0;  //144 / 161 = 0
    16'b10010000_10100010 : OUT <= 0;  //144 / 162 = 0
    16'b10010000_10100011 : OUT <= 0;  //144 / 163 = 0
    16'b10010000_10100100 : OUT <= 0;  //144 / 164 = 0
    16'b10010000_10100101 : OUT <= 0;  //144 / 165 = 0
    16'b10010000_10100110 : OUT <= 0;  //144 / 166 = 0
    16'b10010000_10100111 : OUT <= 0;  //144 / 167 = 0
    16'b10010000_10101000 : OUT <= 0;  //144 / 168 = 0
    16'b10010000_10101001 : OUT <= 0;  //144 / 169 = 0
    16'b10010000_10101010 : OUT <= 0;  //144 / 170 = 0
    16'b10010000_10101011 : OUT <= 0;  //144 / 171 = 0
    16'b10010000_10101100 : OUT <= 0;  //144 / 172 = 0
    16'b10010000_10101101 : OUT <= 0;  //144 / 173 = 0
    16'b10010000_10101110 : OUT <= 0;  //144 / 174 = 0
    16'b10010000_10101111 : OUT <= 0;  //144 / 175 = 0
    16'b10010000_10110000 : OUT <= 0;  //144 / 176 = 0
    16'b10010000_10110001 : OUT <= 0;  //144 / 177 = 0
    16'b10010000_10110010 : OUT <= 0;  //144 / 178 = 0
    16'b10010000_10110011 : OUT <= 0;  //144 / 179 = 0
    16'b10010000_10110100 : OUT <= 0;  //144 / 180 = 0
    16'b10010000_10110101 : OUT <= 0;  //144 / 181 = 0
    16'b10010000_10110110 : OUT <= 0;  //144 / 182 = 0
    16'b10010000_10110111 : OUT <= 0;  //144 / 183 = 0
    16'b10010000_10111000 : OUT <= 0;  //144 / 184 = 0
    16'b10010000_10111001 : OUT <= 0;  //144 / 185 = 0
    16'b10010000_10111010 : OUT <= 0;  //144 / 186 = 0
    16'b10010000_10111011 : OUT <= 0;  //144 / 187 = 0
    16'b10010000_10111100 : OUT <= 0;  //144 / 188 = 0
    16'b10010000_10111101 : OUT <= 0;  //144 / 189 = 0
    16'b10010000_10111110 : OUT <= 0;  //144 / 190 = 0
    16'b10010000_10111111 : OUT <= 0;  //144 / 191 = 0
    16'b10010000_11000000 : OUT <= 0;  //144 / 192 = 0
    16'b10010000_11000001 : OUT <= 0;  //144 / 193 = 0
    16'b10010000_11000010 : OUT <= 0;  //144 / 194 = 0
    16'b10010000_11000011 : OUT <= 0;  //144 / 195 = 0
    16'b10010000_11000100 : OUT <= 0;  //144 / 196 = 0
    16'b10010000_11000101 : OUT <= 0;  //144 / 197 = 0
    16'b10010000_11000110 : OUT <= 0;  //144 / 198 = 0
    16'b10010000_11000111 : OUT <= 0;  //144 / 199 = 0
    16'b10010000_11001000 : OUT <= 0;  //144 / 200 = 0
    16'b10010000_11001001 : OUT <= 0;  //144 / 201 = 0
    16'b10010000_11001010 : OUT <= 0;  //144 / 202 = 0
    16'b10010000_11001011 : OUT <= 0;  //144 / 203 = 0
    16'b10010000_11001100 : OUT <= 0;  //144 / 204 = 0
    16'b10010000_11001101 : OUT <= 0;  //144 / 205 = 0
    16'b10010000_11001110 : OUT <= 0;  //144 / 206 = 0
    16'b10010000_11001111 : OUT <= 0;  //144 / 207 = 0
    16'b10010000_11010000 : OUT <= 0;  //144 / 208 = 0
    16'b10010000_11010001 : OUT <= 0;  //144 / 209 = 0
    16'b10010000_11010010 : OUT <= 0;  //144 / 210 = 0
    16'b10010000_11010011 : OUT <= 0;  //144 / 211 = 0
    16'b10010000_11010100 : OUT <= 0;  //144 / 212 = 0
    16'b10010000_11010101 : OUT <= 0;  //144 / 213 = 0
    16'b10010000_11010110 : OUT <= 0;  //144 / 214 = 0
    16'b10010000_11010111 : OUT <= 0;  //144 / 215 = 0
    16'b10010000_11011000 : OUT <= 0;  //144 / 216 = 0
    16'b10010000_11011001 : OUT <= 0;  //144 / 217 = 0
    16'b10010000_11011010 : OUT <= 0;  //144 / 218 = 0
    16'b10010000_11011011 : OUT <= 0;  //144 / 219 = 0
    16'b10010000_11011100 : OUT <= 0;  //144 / 220 = 0
    16'b10010000_11011101 : OUT <= 0;  //144 / 221 = 0
    16'b10010000_11011110 : OUT <= 0;  //144 / 222 = 0
    16'b10010000_11011111 : OUT <= 0;  //144 / 223 = 0
    16'b10010000_11100000 : OUT <= 0;  //144 / 224 = 0
    16'b10010000_11100001 : OUT <= 0;  //144 / 225 = 0
    16'b10010000_11100010 : OUT <= 0;  //144 / 226 = 0
    16'b10010000_11100011 : OUT <= 0;  //144 / 227 = 0
    16'b10010000_11100100 : OUT <= 0;  //144 / 228 = 0
    16'b10010000_11100101 : OUT <= 0;  //144 / 229 = 0
    16'b10010000_11100110 : OUT <= 0;  //144 / 230 = 0
    16'b10010000_11100111 : OUT <= 0;  //144 / 231 = 0
    16'b10010000_11101000 : OUT <= 0;  //144 / 232 = 0
    16'b10010000_11101001 : OUT <= 0;  //144 / 233 = 0
    16'b10010000_11101010 : OUT <= 0;  //144 / 234 = 0
    16'b10010000_11101011 : OUT <= 0;  //144 / 235 = 0
    16'b10010000_11101100 : OUT <= 0;  //144 / 236 = 0
    16'b10010000_11101101 : OUT <= 0;  //144 / 237 = 0
    16'b10010000_11101110 : OUT <= 0;  //144 / 238 = 0
    16'b10010000_11101111 : OUT <= 0;  //144 / 239 = 0
    16'b10010000_11110000 : OUT <= 0;  //144 / 240 = 0
    16'b10010000_11110001 : OUT <= 0;  //144 / 241 = 0
    16'b10010000_11110010 : OUT <= 0;  //144 / 242 = 0
    16'b10010000_11110011 : OUT <= 0;  //144 / 243 = 0
    16'b10010000_11110100 : OUT <= 0;  //144 / 244 = 0
    16'b10010000_11110101 : OUT <= 0;  //144 / 245 = 0
    16'b10010000_11110110 : OUT <= 0;  //144 / 246 = 0
    16'b10010000_11110111 : OUT <= 0;  //144 / 247 = 0
    16'b10010000_11111000 : OUT <= 0;  //144 / 248 = 0
    16'b10010000_11111001 : OUT <= 0;  //144 / 249 = 0
    16'b10010000_11111010 : OUT <= 0;  //144 / 250 = 0
    16'b10010000_11111011 : OUT <= 0;  //144 / 251 = 0
    16'b10010000_11111100 : OUT <= 0;  //144 / 252 = 0
    16'b10010000_11111101 : OUT <= 0;  //144 / 253 = 0
    16'b10010000_11111110 : OUT <= 0;  //144 / 254 = 0
    16'b10010000_11111111 : OUT <= 0;  //144 / 255 = 0
    16'b10010001_00000000 : OUT <= 0;  //145 / 0 = 0
    16'b10010001_00000001 : OUT <= 145;  //145 / 1 = 145
    16'b10010001_00000010 : OUT <= 72;  //145 / 2 = 72
    16'b10010001_00000011 : OUT <= 48;  //145 / 3 = 48
    16'b10010001_00000100 : OUT <= 36;  //145 / 4 = 36
    16'b10010001_00000101 : OUT <= 29;  //145 / 5 = 29
    16'b10010001_00000110 : OUT <= 24;  //145 / 6 = 24
    16'b10010001_00000111 : OUT <= 20;  //145 / 7 = 20
    16'b10010001_00001000 : OUT <= 18;  //145 / 8 = 18
    16'b10010001_00001001 : OUT <= 16;  //145 / 9 = 16
    16'b10010001_00001010 : OUT <= 14;  //145 / 10 = 14
    16'b10010001_00001011 : OUT <= 13;  //145 / 11 = 13
    16'b10010001_00001100 : OUT <= 12;  //145 / 12 = 12
    16'b10010001_00001101 : OUT <= 11;  //145 / 13 = 11
    16'b10010001_00001110 : OUT <= 10;  //145 / 14 = 10
    16'b10010001_00001111 : OUT <= 9;  //145 / 15 = 9
    16'b10010001_00010000 : OUT <= 9;  //145 / 16 = 9
    16'b10010001_00010001 : OUT <= 8;  //145 / 17 = 8
    16'b10010001_00010010 : OUT <= 8;  //145 / 18 = 8
    16'b10010001_00010011 : OUT <= 7;  //145 / 19 = 7
    16'b10010001_00010100 : OUT <= 7;  //145 / 20 = 7
    16'b10010001_00010101 : OUT <= 6;  //145 / 21 = 6
    16'b10010001_00010110 : OUT <= 6;  //145 / 22 = 6
    16'b10010001_00010111 : OUT <= 6;  //145 / 23 = 6
    16'b10010001_00011000 : OUT <= 6;  //145 / 24 = 6
    16'b10010001_00011001 : OUT <= 5;  //145 / 25 = 5
    16'b10010001_00011010 : OUT <= 5;  //145 / 26 = 5
    16'b10010001_00011011 : OUT <= 5;  //145 / 27 = 5
    16'b10010001_00011100 : OUT <= 5;  //145 / 28 = 5
    16'b10010001_00011101 : OUT <= 5;  //145 / 29 = 5
    16'b10010001_00011110 : OUT <= 4;  //145 / 30 = 4
    16'b10010001_00011111 : OUT <= 4;  //145 / 31 = 4
    16'b10010001_00100000 : OUT <= 4;  //145 / 32 = 4
    16'b10010001_00100001 : OUT <= 4;  //145 / 33 = 4
    16'b10010001_00100010 : OUT <= 4;  //145 / 34 = 4
    16'b10010001_00100011 : OUT <= 4;  //145 / 35 = 4
    16'b10010001_00100100 : OUT <= 4;  //145 / 36 = 4
    16'b10010001_00100101 : OUT <= 3;  //145 / 37 = 3
    16'b10010001_00100110 : OUT <= 3;  //145 / 38 = 3
    16'b10010001_00100111 : OUT <= 3;  //145 / 39 = 3
    16'b10010001_00101000 : OUT <= 3;  //145 / 40 = 3
    16'b10010001_00101001 : OUT <= 3;  //145 / 41 = 3
    16'b10010001_00101010 : OUT <= 3;  //145 / 42 = 3
    16'b10010001_00101011 : OUT <= 3;  //145 / 43 = 3
    16'b10010001_00101100 : OUT <= 3;  //145 / 44 = 3
    16'b10010001_00101101 : OUT <= 3;  //145 / 45 = 3
    16'b10010001_00101110 : OUT <= 3;  //145 / 46 = 3
    16'b10010001_00101111 : OUT <= 3;  //145 / 47 = 3
    16'b10010001_00110000 : OUT <= 3;  //145 / 48 = 3
    16'b10010001_00110001 : OUT <= 2;  //145 / 49 = 2
    16'b10010001_00110010 : OUT <= 2;  //145 / 50 = 2
    16'b10010001_00110011 : OUT <= 2;  //145 / 51 = 2
    16'b10010001_00110100 : OUT <= 2;  //145 / 52 = 2
    16'b10010001_00110101 : OUT <= 2;  //145 / 53 = 2
    16'b10010001_00110110 : OUT <= 2;  //145 / 54 = 2
    16'b10010001_00110111 : OUT <= 2;  //145 / 55 = 2
    16'b10010001_00111000 : OUT <= 2;  //145 / 56 = 2
    16'b10010001_00111001 : OUT <= 2;  //145 / 57 = 2
    16'b10010001_00111010 : OUT <= 2;  //145 / 58 = 2
    16'b10010001_00111011 : OUT <= 2;  //145 / 59 = 2
    16'b10010001_00111100 : OUT <= 2;  //145 / 60 = 2
    16'b10010001_00111101 : OUT <= 2;  //145 / 61 = 2
    16'b10010001_00111110 : OUT <= 2;  //145 / 62 = 2
    16'b10010001_00111111 : OUT <= 2;  //145 / 63 = 2
    16'b10010001_01000000 : OUT <= 2;  //145 / 64 = 2
    16'b10010001_01000001 : OUT <= 2;  //145 / 65 = 2
    16'b10010001_01000010 : OUT <= 2;  //145 / 66 = 2
    16'b10010001_01000011 : OUT <= 2;  //145 / 67 = 2
    16'b10010001_01000100 : OUT <= 2;  //145 / 68 = 2
    16'b10010001_01000101 : OUT <= 2;  //145 / 69 = 2
    16'b10010001_01000110 : OUT <= 2;  //145 / 70 = 2
    16'b10010001_01000111 : OUT <= 2;  //145 / 71 = 2
    16'b10010001_01001000 : OUT <= 2;  //145 / 72 = 2
    16'b10010001_01001001 : OUT <= 1;  //145 / 73 = 1
    16'b10010001_01001010 : OUT <= 1;  //145 / 74 = 1
    16'b10010001_01001011 : OUT <= 1;  //145 / 75 = 1
    16'b10010001_01001100 : OUT <= 1;  //145 / 76 = 1
    16'b10010001_01001101 : OUT <= 1;  //145 / 77 = 1
    16'b10010001_01001110 : OUT <= 1;  //145 / 78 = 1
    16'b10010001_01001111 : OUT <= 1;  //145 / 79 = 1
    16'b10010001_01010000 : OUT <= 1;  //145 / 80 = 1
    16'b10010001_01010001 : OUT <= 1;  //145 / 81 = 1
    16'b10010001_01010010 : OUT <= 1;  //145 / 82 = 1
    16'b10010001_01010011 : OUT <= 1;  //145 / 83 = 1
    16'b10010001_01010100 : OUT <= 1;  //145 / 84 = 1
    16'b10010001_01010101 : OUT <= 1;  //145 / 85 = 1
    16'b10010001_01010110 : OUT <= 1;  //145 / 86 = 1
    16'b10010001_01010111 : OUT <= 1;  //145 / 87 = 1
    16'b10010001_01011000 : OUT <= 1;  //145 / 88 = 1
    16'b10010001_01011001 : OUT <= 1;  //145 / 89 = 1
    16'b10010001_01011010 : OUT <= 1;  //145 / 90 = 1
    16'b10010001_01011011 : OUT <= 1;  //145 / 91 = 1
    16'b10010001_01011100 : OUT <= 1;  //145 / 92 = 1
    16'b10010001_01011101 : OUT <= 1;  //145 / 93 = 1
    16'b10010001_01011110 : OUT <= 1;  //145 / 94 = 1
    16'b10010001_01011111 : OUT <= 1;  //145 / 95 = 1
    16'b10010001_01100000 : OUT <= 1;  //145 / 96 = 1
    16'b10010001_01100001 : OUT <= 1;  //145 / 97 = 1
    16'b10010001_01100010 : OUT <= 1;  //145 / 98 = 1
    16'b10010001_01100011 : OUT <= 1;  //145 / 99 = 1
    16'b10010001_01100100 : OUT <= 1;  //145 / 100 = 1
    16'b10010001_01100101 : OUT <= 1;  //145 / 101 = 1
    16'b10010001_01100110 : OUT <= 1;  //145 / 102 = 1
    16'b10010001_01100111 : OUT <= 1;  //145 / 103 = 1
    16'b10010001_01101000 : OUT <= 1;  //145 / 104 = 1
    16'b10010001_01101001 : OUT <= 1;  //145 / 105 = 1
    16'b10010001_01101010 : OUT <= 1;  //145 / 106 = 1
    16'b10010001_01101011 : OUT <= 1;  //145 / 107 = 1
    16'b10010001_01101100 : OUT <= 1;  //145 / 108 = 1
    16'b10010001_01101101 : OUT <= 1;  //145 / 109 = 1
    16'b10010001_01101110 : OUT <= 1;  //145 / 110 = 1
    16'b10010001_01101111 : OUT <= 1;  //145 / 111 = 1
    16'b10010001_01110000 : OUT <= 1;  //145 / 112 = 1
    16'b10010001_01110001 : OUT <= 1;  //145 / 113 = 1
    16'b10010001_01110010 : OUT <= 1;  //145 / 114 = 1
    16'b10010001_01110011 : OUT <= 1;  //145 / 115 = 1
    16'b10010001_01110100 : OUT <= 1;  //145 / 116 = 1
    16'b10010001_01110101 : OUT <= 1;  //145 / 117 = 1
    16'b10010001_01110110 : OUT <= 1;  //145 / 118 = 1
    16'b10010001_01110111 : OUT <= 1;  //145 / 119 = 1
    16'b10010001_01111000 : OUT <= 1;  //145 / 120 = 1
    16'b10010001_01111001 : OUT <= 1;  //145 / 121 = 1
    16'b10010001_01111010 : OUT <= 1;  //145 / 122 = 1
    16'b10010001_01111011 : OUT <= 1;  //145 / 123 = 1
    16'b10010001_01111100 : OUT <= 1;  //145 / 124 = 1
    16'b10010001_01111101 : OUT <= 1;  //145 / 125 = 1
    16'b10010001_01111110 : OUT <= 1;  //145 / 126 = 1
    16'b10010001_01111111 : OUT <= 1;  //145 / 127 = 1
    16'b10010001_10000000 : OUT <= 1;  //145 / 128 = 1
    16'b10010001_10000001 : OUT <= 1;  //145 / 129 = 1
    16'b10010001_10000010 : OUT <= 1;  //145 / 130 = 1
    16'b10010001_10000011 : OUT <= 1;  //145 / 131 = 1
    16'b10010001_10000100 : OUT <= 1;  //145 / 132 = 1
    16'b10010001_10000101 : OUT <= 1;  //145 / 133 = 1
    16'b10010001_10000110 : OUT <= 1;  //145 / 134 = 1
    16'b10010001_10000111 : OUT <= 1;  //145 / 135 = 1
    16'b10010001_10001000 : OUT <= 1;  //145 / 136 = 1
    16'b10010001_10001001 : OUT <= 1;  //145 / 137 = 1
    16'b10010001_10001010 : OUT <= 1;  //145 / 138 = 1
    16'b10010001_10001011 : OUT <= 1;  //145 / 139 = 1
    16'b10010001_10001100 : OUT <= 1;  //145 / 140 = 1
    16'b10010001_10001101 : OUT <= 1;  //145 / 141 = 1
    16'b10010001_10001110 : OUT <= 1;  //145 / 142 = 1
    16'b10010001_10001111 : OUT <= 1;  //145 / 143 = 1
    16'b10010001_10010000 : OUT <= 1;  //145 / 144 = 1
    16'b10010001_10010001 : OUT <= 1;  //145 / 145 = 1
    16'b10010001_10010010 : OUT <= 0;  //145 / 146 = 0
    16'b10010001_10010011 : OUT <= 0;  //145 / 147 = 0
    16'b10010001_10010100 : OUT <= 0;  //145 / 148 = 0
    16'b10010001_10010101 : OUT <= 0;  //145 / 149 = 0
    16'b10010001_10010110 : OUT <= 0;  //145 / 150 = 0
    16'b10010001_10010111 : OUT <= 0;  //145 / 151 = 0
    16'b10010001_10011000 : OUT <= 0;  //145 / 152 = 0
    16'b10010001_10011001 : OUT <= 0;  //145 / 153 = 0
    16'b10010001_10011010 : OUT <= 0;  //145 / 154 = 0
    16'b10010001_10011011 : OUT <= 0;  //145 / 155 = 0
    16'b10010001_10011100 : OUT <= 0;  //145 / 156 = 0
    16'b10010001_10011101 : OUT <= 0;  //145 / 157 = 0
    16'b10010001_10011110 : OUT <= 0;  //145 / 158 = 0
    16'b10010001_10011111 : OUT <= 0;  //145 / 159 = 0
    16'b10010001_10100000 : OUT <= 0;  //145 / 160 = 0
    16'b10010001_10100001 : OUT <= 0;  //145 / 161 = 0
    16'b10010001_10100010 : OUT <= 0;  //145 / 162 = 0
    16'b10010001_10100011 : OUT <= 0;  //145 / 163 = 0
    16'b10010001_10100100 : OUT <= 0;  //145 / 164 = 0
    16'b10010001_10100101 : OUT <= 0;  //145 / 165 = 0
    16'b10010001_10100110 : OUT <= 0;  //145 / 166 = 0
    16'b10010001_10100111 : OUT <= 0;  //145 / 167 = 0
    16'b10010001_10101000 : OUT <= 0;  //145 / 168 = 0
    16'b10010001_10101001 : OUT <= 0;  //145 / 169 = 0
    16'b10010001_10101010 : OUT <= 0;  //145 / 170 = 0
    16'b10010001_10101011 : OUT <= 0;  //145 / 171 = 0
    16'b10010001_10101100 : OUT <= 0;  //145 / 172 = 0
    16'b10010001_10101101 : OUT <= 0;  //145 / 173 = 0
    16'b10010001_10101110 : OUT <= 0;  //145 / 174 = 0
    16'b10010001_10101111 : OUT <= 0;  //145 / 175 = 0
    16'b10010001_10110000 : OUT <= 0;  //145 / 176 = 0
    16'b10010001_10110001 : OUT <= 0;  //145 / 177 = 0
    16'b10010001_10110010 : OUT <= 0;  //145 / 178 = 0
    16'b10010001_10110011 : OUT <= 0;  //145 / 179 = 0
    16'b10010001_10110100 : OUT <= 0;  //145 / 180 = 0
    16'b10010001_10110101 : OUT <= 0;  //145 / 181 = 0
    16'b10010001_10110110 : OUT <= 0;  //145 / 182 = 0
    16'b10010001_10110111 : OUT <= 0;  //145 / 183 = 0
    16'b10010001_10111000 : OUT <= 0;  //145 / 184 = 0
    16'b10010001_10111001 : OUT <= 0;  //145 / 185 = 0
    16'b10010001_10111010 : OUT <= 0;  //145 / 186 = 0
    16'b10010001_10111011 : OUT <= 0;  //145 / 187 = 0
    16'b10010001_10111100 : OUT <= 0;  //145 / 188 = 0
    16'b10010001_10111101 : OUT <= 0;  //145 / 189 = 0
    16'b10010001_10111110 : OUT <= 0;  //145 / 190 = 0
    16'b10010001_10111111 : OUT <= 0;  //145 / 191 = 0
    16'b10010001_11000000 : OUT <= 0;  //145 / 192 = 0
    16'b10010001_11000001 : OUT <= 0;  //145 / 193 = 0
    16'b10010001_11000010 : OUT <= 0;  //145 / 194 = 0
    16'b10010001_11000011 : OUT <= 0;  //145 / 195 = 0
    16'b10010001_11000100 : OUT <= 0;  //145 / 196 = 0
    16'b10010001_11000101 : OUT <= 0;  //145 / 197 = 0
    16'b10010001_11000110 : OUT <= 0;  //145 / 198 = 0
    16'b10010001_11000111 : OUT <= 0;  //145 / 199 = 0
    16'b10010001_11001000 : OUT <= 0;  //145 / 200 = 0
    16'b10010001_11001001 : OUT <= 0;  //145 / 201 = 0
    16'b10010001_11001010 : OUT <= 0;  //145 / 202 = 0
    16'b10010001_11001011 : OUT <= 0;  //145 / 203 = 0
    16'b10010001_11001100 : OUT <= 0;  //145 / 204 = 0
    16'b10010001_11001101 : OUT <= 0;  //145 / 205 = 0
    16'b10010001_11001110 : OUT <= 0;  //145 / 206 = 0
    16'b10010001_11001111 : OUT <= 0;  //145 / 207 = 0
    16'b10010001_11010000 : OUT <= 0;  //145 / 208 = 0
    16'b10010001_11010001 : OUT <= 0;  //145 / 209 = 0
    16'b10010001_11010010 : OUT <= 0;  //145 / 210 = 0
    16'b10010001_11010011 : OUT <= 0;  //145 / 211 = 0
    16'b10010001_11010100 : OUT <= 0;  //145 / 212 = 0
    16'b10010001_11010101 : OUT <= 0;  //145 / 213 = 0
    16'b10010001_11010110 : OUT <= 0;  //145 / 214 = 0
    16'b10010001_11010111 : OUT <= 0;  //145 / 215 = 0
    16'b10010001_11011000 : OUT <= 0;  //145 / 216 = 0
    16'b10010001_11011001 : OUT <= 0;  //145 / 217 = 0
    16'b10010001_11011010 : OUT <= 0;  //145 / 218 = 0
    16'b10010001_11011011 : OUT <= 0;  //145 / 219 = 0
    16'b10010001_11011100 : OUT <= 0;  //145 / 220 = 0
    16'b10010001_11011101 : OUT <= 0;  //145 / 221 = 0
    16'b10010001_11011110 : OUT <= 0;  //145 / 222 = 0
    16'b10010001_11011111 : OUT <= 0;  //145 / 223 = 0
    16'b10010001_11100000 : OUT <= 0;  //145 / 224 = 0
    16'b10010001_11100001 : OUT <= 0;  //145 / 225 = 0
    16'b10010001_11100010 : OUT <= 0;  //145 / 226 = 0
    16'b10010001_11100011 : OUT <= 0;  //145 / 227 = 0
    16'b10010001_11100100 : OUT <= 0;  //145 / 228 = 0
    16'b10010001_11100101 : OUT <= 0;  //145 / 229 = 0
    16'b10010001_11100110 : OUT <= 0;  //145 / 230 = 0
    16'b10010001_11100111 : OUT <= 0;  //145 / 231 = 0
    16'b10010001_11101000 : OUT <= 0;  //145 / 232 = 0
    16'b10010001_11101001 : OUT <= 0;  //145 / 233 = 0
    16'b10010001_11101010 : OUT <= 0;  //145 / 234 = 0
    16'b10010001_11101011 : OUT <= 0;  //145 / 235 = 0
    16'b10010001_11101100 : OUT <= 0;  //145 / 236 = 0
    16'b10010001_11101101 : OUT <= 0;  //145 / 237 = 0
    16'b10010001_11101110 : OUT <= 0;  //145 / 238 = 0
    16'b10010001_11101111 : OUT <= 0;  //145 / 239 = 0
    16'b10010001_11110000 : OUT <= 0;  //145 / 240 = 0
    16'b10010001_11110001 : OUT <= 0;  //145 / 241 = 0
    16'b10010001_11110010 : OUT <= 0;  //145 / 242 = 0
    16'b10010001_11110011 : OUT <= 0;  //145 / 243 = 0
    16'b10010001_11110100 : OUT <= 0;  //145 / 244 = 0
    16'b10010001_11110101 : OUT <= 0;  //145 / 245 = 0
    16'b10010001_11110110 : OUT <= 0;  //145 / 246 = 0
    16'b10010001_11110111 : OUT <= 0;  //145 / 247 = 0
    16'b10010001_11111000 : OUT <= 0;  //145 / 248 = 0
    16'b10010001_11111001 : OUT <= 0;  //145 / 249 = 0
    16'b10010001_11111010 : OUT <= 0;  //145 / 250 = 0
    16'b10010001_11111011 : OUT <= 0;  //145 / 251 = 0
    16'b10010001_11111100 : OUT <= 0;  //145 / 252 = 0
    16'b10010001_11111101 : OUT <= 0;  //145 / 253 = 0
    16'b10010001_11111110 : OUT <= 0;  //145 / 254 = 0
    16'b10010001_11111111 : OUT <= 0;  //145 / 255 = 0
    16'b10010010_00000000 : OUT <= 0;  //146 / 0 = 0
    16'b10010010_00000001 : OUT <= 146;  //146 / 1 = 146
    16'b10010010_00000010 : OUT <= 73;  //146 / 2 = 73
    16'b10010010_00000011 : OUT <= 48;  //146 / 3 = 48
    16'b10010010_00000100 : OUT <= 36;  //146 / 4 = 36
    16'b10010010_00000101 : OUT <= 29;  //146 / 5 = 29
    16'b10010010_00000110 : OUT <= 24;  //146 / 6 = 24
    16'b10010010_00000111 : OUT <= 20;  //146 / 7 = 20
    16'b10010010_00001000 : OUT <= 18;  //146 / 8 = 18
    16'b10010010_00001001 : OUT <= 16;  //146 / 9 = 16
    16'b10010010_00001010 : OUT <= 14;  //146 / 10 = 14
    16'b10010010_00001011 : OUT <= 13;  //146 / 11 = 13
    16'b10010010_00001100 : OUT <= 12;  //146 / 12 = 12
    16'b10010010_00001101 : OUT <= 11;  //146 / 13 = 11
    16'b10010010_00001110 : OUT <= 10;  //146 / 14 = 10
    16'b10010010_00001111 : OUT <= 9;  //146 / 15 = 9
    16'b10010010_00010000 : OUT <= 9;  //146 / 16 = 9
    16'b10010010_00010001 : OUT <= 8;  //146 / 17 = 8
    16'b10010010_00010010 : OUT <= 8;  //146 / 18 = 8
    16'b10010010_00010011 : OUT <= 7;  //146 / 19 = 7
    16'b10010010_00010100 : OUT <= 7;  //146 / 20 = 7
    16'b10010010_00010101 : OUT <= 6;  //146 / 21 = 6
    16'b10010010_00010110 : OUT <= 6;  //146 / 22 = 6
    16'b10010010_00010111 : OUT <= 6;  //146 / 23 = 6
    16'b10010010_00011000 : OUT <= 6;  //146 / 24 = 6
    16'b10010010_00011001 : OUT <= 5;  //146 / 25 = 5
    16'b10010010_00011010 : OUT <= 5;  //146 / 26 = 5
    16'b10010010_00011011 : OUT <= 5;  //146 / 27 = 5
    16'b10010010_00011100 : OUT <= 5;  //146 / 28 = 5
    16'b10010010_00011101 : OUT <= 5;  //146 / 29 = 5
    16'b10010010_00011110 : OUT <= 4;  //146 / 30 = 4
    16'b10010010_00011111 : OUT <= 4;  //146 / 31 = 4
    16'b10010010_00100000 : OUT <= 4;  //146 / 32 = 4
    16'b10010010_00100001 : OUT <= 4;  //146 / 33 = 4
    16'b10010010_00100010 : OUT <= 4;  //146 / 34 = 4
    16'b10010010_00100011 : OUT <= 4;  //146 / 35 = 4
    16'b10010010_00100100 : OUT <= 4;  //146 / 36 = 4
    16'b10010010_00100101 : OUT <= 3;  //146 / 37 = 3
    16'b10010010_00100110 : OUT <= 3;  //146 / 38 = 3
    16'b10010010_00100111 : OUT <= 3;  //146 / 39 = 3
    16'b10010010_00101000 : OUT <= 3;  //146 / 40 = 3
    16'b10010010_00101001 : OUT <= 3;  //146 / 41 = 3
    16'b10010010_00101010 : OUT <= 3;  //146 / 42 = 3
    16'b10010010_00101011 : OUT <= 3;  //146 / 43 = 3
    16'b10010010_00101100 : OUT <= 3;  //146 / 44 = 3
    16'b10010010_00101101 : OUT <= 3;  //146 / 45 = 3
    16'b10010010_00101110 : OUT <= 3;  //146 / 46 = 3
    16'b10010010_00101111 : OUT <= 3;  //146 / 47 = 3
    16'b10010010_00110000 : OUT <= 3;  //146 / 48 = 3
    16'b10010010_00110001 : OUT <= 2;  //146 / 49 = 2
    16'b10010010_00110010 : OUT <= 2;  //146 / 50 = 2
    16'b10010010_00110011 : OUT <= 2;  //146 / 51 = 2
    16'b10010010_00110100 : OUT <= 2;  //146 / 52 = 2
    16'b10010010_00110101 : OUT <= 2;  //146 / 53 = 2
    16'b10010010_00110110 : OUT <= 2;  //146 / 54 = 2
    16'b10010010_00110111 : OUT <= 2;  //146 / 55 = 2
    16'b10010010_00111000 : OUT <= 2;  //146 / 56 = 2
    16'b10010010_00111001 : OUT <= 2;  //146 / 57 = 2
    16'b10010010_00111010 : OUT <= 2;  //146 / 58 = 2
    16'b10010010_00111011 : OUT <= 2;  //146 / 59 = 2
    16'b10010010_00111100 : OUT <= 2;  //146 / 60 = 2
    16'b10010010_00111101 : OUT <= 2;  //146 / 61 = 2
    16'b10010010_00111110 : OUT <= 2;  //146 / 62 = 2
    16'b10010010_00111111 : OUT <= 2;  //146 / 63 = 2
    16'b10010010_01000000 : OUT <= 2;  //146 / 64 = 2
    16'b10010010_01000001 : OUT <= 2;  //146 / 65 = 2
    16'b10010010_01000010 : OUT <= 2;  //146 / 66 = 2
    16'b10010010_01000011 : OUT <= 2;  //146 / 67 = 2
    16'b10010010_01000100 : OUT <= 2;  //146 / 68 = 2
    16'b10010010_01000101 : OUT <= 2;  //146 / 69 = 2
    16'b10010010_01000110 : OUT <= 2;  //146 / 70 = 2
    16'b10010010_01000111 : OUT <= 2;  //146 / 71 = 2
    16'b10010010_01001000 : OUT <= 2;  //146 / 72 = 2
    16'b10010010_01001001 : OUT <= 2;  //146 / 73 = 2
    16'b10010010_01001010 : OUT <= 1;  //146 / 74 = 1
    16'b10010010_01001011 : OUT <= 1;  //146 / 75 = 1
    16'b10010010_01001100 : OUT <= 1;  //146 / 76 = 1
    16'b10010010_01001101 : OUT <= 1;  //146 / 77 = 1
    16'b10010010_01001110 : OUT <= 1;  //146 / 78 = 1
    16'b10010010_01001111 : OUT <= 1;  //146 / 79 = 1
    16'b10010010_01010000 : OUT <= 1;  //146 / 80 = 1
    16'b10010010_01010001 : OUT <= 1;  //146 / 81 = 1
    16'b10010010_01010010 : OUT <= 1;  //146 / 82 = 1
    16'b10010010_01010011 : OUT <= 1;  //146 / 83 = 1
    16'b10010010_01010100 : OUT <= 1;  //146 / 84 = 1
    16'b10010010_01010101 : OUT <= 1;  //146 / 85 = 1
    16'b10010010_01010110 : OUT <= 1;  //146 / 86 = 1
    16'b10010010_01010111 : OUT <= 1;  //146 / 87 = 1
    16'b10010010_01011000 : OUT <= 1;  //146 / 88 = 1
    16'b10010010_01011001 : OUT <= 1;  //146 / 89 = 1
    16'b10010010_01011010 : OUT <= 1;  //146 / 90 = 1
    16'b10010010_01011011 : OUT <= 1;  //146 / 91 = 1
    16'b10010010_01011100 : OUT <= 1;  //146 / 92 = 1
    16'b10010010_01011101 : OUT <= 1;  //146 / 93 = 1
    16'b10010010_01011110 : OUT <= 1;  //146 / 94 = 1
    16'b10010010_01011111 : OUT <= 1;  //146 / 95 = 1
    16'b10010010_01100000 : OUT <= 1;  //146 / 96 = 1
    16'b10010010_01100001 : OUT <= 1;  //146 / 97 = 1
    16'b10010010_01100010 : OUT <= 1;  //146 / 98 = 1
    16'b10010010_01100011 : OUT <= 1;  //146 / 99 = 1
    16'b10010010_01100100 : OUT <= 1;  //146 / 100 = 1
    16'b10010010_01100101 : OUT <= 1;  //146 / 101 = 1
    16'b10010010_01100110 : OUT <= 1;  //146 / 102 = 1
    16'b10010010_01100111 : OUT <= 1;  //146 / 103 = 1
    16'b10010010_01101000 : OUT <= 1;  //146 / 104 = 1
    16'b10010010_01101001 : OUT <= 1;  //146 / 105 = 1
    16'b10010010_01101010 : OUT <= 1;  //146 / 106 = 1
    16'b10010010_01101011 : OUT <= 1;  //146 / 107 = 1
    16'b10010010_01101100 : OUT <= 1;  //146 / 108 = 1
    16'b10010010_01101101 : OUT <= 1;  //146 / 109 = 1
    16'b10010010_01101110 : OUT <= 1;  //146 / 110 = 1
    16'b10010010_01101111 : OUT <= 1;  //146 / 111 = 1
    16'b10010010_01110000 : OUT <= 1;  //146 / 112 = 1
    16'b10010010_01110001 : OUT <= 1;  //146 / 113 = 1
    16'b10010010_01110010 : OUT <= 1;  //146 / 114 = 1
    16'b10010010_01110011 : OUT <= 1;  //146 / 115 = 1
    16'b10010010_01110100 : OUT <= 1;  //146 / 116 = 1
    16'b10010010_01110101 : OUT <= 1;  //146 / 117 = 1
    16'b10010010_01110110 : OUT <= 1;  //146 / 118 = 1
    16'b10010010_01110111 : OUT <= 1;  //146 / 119 = 1
    16'b10010010_01111000 : OUT <= 1;  //146 / 120 = 1
    16'b10010010_01111001 : OUT <= 1;  //146 / 121 = 1
    16'b10010010_01111010 : OUT <= 1;  //146 / 122 = 1
    16'b10010010_01111011 : OUT <= 1;  //146 / 123 = 1
    16'b10010010_01111100 : OUT <= 1;  //146 / 124 = 1
    16'b10010010_01111101 : OUT <= 1;  //146 / 125 = 1
    16'b10010010_01111110 : OUT <= 1;  //146 / 126 = 1
    16'b10010010_01111111 : OUT <= 1;  //146 / 127 = 1
    16'b10010010_10000000 : OUT <= 1;  //146 / 128 = 1
    16'b10010010_10000001 : OUT <= 1;  //146 / 129 = 1
    16'b10010010_10000010 : OUT <= 1;  //146 / 130 = 1
    16'b10010010_10000011 : OUT <= 1;  //146 / 131 = 1
    16'b10010010_10000100 : OUT <= 1;  //146 / 132 = 1
    16'b10010010_10000101 : OUT <= 1;  //146 / 133 = 1
    16'b10010010_10000110 : OUT <= 1;  //146 / 134 = 1
    16'b10010010_10000111 : OUT <= 1;  //146 / 135 = 1
    16'b10010010_10001000 : OUT <= 1;  //146 / 136 = 1
    16'b10010010_10001001 : OUT <= 1;  //146 / 137 = 1
    16'b10010010_10001010 : OUT <= 1;  //146 / 138 = 1
    16'b10010010_10001011 : OUT <= 1;  //146 / 139 = 1
    16'b10010010_10001100 : OUT <= 1;  //146 / 140 = 1
    16'b10010010_10001101 : OUT <= 1;  //146 / 141 = 1
    16'b10010010_10001110 : OUT <= 1;  //146 / 142 = 1
    16'b10010010_10001111 : OUT <= 1;  //146 / 143 = 1
    16'b10010010_10010000 : OUT <= 1;  //146 / 144 = 1
    16'b10010010_10010001 : OUT <= 1;  //146 / 145 = 1
    16'b10010010_10010010 : OUT <= 1;  //146 / 146 = 1
    16'b10010010_10010011 : OUT <= 0;  //146 / 147 = 0
    16'b10010010_10010100 : OUT <= 0;  //146 / 148 = 0
    16'b10010010_10010101 : OUT <= 0;  //146 / 149 = 0
    16'b10010010_10010110 : OUT <= 0;  //146 / 150 = 0
    16'b10010010_10010111 : OUT <= 0;  //146 / 151 = 0
    16'b10010010_10011000 : OUT <= 0;  //146 / 152 = 0
    16'b10010010_10011001 : OUT <= 0;  //146 / 153 = 0
    16'b10010010_10011010 : OUT <= 0;  //146 / 154 = 0
    16'b10010010_10011011 : OUT <= 0;  //146 / 155 = 0
    16'b10010010_10011100 : OUT <= 0;  //146 / 156 = 0
    16'b10010010_10011101 : OUT <= 0;  //146 / 157 = 0
    16'b10010010_10011110 : OUT <= 0;  //146 / 158 = 0
    16'b10010010_10011111 : OUT <= 0;  //146 / 159 = 0
    16'b10010010_10100000 : OUT <= 0;  //146 / 160 = 0
    16'b10010010_10100001 : OUT <= 0;  //146 / 161 = 0
    16'b10010010_10100010 : OUT <= 0;  //146 / 162 = 0
    16'b10010010_10100011 : OUT <= 0;  //146 / 163 = 0
    16'b10010010_10100100 : OUT <= 0;  //146 / 164 = 0
    16'b10010010_10100101 : OUT <= 0;  //146 / 165 = 0
    16'b10010010_10100110 : OUT <= 0;  //146 / 166 = 0
    16'b10010010_10100111 : OUT <= 0;  //146 / 167 = 0
    16'b10010010_10101000 : OUT <= 0;  //146 / 168 = 0
    16'b10010010_10101001 : OUT <= 0;  //146 / 169 = 0
    16'b10010010_10101010 : OUT <= 0;  //146 / 170 = 0
    16'b10010010_10101011 : OUT <= 0;  //146 / 171 = 0
    16'b10010010_10101100 : OUT <= 0;  //146 / 172 = 0
    16'b10010010_10101101 : OUT <= 0;  //146 / 173 = 0
    16'b10010010_10101110 : OUT <= 0;  //146 / 174 = 0
    16'b10010010_10101111 : OUT <= 0;  //146 / 175 = 0
    16'b10010010_10110000 : OUT <= 0;  //146 / 176 = 0
    16'b10010010_10110001 : OUT <= 0;  //146 / 177 = 0
    16'b10010010_10110010 : OUT <= 0;  //146 / 178 = 0
    16'b10010010_10110011 : OUT <= 0;  //146 / 179 = 0
    16'b10010010_10110100 : OUT <= 0;  //146 / 180 = 0
    16'b10010010_10110101 : OUT <= 0;  //146 / 181 = 0
    16'b10010010_10110110 : OUT <= 0;  //146 / 182 = 0
    16'b10010010_10110111 : OUT <= 0;  //146 / 183 = 0
    16'b10010010_10111000 : OUT <= 0;  //146 / 184 = 0
    16'b10010010_10111001 : OUT <= 0;  //146 / 185 = 0
    16'b10010010_10111010 : OUT <= 0;  //146 / 186 = 0
    16'b10010010_10111011 : OUT <= 0;  //146 / 187 = 0
    16'b10010010_10111100 : OUT <= 0;  //146 / 188 = 0
    16'b10010010_10111101 : OUT <= 0;  //146 / 189 = 0
    16'b10010010_10111110 : OUT <= 0;  //146 / 190 = 0
    16'b10010010_10111111 : OUT <= 0;  //146 / 191 = 0
    16'b10010010_11000000 : OUT <= 0;  //146 / 192 = 0
    16'b10010010_11000001 : OUT <= 0;  //146 / 193 = 0
    16'b10010010_11000010 : OUT <= 0;  //146 / 194 = 0
    16'b10010010_11000011 : OUT <= 0;  //146 / 195 = 0
    16'b10010010_11000100 : OUT <= 0;  //146 / 196 = 0
    16'b10010010_11000101 : OUT <= 0;  //146 / 197 = 0
    16'b10010010_11000110 : OUT <= 0;  //146 / 198 = 0
    16'b10010010_11000111 : OUT <= 0;  //146 / 199 = 0
    16'b10010010_11001000 : OUT <= 0;  //146 / 200 = 0
    16'b10010010_11001001 : OUT <= 0;  //146 / 201 = 0
    16'b10010010_11001010 : OUT <= 0;  //146 / 202 = 0
    16'b10010010_11001011 : OUT <= 0;  //146 / 203 = 0
    16'b10010010_11001100 : OUT <= 0;  //146 / 204 = 0
    16'b10010010_11001101 : OUT <= 0;  //146 / 205 = 0
    16'b10010010_11001110 : OUT <= 0;  //146 / 206 = 0
    16'b10010010_11001111 : OUT <= 0;  //146 / 207 = 0
    16'b10010010_11010000 : OUT <= 0;  //146 / 208 = 0
    16'b10010010_11010001 : OUT <= 0;  //146 / 209 = 0
    16'b10010010_11010010 : OUT <= 0;  //146 / 210 = 0
    16'b10010010_11010011 : OUT <= 0;  //146 / 211 = 0
    16'b10010010_11010100 : OUT <= 0;  //146 / 212 = 0
    16'b10010010_11010101 : OUT <= 0;  //146 / 213 = 0
    16'b10010010_11010110 : OUT <= 0;  //146 / 214 = 0
    16'b10010010_11010111 : OUT <= 0;  //146 / 215 = 0
    16'b10010010_11011000 : OUT <= 0;  //146 / 216 = 0
    16'b10010010_11011001 : OUT <= 0;  //146 / 217 = 0
    16'b10010010_11011010 : OUT <= 0;  //146 / 218 = 0
    16'b10010010_11011011 : OUT <= 0;  //146 / 219 = 0
    16'b10010010_11011100 : OUT <= 0;  //146 / 220 = 0
    16'b10010010_11011101 : OUT <= 0;  //146 / 221 = 0
    16'b10010010_11011110 : OUT <= 0;  //146 / 222 = 0
    16'b10010010_11011111 : OUT <= 0;  //146 / 223 = 0
    16'b10010010_11100000 : OUT <= 0;  //146 / 224 = 0
    16'b10010010_11100001 : OUT <= 0;  //146 / 225 = 0
    16'b10010010_11100010 : OUT <= 0;  //146 / 226 = 0
    16'b10010010_11100011 : OUT <= 0;  //146 / 227 = 0
    16'b10010010_11100100 : OUT <= 0;  //146 / 228 = 0
    16'b10010010_11100101 : OUT <= 0;  //146 / 229 = 0
    16'b10010010_11100110 : OUT <= 0;  //146 / 230 = 0
    16'b10010010_11100111 : OUT <= 0;  //146 / 231 = 0
    16'b10010010_11101000 : OUT <= 0;  //146 / 232 = 0
    16'b10010010_11101001 : OUT <= 0;  //146 / 233 = 0
    16'b10010010_11101010 : OUT <= 0;  //146 / 234 = 0
    16'b10010010_11101011 : OUT <= 0;  //146 / 235 = 0
    16'b10010010_11101100 : OUT <= 0;  //146 / 236 = 0
    16'b10010010_11101101 : OUT <= 0;  //146 / 237 = 0
    16'b10010010_11101110 : OUT <= 0;  //146 / 238 = 0
    16'b10010010_11101111 : OUT <= 0;  //146 / 239 = 0
    16'b10010010_11110000 : OUT <= 0;  //146 / 240 = 0
    16'b10010010_11110001 : OUT <= 0;  //146 / 241 = 0
    16'b10010010_11110010 : OUT <= 0;  //146 / 242 = 0
    16'b10010010_11110011 : OUT <= 0;  //146 / 243 = 0
    16'b10010010_11110100 : OUT <= 0;  //146 / 244 = 0
    16'b10010010_11110101 : OUT <= 0;  //146 / 245 = 0
    16'b10010010_11110110 : OUT <= 0;  //146 / 246 = 0
    16'b10010010_11110111 : OUT <= 0;  //146 / 247 = 0
    16'b10010010_11111000 : OUT <= 0;  //146 / 248 = 0
    16'b10010010_11111001 : OUT <= 0;  //146 / 249 = 0
    16'b10010010_11111010 : OUT <= 0;  //146 / 250 = 0
    16'b10010010_11111011 : OUT <= 0;  //146 / 251 = 0
    16'b10010010_11111100 : OUT <= 0;  //146 / 252 = 0
    16'b10010010_11111101 : OUT <= 0;  //146 / 253 = 0
    16'b10010010_11111110 : OUT <= 0;  //146 / 254 = 0
    16'b10010010_11111111 : OUT <= 0;  //146 / 255 = 0
    16'b10010011_00000000 : OUT <= 0;  //147 / 0 = 0
    16'b10010011_00000001 : OUT <= 147;  //147 / 1 = 147
    16'b10010011_00000010 : OUT <= 73;  //147 / 2 = 73
    16'b10010011_00000011 : OUT <= 49;  //147 / 3 = 49
    16'b10010011_00000100 : OUT <= 36;  //147 / 4 = 36
    16'b10010011_00000101 : OUT <= 29;  //147 / 5 = 29
    16'b10010011_00000110 : OUT <= 24;  //147 / 6 = 24
    16'b10010011_00000111 : OUT <= 21;  //147 / 7 = 21
    16'b10010011_00001000 : OUT <= 18;  //147 / 8 = 18
    16'b10010011_00001001 : OUT <= 16;  //147 / 9 = 16
    16'b10010011_00001010 : OUT <= 14;  //147 / 10 = 14
    16'b10010011_00001011 : OUT <= 13;  //147 / 11 = 13
    16'b10010011_00001100 : OUT <= 12;  //147 / 12 = 12
    16'b10010011_00001101 : OUT <= 11;  //147 / 13 = 11
    16'b10010011_00001110 : OUT <= 10;  //147 / 14 = 10
    16'b10010011_00001111 : OUT <= 9;  //147 / 15 = 9
    16'b10010011_00010000 : OUT <= 9;  //147 / 16 = 9
    16'b10010011_00010001 : OUT <= 8;  //147 / 17 = 8
    16'b10010011_00010010 : OUT <= 8;  //147 / 18 = 8
    16'b10010011_00010011 : OUT <= 7;  //147 / 19 = 7
    16'b10010011_00010100 : OUT <= 7;  //147 / 20 = 7
    16'b10010011_00010101 : OUT <= 7;  //147 / 21 = 7
    16'b10010011_00010110 : OUT <= 6;  //147 / 22 = 6
    16'b10010011_00010111 : OUT <= 6;  //147 / 23 = 6
    16'b10010011_00011000 : OUT <= 6;  //147 / 24 = 6
    16'b10010011_00011001 : OUT <= 5;  //147 / 25 = 5
    16'b10010011_00011010 : OUT <= 5;  //147 / 26 = 5
    16'b10010011_00011011 : OUT <= 5;  //147 / 27 = 5
    16'b10010011_00011100 : OUT <= 5;  //147 / 28 = 5
    16'b10010011_00011101 : OUT <= 5;  //147 / 29 = 5
    16'b10010011_00011110 : OUT <= 4;  //147 / 30 = 4
    16'b10010011_00011111 : OUT <= 4;  //147 / 31 = 4
    16'b10010011_00100000 : OUT <= 4;  //147 / 32 = 4
    16'b10010011_00100001 : OUT <= 4;  //147 / 33 = 4
    16'b10010011_00100010 : OUT <= 4;  //147 / 34 = 4
    16'b10010011_00100011 : OUT <= 4;  //147 / 35 = 4
    16'b10010011_00100100 : OUT <= 4;  //147 / 36 = 4
    16'b10010011_00100101 : OUT <= 3;  //147 / 37 = 3
    16'b10010011_00100110 : OUT <= 3;  //147 / 38 = 3
    16'b10010011_00100111 : OUT <= 3;  //147 / 39 = 3
    16'b10010011_00101000 : OUT <= 3;  //147 / 40 = 3
    16'b10010011_00101001 : OUT <= 3;  //147 / 41 = 3
    16'b10010011_00101010 : OUT <= 3;  //147 / 42 = 3
    16'b10010011_00101011 : OUT <= 3;  //147 / 43 = 3
    16'b10010011_00101100 : OUT <= 3;  //147 / 44 = 3
    16'b10010011_00101101 : OUT <= 3;  //147 / 45 = 3
    16'b10010011_00101110 : OUT <= 3;  //147 / 46 = 3
    16'b10010011_00101111 : OUT <= 3;  //147 / 47 = 3
    16'b10010011_00110000 : OUT <= 3;  //147 / 48 = 3
    16'b10010011_00110001 : OUT <= 3;  //147 / 49 = 3
    16'b10010011_00110010 : OUT <= 2;  //147 / 50 = 2
    16'b10010011_00110011 : OUT <= 2;  //147 / 51 = 2
    16'b10010011_00110100 : OUT <= 2;  //147 / 52 = 2
    16'b10010011_00110101 : OUT <= 2;  //147 / 53 = 2
    16'b10010011_00110110 : OUT <= 2;  //147 / 54 = 2
    16'b10010011_00110111 : OUT <= 2;  //147 / 55 = 2
    16'b10010011_00111000 : OUT <= 2;  //147 / 56 = 2
    16'b10010011_00111001 : OUT <= 2;  //147 / 57 = 2
    16'b10010011_00111010 : OUT <= 2;  //147 / 58 = 2
    16'b10010011_00111011 : OUT <= 2;  //147 / 59 = 2
    16'b10010011_00111100 : OUT <= 2;  //147 / 60 = 2
    16'b10010011_00111101 : OUT <= 2;  //147 / 61 = 2
    16'b10010011_00111110 : OUT <= 2;  //147 / 62 = 2
    16'b10010011_00111111 : OUT <= 2;  //147 / 63 = 2
    16'b10010011_01000000 : OUT <= 2;  //147 / 64 = 2
    16'b10010011_01000001 : OUT <= 2;  //147 / 65 = 2
    16'b10010011_01000010 : OUT <= 2;  //147 / 66 = 2
    16'b10010011_01000011 : OUT <= 2;  //147 / 67 = 2
    16'b10010011_01000100 : OUT <= 2;  //147 / 68 = 2
    16'b10010011_01000101 : OUT <= 2;  //147 / 69 = 2
    16'b10010011_01000110 : OUT <= 2;  //147 / 70 = 2
    16'b10010011_01000111 : OUT <= 2;  //147 / 71 = 2
    16'b10010011_01001000 : OUT <= 2;  //147 / 72 = 2
    16'b10010011_01001001 : OUT <= 2;  //147 / 73 = 2
    16'b10010011_01001010 : OUT <= 1;  //147 / 74 = 1
    16'b10010011_01001011 : OUT <= 1;  //147 / 75 = 1
    16'b10010011_01001100 : OUT <= 1;  //147 / 76 = 1
    16'b10010011_01001101 : OUT <= 1;  //147 / 77 = 1
    16'b10010011_01001110 : OUT <= 1;  //147 / 78 = 1
    16'b10010011_01001111 : OUT <= 1;  //147 / 79 = 1
    16'b10010011_01010000 : OUT <= 1;  //147 / 80 = 1
    16'b10010011_01010001 : OUT <= 1;  //147 / 81 = 1
    16'b10010011_01010010 : OUT <= 1;  //147 / 82 = 1
    16'b10010011_01010011 : OUT <= 1;  //147 / 83 = 1
    16'b10010011_01010100 : OUT <= 1;  //147 / 84 = 1
    16'b10010011_01010101 : OUT <= 1;  //147 / 85 = 1
    16'b10010011_01010110 : OUT <= 1;  //147 / 86 = 1
    16'b10010011_01010111 : OUT <= 1;  //147 / 87 = 1
    16'b10010011_01011000 : OUT <= 1;  //147 / 88 = 1
    16'b10010011_01011001 : OUT <= 1;  //147 / 89 = 1
    16'b10010011_01011010 : OUT <= 1;  //147 / 90 = 1
    16'b10010011_01011011 : OUT <= 1;  //147 / 91 = 1
    16'b10010011_01011100 : OUT <= 1;  //147 / 92 = 1
    16'b10010011_01011101 : OUT <= 1;  //147 / 93 = 1
    16'b10010011_01011110 : OUT <= 1;  //147 / 94 = 1
    16'b10010011_01011111 : OUT <= 1;  //147 / 95 = 1
    16'b10010011_01100000 : OUT <= 1;  //147 / 96 = 1
    16'b10010011_01100001 : OUT <= 1;  //147 / 97 = 1
    16'b10010011_01100010 : OUT <= 1;  //147 / 98 = 1
    16'b10010011_01100011 : OUT <= 1;  //147 / 99 = 1
    16'b10010011_01100100 : OUT <= 1;  //147 / 100 = 1
    16'b10010011_01100101 : OUT <= 1;  //147 / 101 = 1
    16'b10010011_01100110 : OUT <= 1;  //147 / 102 = 1
    16'b10010011_01100111 : OUT <= 1;  //147 / 103 = 1
    16'b10010011_01101000 : OUT <= 1;  //147 / 104 = 1
    16'b10010011_01101001 : OUT <= 1;  //147 / 105 = 1
    16'b10010011_01101010 : OUT <= 1;  //147 / 106 = 1
    16'b10010011_01101011 : OUT <= 1;  //147 / 107 = 1
    16'b10010011_01101100 : OUT <= 1;  //147 / 108 = 1
    16'b10010011_01101101 : OUT <= 1;  //147 / 109 = 1
    16'b10010011_01101110 : OUT <= 1;  //147 / 110 = 1
    16'b10010011_01101111 : OUT <= 1;  //147 / 111 = 1
    16'b10010011_01110000 : OUT <= 1;  //147 / 112 = 1
    16'b10010011_01110001 : OUT <= 1;  //147 / 113 = 1
    16'b10010011_01110010 : OUT <= 1;  //147 / 114 = 1
    16'b10010011_01110011 : OUT <= 1;  //147 / 115 = 1
    16'b10010011_01110100 : OUT <= 1;  //147 / 116 = 1
    16'b10010011_01110101 : OUT <= 1;  //147 / 117 = 1
    16'b10010011_01110110 : OUT <= 1;  //147 / 118 = 1
    16'b10010011_01110111 : OUT <= 1;  //147 / 119 = 1
    16'b10010011_01111000 : OUT <= 1;  //147 / 120 = 1
    16'b10010011_01111001 : OUT <= 1;  //147 / 121 = 1
    16'b10010011_01111010 : OUT <= 1;  //147 / 122 = 1
    16'b10010011_01111011 : OUT <= 1;  //147 / 123 = 1
    16'b10010011_01111100 : OUT <= 1;  //147 / 124 = 1
    16'b10010011_01111101 : OUT <= 1;  //147 / 125 = 1
    16'b10010011_01111110 : OUT <= 1;  //147 / 126 = 1
    16'b10010011_01111111 : OUT <= 1;  //147 / 127 = 1
    16'b10010011_10000000 : OUT <= 1;  //147 / 128 = 1
    16'b10010011_10000001 : OUT <= 1;  //147 / 129 = 1
    16'b10010011_10000010 : OUT <= 1;  //147 / 130 = 1
    16'b10010011_10000011 : OUT <= 1;  //147 / 131 = 1
    16'b10010011_10000100 : OUT <= 1;  //147 / 132 = 1
    16'b10010011_10000101 : OUT <= 1;  //147 / 133 = 1
    16'b10010011_10000110 : OUT <= 1;  //147 / 134 = 1
    16'b10010011_10000111 : OUT <= 1;  //147 / 135 = 1
    16'b10010011_10001000 : OUT <= 1;  //147 / 136 = 1
    16'b10010011_10001001 : OUT <= 1;  //147 / 137 = 1
    16'b10010011_10001010 : OUT <= 1;  //147 / 138 = 1
    16'b10010011_10001011 : OUT <= 1;  //147 / 139 = 1
    16'b10010011_10001100 : OUT <= 1;  //147 / 140 = 1
    16'b10010011_10001101 : OUT <= 1;  //147 / 141 = 1
    16'b10010011_10001110 : OUT <= 1;  //147 / 142 = 1
    16'b10010011_10001111 : OUT <= 1;  //147 / 143 = 1
    16'b10010011_10010000 : OUT <= 1;  //147 / 144 = 1
    16'b10010011_10010001 : OUT <= 1;  //147 / 145 = 1
    16'b10010011_10010010 : OUT <= 1;  //147 / 146 = 1
    16'b10010011_10010011 : OUT <= 1;  //147 / 147 = 1
    16'b10010011_10010100 : OUT <= 0;  //147 / 148 = 0
    16'b10010011_10010101 : OUT <= 0;  //147 / 149 = 0
    16'b10010011_10010110 : OUT <= 0;  //147 / 150 = 0
    16'b10010011_10010111 : OUT <= 0;  //147 / 151 = 0
    16'b10010011_10011000 : OUT <= 0;  //147 / 152 = 0
    16'b10010011_10011001 : OUT <= 0;  //147 / 153 = 0
    16'b10010011_10011010 : OUT <= 0;  //147 / 154 = 0
    16'b10010011_10011011 : OUT <= 0;  //147 / 155 = 0
    16'b10010011_10011100 : OUT <= 0;  //147 / 156 = 0
    16'b10010011_10011101 : OUT <= 0;  //147 / 157 = 0
    16'b10010011_10011110 : OUT <= 0;  //147 / 158 = 0
    16'b10010011_10011111 : OUT <= 0;  //147 / 159 = 0
    16'b10010011_10100000 : OUT <= 0;  //147 / 160 = 0
    16'b10010011_10100001 : OUT <= 0;  //147 / 161 = 0
    16'b10010011_10100010 : OUT <= 0;  //147 / 162 = 0
    16'b10010011_10100011 : OUT <= 0;  //147 / 163 = 0
    16'b10010011_10100100 : OUT <= 0;  //147 / 164 = 0
    16'b10010011_10100101 : OUT <= 0;  //147 / 165 = 0
    16'b10010011_10100110 : OUT <= 0;  //147 / 166 = 0
    16'b10010011_10100111 : OUT <= 0;  //147 / 167 = 0
    16'b10010011_10101000 : OUT <= 0;  //147 / 168 = 0
    16'b10010011_10101001 : OUT <= 0;  //147 / 169 = 0
    16'b10010011_10101010 : OUT <= 0;  //147 / 170 = 0
    16'b10010011_10101011 : OUT <= 0;  //147 / 171 = 0
    16'b10010011_10101100 : OUT <= 0;  //147 / 172 = 0
    16'b10010011_10101101 : OUT <= 0;  //147 / 173 = 0
    16'b10010011_10101110 : OUT <= 0;  //147 / 174 = 0
    16'b10010011_10101111 : OUT <= 0;  //147 / 175 = 0
    16'b10010011_10110000 : OUT <= 0;  //147 / 176 = 0
    16'b10010011_10110001 : OUT <= 0;  //147 / 177 = 0
    16'b10010011_10110010 : OUT <= 0;  //147 / 178 = 0
    16'b10010011_10110011 : OUT <= 0;  //147 / 179 = 0
    16'b10010011_10110100 : OUT <= 0;  //147 / 180 = 0
    16'b10010011_10110101 : OUT <= 0;  //147 / 181 = 0
    16'b10010011_10110110 : OUT <= 0;  //147 / 182 = 0
    16'b10010011_10110111 : OUT <= 0;  //147 / 183 = 0
    16'b10010011_10111000 : OUT <= 0;  //147 / 184 = 0
    16'b10010011_10111001 : OUT <= 0;  //147 / 185 = 0
    16'b10010011_10111010 : OUT <= 0;  //147 / 186 = 0
    16'b10010011_10111011 : OUT <= 0;  //147 / 187 = 0
    16'b10010011_10111100 : OUT <= 0;  //147 / 188 = 0
    16'b10010011_10111101 : OUT <= 0;  //147 / 189 = 0
    16'b10010011_10111110 : OUT <= 0;  //147 / 190 = 0
    16'b10010011_10111111 : OUT <= 0;  //147 / 191 = 0
    16'b10010011_11000000 : OUT <= 0;  //147 / 192 = 0
    16'b10010011_11000001 : OUT <= 0;  //147 / 193 = 0
    16'b10010011_11000010 : OUT <= 0;  //147 / 194 = 0
    16'b10010011_11000011 : OUT <= 0;  //147 / 195 = 0
    16'b10010011_11000100 : OUT <= 0;  //147 / 196 = 0
    16'b10010011_11000101 : OUT <= 0;  //147 / 197 = 0
    16'b10010011_11000110 : OUT <= 0;  //147 / 198 = 0
    16'b10010011_11000111 : OUT <= 0;  //147 / 199 = 0
    16'b10010011_11001000 : OUT <= 0;  //147 / 200 = 0
    16'b10010011_11001001 : OUT <= 0;  //147 / 201 = 0
    16'b10010011_11001010 : OUT <= 0;  //147 / 202 = 0
    16'b10010011_11001011 : OUT <= 0;  //147 / 203 = 0
    16'b10010011_11001100 : OUT <= 0;  //147 / 204 = 0
    16'b10010011_11001101 : OUT <= 0;  //147 / 205 = 0
    16'b10010011_11001110 : OUT <= 0;  //147 / 206 = 0
    16'b10010011_11001111 : OUT <= 0;  //147 / 207 = 0
    16'b10010011_11010000 : OUT <= 0;  //147 / 208 = 0
    16'b10010011_11010001 : OUT <= 0;  //147 / 209 = 0
    16'b10010011_11010010 : OUT <= 0;  //147 / 210 = 0
    16'b10010011_11010011 : OUT <= 0;  //147 / 211 = 0
    16'b10010011_11010100 : OUT <= 0;  //147 / 212 = 0
    16'b10010011_11010101 : OUT <= 0;  //147 / 213 = 0
    16'b10010011_11010110 : OUT <= 0;  //147 / 214 = 0
    16'b10010011_11010111 : OUT <= 0;  //147 / 215 = 0
    16'b10010011_11011000 : OUT <= 0;  //147 / 216 = 0
    16'b10010011_11011001 : OUT <= 0;  //147 / 217 = 0
    16'b10010011_11011010 : OUT <= 0;  //147 / 218 = 0
    16'b10010011_11011011 : OUT <= 0;  //147 / 219 = 0
    16'b10010011_11011100 : OUT <= 0;  //147 / 220 = 0
    16'b10010011_11011101 : OUT <= 0;  //147 / 221 = 0
    16'b10010011_11011110 : OUT <= 0;  //147 / 222 = 0
    16'b10010011_11011111 : OUT <= 0;  //147 / 223 = 0
    16'b10010011_11100000 : OUT <= 0;  //147 / 224 = 0
    16'b10010011_11100001 : OUT <= 0;  //147 / 225 = 0
    16'b10010011_11100010 : OUT <= 0;  //147 / 226 = 0
    16'b10010011_11100011 : OUT <= 0;  //147 / 227 = 0
    16'b10010011_11100100 : OUT <= 0;  //147 / 228 = 0
    16'b10010011_11100101 : OUT <= 0;  //147 / 229 = 0
    16'b10010011_11100110 : OUT <= 0;  //147 / 230 = 0
    16'b10010011_11100111 : OUT <= 0;  //147 / 231 = 0
    16'b10010011_11101000 : OUT <= 0;  //147 / 232 = 0
    16'b10010011_11101001 : OUT <= 0;  //147 / 233 = 0
    16'b10010011_11101010 : OUT <= 0;  //147 / 234 = 0
    16'b10010011_11101011 : OUT <= 0;  //147 / 235 = 0
    16'b10010011_11101100 : OUT <= 0;  //147 / 236 = 0
    16'b10010011_11101101 : OUT <= 0;  //147 / 237 = 0
    16'b10010011_11101110 : OUT <= 0;  //147 / 238 = 0
    16'b10010011_11101111 : OUT <= 0;  //147 / 239 = 0
    16'b10010011_11110000 : OUT <= 0;  //147 / 240 = 0
    16'b10010011_11110001 : OUT <= 0;  //147 / 241 = 0
    16'b10010011_11110010 : OUT <= 0;  //147 / 242 = 0
    16'b10010011_11110011 : OUT <= 0;  //147 / 243 = 0
    16'b10010011_11110100 : OUT <= 0;  //147 / 244 = 0
    16'b10010011_11110101 : OUT <= 0;  //147 / 245 = 0
    16'b10010011_11110110 : OUT <= 0;  //147 / 246 = 0
    16'b10010011_11110111 : OUT <= 0;  //147 / 247 = 0
    16'b10010011_11111000 : OUT <= 0;  //147 / 248 = 0
    16'b10010011_11111001 : OUT <= 0;  //147 / 249 = 0
    16'b10010011_11111010 : OUT <= 0;  //147 / 250 = 0
    16'b10010011_11111011 : OUT <= 0;  //147 / 251 = 0
    16'b10010011_11111100 : OUT <= 0;  //147 / 252 = 0
    16'b10010011_11111101 : OUT <= 0;  //147 / 253 = 0
    16'b10010011_11111110 : OUT <= 0;  //147 / 254 = 0
    16'b10010011_11111111 : OUT <= 0;  //147 / 255 = 0
    16'b10010100_00000000 : OUT <= 0;  //148 / 0 = 0
    16'b10010100_00000001 : OUT <= 148;  //148 / 1 = 148
    16'b10010100_00000010 : OUT <= 74;  //148 / 2 = 74
    16'b10010100_00000011 : OUT <= 49;  //148 / 3 = 49
    16'b10010100_00000100 : OUT <= 37;  //148 / 4 = 37
    16'b10010100_00000101 : OUT <= 29;  //148 / 5 = 29
    16'b10010100_00000110 : OUT <= 24;  //148 / 6 = 24
    16'b10010100_00000111 : OUT <= 21;  //148 / 7 = 21
    16'b10010100_00001000 : OUT <= 18;  //148 / 8 = 18
    16'b10010100_00001001 : OUT <= 16;  //148 / 9 = 16
    16'b10010100_00001010 : OUT <= 14;  //148 / 10 = 14
    16'b10010100_00001011 : OUT <= 13;  //148 / 11 = 13
    16'b10010100_00001100 : OUT <= 12;  //148 / 12 = 12
    16'b10010100_00001101 : OUT <= 11;  //148 / 13 = 11
    16'b10010100_00001110 : OUT <= 10;  //148 / 14 = 10
    16'b10010100_00001111 : OUT <= 9;  //148 / 15 = 9
    16'b10010100_00010000 : OUT <= 9;  //148 / 16 = 9
    16'b10010100_00010001 : OUT <= 8;  //148 / 17 = 8
    16'b10010100_00010010 : OUT <= 8;  //148 / 18 = 8
    16'b10010100_00010011 : OUT <= 7;  //148 / 19 = 7
    16'b10010100_00010100 : OUT <= 7;  //148 / 20 = 7
    16'b10010100_00010101 : OUT <= 7;  //148 / 21 = 7
    16'b10010100_00010110 : OUT <= 6;  //148 / 22 = 6
    16'b10010100_00010111 : OUT <= 6;  //148 / 23 = 6
    16'b10010100_00011000 : OUT <= 6;  //148 / 24 = 6
    16'b10010100_00011001 : OUT <= 5;  //148 / 25 = 5
    16'b10010100_00011010 : OUT <= 5;  //148 / 26 = 5
    16'b10010100_00011011 : OUT <= 5;  //148 / 27 = 5
    16'b10010100_00011100 : OUT <= 5;  //148 / 28 = 5
    16'b10010100_00011101 : OUT <= 5;  //148 / 29 = 5
    16'b10010100_00011110 : OUT <= 4;  //148 / 30 = 4
    16'b10010100_00011111 : OUT <= 4;  //148 / 31 = 4
    16'b10010100_00100000 : OUT <= 4;  //148 / 32 = 4
    16'b10010100_00100001 : OUT <= 4;  //148 / 33 = 4
    16'b10010100_00100010 : OUT <= 4;  //148 / 34 = 4
    16'b10010100_00100011 : OUT <= 4;  //148 / 35 = 4
    16'b10010100_00100100 : OUT <= 4;  //148 / 36 = 4
    16'b10010100_00100101 : OUT <= 4;  //148 / 37 = 4
    16'b10010100_00100110 : OUT <= 3;  //148 / 38 = 3
    16'b10010100_00100111 : OUT <= 3;  //148 / 39 = 3
    16'b10010100_00101000 : OUT <= 3;  //148 / 40 = 3
    16'b10010100_00101001 : OUT <= 3;  //148 / 41 = 3
    16'b10010100_00101010 : OUT <= 3;  //148 / 42 = 3
    16'b10010100_00101011 : OUT <= 3;  //148 / 43 = 3
    16'b10010100_00101100 : OUT <= 3;  //148 / 44 = 3
    16'b10010100_00101101 : OUT <= 3;  //148 / 45 = 3
    16'b10010100_00101110 : OUT <= 3;  //148 / 46 = 3
    16'b10010100_00101111 : OUT <= 3;  //148 / 47 = 3
    16'b10010100_00110000 : OUT <= 3;  //148 / 48 = 3
    16'b10010100_00110001 : OUT <= 3;  //148 / 49 = 3
    16'b10010100_00110010 : OUT <= 2;  //148 / 50 = 2
    16'b10010100_00110011 : OUT <= 2;  //148 / 51 = 2
    16'b10010100_00110100 : OUT <= 2;  //148 / 52 = 2
    16'b10010100_00110101 : OUT <= 2;  //148 / 53 = 2
    16'b10010100_00110110 : OUT <= 2;  //148 / 54 = 2
    16'b10010100_00110111 : OUT <= 2;  //148 / 55 = 2
    16'b10010100_00111000 : OUT <= 2;  //148 / 56 = 2
    16'b10010100_00111001 : OUT <= 2;  //148 / 57 = 2
    16'b10010100_00111010 : OUT <= 2;  //148 / 58 = 2
    16'b10010100_00111011 : OUT <= 2;  //148 / 59 = 2
    16'b10010100_00111100 : OUT <= 2;  //148 / 60 = 2
    16'b10010100_00111101 : OUT <= 2;  //148 / 61 = 2
    16'b10010100_00111110 : OUT <= 2;  //148 / 62 = 2
    16'b10010100_00111111 : OUT <= 2;  //148 / 63 = 2
    16'b10010100_01000000 : OUT <= 2;  //148 / 64 = 2
    16'b10010100_01000001 : OUT <= 2;  //148 / 65 = 2
    16'b10010100_01000010 : OUT <= 2;  //148 / 66 = 2
    16'b10010100_01000011 : OUT <= 2;  //148 / 67 = 2
    16'b10010100_01000100 : OUT <= 2;  //148 / 68 = 2
    16'b10010100_01000101 : OUT <= 2;  //148 / 69 = 2
    16'b10010100_01000110 : OUT <= 2;  //148 / 70 = 2
    16'b10010100_01000111 : OUT <= 2;  //148 / 71 = 2
    16'b10010100_01001000 : OUT <= 2;  //148 / 72 = 2
    16'b10010100_01001001 : OUT <= 2;  //148 / 73 = 2
    16'b10010100_01001010 : OUT <= 2;  //148 / 74 = 2
    16'b10010100_01001011 : OUT <= 1;  //148 / 75 = 1
    16'b10010100_01001100 : OUT <= 1;  //148 / 76 = 1
    16'b10010100_01001101 : OUT <= 1;  //148 / 77 = 1
    16'b10010100_01001110 : OUT <= 1;  //148 / 78 = 1
    16'b10010100_01001111 : OUT <= 1;  //148 / 79 = 1
    16'b10010100_01010000 : OUT <= 1;  //148 / 80 = 1
    16'b10010100_01010001 : OUT <= 1;  //148 / 81 = 1
    16'b10010100_01010010 : OUT <= 1;  //148 / 82 = 1
    16'b10010100_01010011 : OUT <= 1;  //148 / 83 = 1
    16'b10010100_01010100 : OUT <= 1;  //148 / 84 = 1
    16'b10010100_01010101 : OUT <= 1;  //148 / 85 = 1
    16'b10010100_01010110 : OUT <= 1;  //148 / 86 = 1
    16'b10010100_01010111 : OUT <= 1;  //148 / 87 = 1
    16'b10010100_01011000 : OUT <= 1;  //148 / 88 = 1
    16'b10010100_01011001 : OUT <= 1;  //148 / 89 = 1
    16'b10010100_01011010 : OUT <= 1;  //148 / 90 = 1
    16'b10010100_01011011 : OUT <= 1;  //148 / 91 = 1
    16'b10010100_01011100 : OUT <= 1;  //148 / 92 = 1
    16'b10010100_01011101 : OUT <= 1;  //148 / 93 = 1
    16'b10010100_01011110 : OUT <= 1;  //148 / 94 = 1
    16'b10010100_01011111 : OUT <= 1;  //148 / 95 = 1
    16'b10010100_01100000 : OUT <= 1;  //148 / 96 = 1
    16'b10010100_01100001 : OUT <= 1;  //148 / 97 = 1
    16'b10010100_01100010 : OUT <= 1;  //148 / 98 = 1
    16'b10010100_01100011 : OUT <= 1;  //148 / 99 = 1
    16'b10010100_01100100 : OUT <= 1;  //148 / 100 = 1
    16'b10010100_01100101 : OUT <= 1;  //148 / 101 = 1
    16'b10010100_01100110 : OUT <= 1;  //148 / 102 = 1
    16'b10010100_01100111 : OUT <= 1;  //148 / 103 = 1
    16'b10010100_01101000 : OUT <= 1;  //148 / 104 = 1
    16'b10010100_01101001 : OUT <= 1;  //148 / 105 = 1
    16'b10010100_01101010 : OUT <= 1;  //148 / 106 = 1
    16'b10010100_01101011 : OUT <= 1;  //148 / 107 = 1
    16'b10010100_01101100 : OUT <= 1;  //148 / 108 = 1
    16'b10010100_01101101 : OUT <= 1;  //148 / 109 = 1
    16'b10010100_01101110 : OUT <= 1;  //148 / 110 = 1
    16'b10010100_01101111 : OUT <= 1;  //148 / 111 = 1
    16'b10010100_01110000 : OUT <= 1;  //148 / 112 = 1
    16'b10010100_01110001 : OUT <= 1;  //148 / 113 = 1
    16'b10010100_01110010 : OUT <= 1;  //148 / 114 = 1
    16'b10010100_01110011 : OUT <= 1;  //148 / 115 = 1
    16'b10010100_01110100 : OUT <= 1;  //148 / 116 = 1
    16'b10010100_01110101 : OUT <= 1;  //148 / 117 = 1
    16'b10010100_01110110 : OUT <= 1;  //148 / 118 = 1
    16'b10010100_01110111 : OUT <= 1;  //148 / 119 = 1
    16'b10010100_01111000 : OUT <= 1;  //148 / 120 = 1
    16'b10010100_01111001 : OUT <= 1;  //148 / 121 = 1
    16'b10010100_01111010 : OUT <= 1;  //148 / 122 = 1
    16'b10010100_01111011 : OUT <= 1;  //148 / 123 = 1
    16'b10010100_01111100 : OUT <= 1;  //148 / 124 = 1
    16'b10010100_01111101 : OUT <= 1;  //148 / 125 = 1
    16'b10010100_01111110 : OUT <= 1;  //148 / 126 = 1
    16'b10010100_01111111 : OUT <= 1;  //148 / 127 = 1
    16'b10010100_10000000 : OUT <= 1;  //148 / 128 = 1
    16'b10010100_10000001 : OUT <= 1;  //148 / 129 = 1
    16'b10010100_10000010 : OUT <= 1;  //148 / 130 = 1
    16'b10010100_10000011 : OUT <= 1;  //148 / 131 = 1
    16'b10010100_10000100 : OUT <= 1;  //148 / 132 = 1
    16'b10010100_10000101 : OUT <= 1;  //148 / 133 = 1
    16'b10010100_10000110 : OUT <= 1;  //148 / 134 = 1
    16'b10010100_10000111 : OUT <= 1;  //148 / 135 = 1
    16'b10010100_10001000 : OUT <= 1;  //148 / 136 = 1
    16'b10010100_10001001 : OUT <= 1;  //148 / 137 = 1
    16'b10010100_10001010 : OUT <= 1;  //148 / 138 = 1
    16'b10010100_10001011 : OUT <= 1;  //148 / 139 = 1
    16'b10010100_10001100 : OUT <= 1;  //148 / 140 = 1
    16'b10010100_10001101 : OUT <= 1;  //148 / 141 = 1
    16'b10010100_10001110 : OUT <= 1;  //148 / 142 = 1
    16'b10010100_10001111 : OUT <= 1;  //148 / 143 = 1
    16'b10010100_10010000 : OUT <= 1;  //148 / 144 = 1
    16'b10010100_10010001 : OUT <= 1;  //148 / 145 = 1
    16'b10010100_10010010 : OUT <= 1;  //148 / 146 = 1
    16'b10010100_10010011 : OUT <= 1;  //148 / 147 = 1
    16'b10010100_10010100 : OUT <= 1;  //148 / 148 = 1
    16'b10010100_10010101 : OUT <= 0;  //148 / 149 = 0
    16'b10010100_10010110 : OUT <= 0;  //148 / 150 = 0
    16'b10010100_10010111 : OUT <= 0;  //148 / 151 = 0
    16'b10010100_10011000 : OUT <= 0;  //148 / 152 = 0
    16'b10010100_10011001 : OUT <= 0;  //148 / 153 = 0
    16'b10010100_10011010 : OUT <= 0;  //148 / 154 = 0
    16'b10010100_10011011 : OUT <= 0;  //148 / 155 = 0
    16'b10010100_10011100 : OUT <= 0;  //148 / 156 = 0
    16'b10010100_10011101 : OUT <= 0;  //148 / 157 = 0
    16'b10010100_10011110 : OUT <= 0;  //148 / 158 = 0
    16'b10010100_10011111 : OUT <= 0;  //148 / 159 = 0
    16'b10010100_10100000 : OUT <= 0;  //148 / 160 = 0
    16'b10010100_10100001 : OUT <= 0;  //148 / 161 = 0
    16'b10010100_10100010 : OUT <= 0;  //148 / 162 = 0
    16'b10010100_10100011 : OUT <= 0;  //148 / 163 = 0
    16'b10010100_10100100 : OUT <= 0;  //148 / 164 = 0
    16'b10010100_10100101 : OUT <= 0;  //148 / 165 = 0
    16'b10010100_10100110 : OUT <= 0;  //148 / 166 = 0
    16'b10010100_10100111 : OUT <= 0;  //148 / 167 = 0
    16'b10010100_10101000 : OUT <= 0;  //148 / 168 = 0
    16'b10010100_10101001 : OUT <= 0;  //148 / 169 = 0
    16'b10010100_10101010 : OUT <= 0;  //148 / 170 = 0
    16'b10010100_10101011 : OUT <= 0;  //148 / 171 = 0
    16'b10010100_10101100 : OUT <= 0;  //148 / 172 = 0
    16'b10010100_10101101 : OUT <= 0;  //148 / 173 = 0
    16'b10010100_10101110 : OUT <= 0;  //148 / 174 = 0
    16'b10010100_10101111 : OUT <= 0;  //148 / 175 = 0
    16'b10010100_10110000 : OUT <= 0;  //148 / 176 = 0
    16'b10010100_10110001 : OUT <= 0;  //148 / 177 = 0
    16'b10010100_10110010 : OUT <= 0;  //148 / 178 = 0
    16'b10010100_10110011 : OUT <= 0;  //148 / 179 = 0
    16'b10010100_10110100 : OUT <= 0;  //148 / 180 = 0
    16'b10010100_10110101 : OUT <= 0;  //148 / 181 = 0
    16'b10010100_10110110 : OUT <= 0;  //148 / 182 = 0
    16'b10010100_10110111 : OUT <= 0;  //148 / 183 = 0
    16'b10010100_10111000 : OUT <= 0;  //148 / 184 = 0
    16'b10010100_10111001 : OUT <= 0;  //148 / 185 = 0
    16'b10010100_10111010 : OUT <= 0;  //148 / 186 = 0
    16'b10010100_10111011 : OUT <= 0;  //148 / 187 = 0
    16'b10010100_10111100 : OUT <= 0;  //148 / 188 = 0
    16'b10010100_10111101 : OUT <= 0;  //148 / 189 = 0
    16'b10010100_10111110 : OUT <= 0;  //148 / 190 = 0
    16'b10010100_10111111 : OUT <= 0;  //148 / 191 = 0
    16'b10010100_11000000 : OUT <= 0;  //148 / 192 = 0
    16'b10010100_11000001 : OUT <= 0;  //148 / 193 = 0
    16'b10010100_11000010 : OUT <= 0;  //148 / 194 = 0
    16'b10010100_11000011 : OUT <= 0;  //148 / 195 = 0
    16'b10010100_11000100 : OUT <= 0;  //148 / 196 = 0
    16'b10010100_11000101 : OUT <= 0;  //148 / 197 = 0
    16'b10010100_11000110 : OUT <= 0;  //148 / 198 = 0
    16'b10010100_11000111 : OUT <= 0;  //148 / 199 = 0
    16'b10010100_11001000 : OUT <= 0;  //148 / 200 = 0
    16'b10010100_11001001 : OUT <= 0;  //148 / 201 = 0
    16'b10010100_11001010 : OUT <= 0;  //148 / 202 = 0
    16'b10010100_11001011 : OUT <= 0;  //148 / 203 = 0
    16'b10010100_11001100 : OUT <= 0;  //148 / 204 = 0
    16'b10010100_11001101 : OUT <= 0;  //148 / 205 = 0
    16'b10010100_11001110 : OUT <= 0;  //148 / 206 = 0
    16'b10010100_11001111 : OUT <= 0;  //148 / 207 = 0
    16'b10010100_11010000 : OUT <= 0;  //148 / 208 = 0
    16'b10010100_11010001 : OUT <= 0;  //148 / 209 = 0
    16'b10010100_11010010 : OUT <= 0;  //148 / 210 = 0
    16'b10010100_11010011 : OUT <= 0;  //148 / 211 = 0
    16'b10010100_11010100 : OUT <= 0;  //148 / 212 = 0
    16'b10010100_11010101 : OUT <= 0;  //148 / 213 = 0
    16'b10010100_11010110 : OUT <= 0;  //148 / 214 = 0
    16'b10010100_11010111 : OUT <= 0;  //148 / 215 = 0
    16'b10010100_11011000 : OUT <= 0;  //148 / 216 = 0
    16'b10010100_11011001 : OUT <= 0;  //148 / 217 = 0
    16'b10010100_11011010 : OUT <= 0;  //148 / 218 = 0
    16'b10010100_11011011 : OUT <= 0;  //148 / 219 = 0
    16'b10010100_11011100 : OUT <= 0;  //148 / 220 = 0
    16'b10010100_11011101 : OUT <= 0;  //148 / 221 = 0
    16'b10010100_11011110 : OUT <= 0;  //148 / 222 = 0
    16'b10010100_11011111 : OUT <= 0;  //148 / 223 = 0
    16'b10010100_11100000 : OUT <= 0;  //148 / 224 = 0
    16'b10010100_11100001 : OUT <= 0;  //148 / 225 = 0
    16'b10010100_11100010 : OUT <= 0;  //148 / 226 = 0
    16'b10010100_11100011 : OUT <= 0;  //148 / 227 = 0
    16'b10010100_11100100 : OUT <= 0;  //148 / 228 = 0
    16'b10010100_11100101 : OUT <= 0;  //148 / 229 = 0
    16'b10010100_11100110 : OUT <= 0;  //148 / 230 = 0
    16'b10010100_11100111 : OUT <= 0;  //148 / 231 = 0
    16'b10010100_11101000 : OUT <= 0;  //148 / 232 = 0
    16'b10010100_11101001 : OUT <= 0;  //148 / 233 = 0
    16'b10010100_11101010 : OUT <= 0;  //148 / 234 = 0
    16'b10010100_11101011 : OUT <= 0;  //148 / 235 = 0
    16'b10010100_11101100 : OUT <= 0;  //148 / 236 = 0
    16'b10010100_11101101 : OUT <= 0;  //148 / 237 = 0
    16'b10010100_11101110 : OUT <= 0;  //148 / 238 = 0
    16'b10010100_11101111 : OUT <= 0;  //148 / 239 = 0
    16'b10010100_11110000 : OUT <= 0;  //148 / 240 = 0
    16'b10010100_11110001 : OUT <= 0;  //148 / 241 = 0
    16'b10010100_11110010 : OUT <= 0;  //148 / 242 = 0
    16'b10010100_11110011 : OUT <= 0;  //148 / 243 = 0
    16'b10010100_11110100 : OUT <= 0;  //148 / 244 = 0
    16'b10010100_11110101 : OUT <= 0;  //148 / 245 = 0
    16'b10010100_11110110 : OUT <= 0;  //148 / 246 = 0
    16'b10010100_11110111 : OUT <= 0;  //148 / 247 = 0
    16'b10010100_11111000 : OUT <= 0;  //148 / 248 = 0
    16'b10010100_11111001 : OUT <= 0;  //148 / 249 = 0
    16'b10010100_11111010 : OUT <= 0;  //148 / 250 = 0
    16'b10010100_11111011 : OUT <= 0;  //148 / 251 = 0
    16'b10010100_11111100 : OUT <= 0;  //148 / 252 = 0
    16'b10010100_11111101 : OUT <= 0;  //148 / 253 = 0
    16'b10010100_11111110 : OUT <= 0;  //148 / 254 = 0
    16'b10010100_11111111 : OUT <= 0;  //148 / 255 = 0
    16'b10010101_00000000 : OUT <= 0;  //149 / 0 = 0
    16'b10010101_00000001 : OUT <= 149;  //149 / 1 = 149
    16'b10010101_00000010 : OUT <= 74;  //149 / 2 = 74
    16'b10010101_00000011 : OUT <= 49;  //149 / 3 = 49
    16'b10010101_00000100 : OUT <= 37;  //149 / 4 = 37
    16'b10010101_00000101 : OUT <= 29;  //149 / 5 = 29
    16'b10010101_00000110 : OUT <= 24;  //149 / 6 = 24
    16'b10010101_00000111 : OUT <= 21;  //149 / 7 = 21
    16'b10010101_00001000 : OUT <= 18;  //149 / 8 = 18
    16'b10010101_00001001 : OUT <= 16;  //149 / 9 = 16
    16'b10010101_00001010 : OUT <= 14;  //149 / 10 = 14
    16'b10010101_00001011 : OUT <= 13;  //149 / 11 = 13
    16'b10010101_00001100 : OUT <= 12;  //149 / 12 = 12
    16'b10010101_00001101 : OUT <= 11;  //149 / 13 = 11
    16'b10010101_00001110 : OUT <= 10;  //149 / 14 = 10
    16'b10010101_00001111 : OUT <= 9;  //149 / 15 = 9
    16'b10010101_00010000 : OUT <= 9;  //149 / 16 = 9
    16'b10010101_00010001 : OUT <= 8;  //149 / 17 = 8
    16'b10010101_00010010 : OUT <= 8;  //149 / 18 = 8
    16'b10010101_00010011 : OUT <= 7;  //149 / 19 = 7
    16'b10010101_00010100 : OUT <= 7;  //149 / 20 = 7
    16'b10010101_00010101 : OUT <= 7;  //149 / 21 = 7
    16'b10010101_00010110 : OUT <= 6;  //149 / 22 = 6
    16'b10010101_00010111 : OUT <= 6;  //149 / 23 = 6
    16'b10010101_00011000 : OUT <= 6;  //149 / 24 = 6
    16'b10010101_00011001 : OUT <= 5;  //149 / 25 = 5
    16'b10010101_00011010 : OUT <= 5;  //149 / 26 = 5
    16'b10010101_00011011 : OUT <= 5;  //149 / 27 = 5
    16'b10010101_00011100 : OUT <= 5;  //149 / 28 = 5
    16'b10010101_00011101 : OUT <= 5;  //149 / 29 = 5
    16'b10010101_00011110 : OUT <= 4;  //149 / 30 = 4
    16'b10010101_00011111 : OUT <= 4;  //149 / 31 = 4
    16'b10010101_00100000 : OUT <= 4;  //149 / 32 = 4
    16'b10010101_00100001 : OUT <= 4;  //149 / 33 = 4
    16'b10010101_00100010 : OUT <= 4;  //149 / 34 = 4
    16'b10010101_00100011 : OUT <= 4;  //149 / 35 = 4
    16'b10010101_00100100 : OUT <= 4;  //149 / 36 = 4
    16'b10010101_00100101 : OUT <= 4;  //149 / 37 = 4
    16'b10010101_00100110 : OUT <= 3;  //149 / 38 = 3
    16'b10010101_00100111 : OUT <= 3;  //149 / 39 = 3
    16'b10010101_00101000 : OUT <= 3;  //149 / 40 = 3
    16'b10010101_00101001 : OUT <= 3;  //149 / 41 = 3
    16'b10010101_00101010 : OUT <= 3;  //149 / 42 = 3
    16'b10010101_00101011 : OUT <= 3;  //149 / 43 = 3
    16'b10010101_00101100 : OUT <= 3;  //149 / 44 = 3
    16'b10010101_00101101 : OUT <= 3;  //149 / 45 = 3
    16'b10010101_00101110 : OUT <= 3;  //149 / 46 = 3
    16'b10010101_00101111 : OUT <= 3;  //149 / 47 = 3
    16'b10010101_00110000 : OUT <= 3;  //149 / 48 = 3
    16'b10010101_00110001 : OUT <= 3;  //149 / 49 = 3
    16'b10010101_00110010 : OUT <= 2;  //149 / 50 = 2
    16'b10010101_00110011 : OUT <= 2;  //149 / 51 = 2
    16'b10010101_00110100 : OUT <= 2;  //149 / 52 = 2
    16'b10010101_00110101 : OUT <= 2;  //149 / 53 = 2
    16'b10010101_00110110 : OUT <= 2;  //149 / 54 = 2
    16'b10010101_00110111 : OUT <= 2;  //149 / 55 = 2
    16'b10010101_00111000 : OUT <= 2;  //149 / 56 = 2
    16'b10010101_00111001 : OUT <= 2;  //149 / 57 = 2
    16'b10010101_00111010 : OUT <= 2;  //149 / 58 = 2
    16'b10010101_00111011 : OUT <= 2;  //149 / 59 = 2
    16'b10010101_00111100 : OUT <= 2;  //149 / 60 = 2
    16'b10010101_00111101 : OUT <= 2;  //149 / 61 = 2
    16'b10010101_00111110 : OUT <= 2;  //149 / 62 = 2
    16'b10010101_00111111 : OUT <= 2;  //149 / 63 = 2
    16'b10010101_01000000 : OUT <= 2;  //149 / 64 = 2
    16'b10010101_01000001 : OUT <= 2;  //149 / 65 = 2
    16'b10010101_01000010 : OUT <= 2;  //149 / 66 = 2
    16'b10010101_01000011 : OUT <= 2;  //149 / 67 = 2
    16'b10010101_01000100 : OUT <= 2;  //149 / 68 = 2
    16'b10010101_01000101 : OUT <= 2;  //149 / 69 = 2
    16'b10010101_01000110 : OUT <= 2;  //149 / 70 = 2
    16'b10010101_01000111 : OUT <= 2;  //149 / 71 = 2
    16'b10010101_01001000 : OUT <= 2;  //149 / 72 = 2
    16'b10010101_01001001 : OUT <= 2;  //149 / 73 = 2
    16'b10010101_01001010 : OUT <= 2;  //149 / 74 = 2
    16'b10010101_01001011 : OUT <= 1;  //149 / 75 = 1
    16'b10010101_01001100 : OUT <= 1;  //149 / 76 = 1
    16'b10010101_01001101 : OUT <= 1;  //149 / 77 = 1
    16'b10010101_01001110 : OUT <= 1;  //149 / 78 = 1
    16'b10010101_01001111 : OUT <= 1;  //149 / 79 = 1
    16'b10010101_01010000 : OUT <= 1;  //149 / 80 = 1
    16'b10010101_01010001 : OUT <= 1;  //149 / 81 = 1
    16'b10010101_01010010 : OUT <= 1;  //149 / 82 = 1
    16'b10010101_01010011 : OUT <= 1;  //149 / 83 = 1
    16'b10010101_01010100 : OUT <= 1;  //149 / 84 = 1
    16'b10010101_01010101 : OUT <= 1;  //149 / 85 = 1
    16'b10010101_01010110 : OUT <= 1;  //149 / 86 = 1
    16'b10010101_01010111 : OUT <= 1;  //149 / 87 = 1
    16'b10010101_01011000 : OUT <= 1;  //149 / 88 = 1
    16'b10010101_01011001 : OUT <= 1;  //149 / 89 = 1
    16'b10010101_01011010 : OUT <= 1;  //149 / 90 = 1
    16'b10010101_01011011 : OUT <= 1;  //149 / 91 = 1
    16'b10010101_01011100 : OUT <= 1;  //149 / 92 = 1
    16'b10010101_01011101 : OUT <= 1;  //149 / 93 = 1
    16'b10010101_01011110 : OUT <= 1;  //149 / 94 = 1
    16'b10010101_01011111 : OUT <= 1;  //149 / 95 = 1
    16'b10010101_01100000 : OUT <= 1;  //149 / 96 = 1
    16'b10010101_01100001 : OUT <= 1;  //149 / 97 = 1
    16'b10010101_01100010 : OUT <= 1;  //149 / 98 = 1
    16'b10010101_01100011 : OUT <= 1;  //149 / 99 = 1
    16'b10010101_01100100 : OUT <= 1;  //149 / 100 = 1
    16'b10010101_01100101 : OUT <= 1;  //149 / 101 = 1
    16'b10010101_01100110 : OUT <= 1;  //149 / 102 = 1
    16'b10010101_01100111 : OUT <= 1;  //149 / 103 = 1
    16'b10010101_01101000 : OUT <= 1;  //149 / 104 = 1
    16'b10010101_01101001 : OUT <= 1;  //149 / 105 = 1
    16'b10010101_01101010 : OUT <= 1;  //149 / 106 = 1
    16'b10010101_01101011 : OUT <= 1;  //149 / 107 = 1
    16'b10010101_01101100 : OUT <= 1;  //149 / 108 = 1
    16'b10010101_01101101 : OUT <= 1;  //149 / 109 = 1
    16'b10010101_01101110 : OUT <= 1;  //149 / 110 = 1
    16'b10010101_01101111 : OUT <= 1;  //149 / 111 = 1
    16'b10010101_01110000 : OUT <= 1;  //149 / 112 = 1
    16'b10010101_01110001 : OUT <= 1;  //149 / 113 = 1
    16'b10010101_01110010 : OUT <= 1;  //149 / 114 = 1
    16'b10010101_01110011 : OUT <= 1;  //149 / 115 = 1
    16'b10010101_01110100 : OUT <= 1;  //149 / 116 = 1
    16'b10010101_01110101 : OUT <= 1;  //149 / 117 = 1
    16'b10010101_01110110 : OUT <= 1;  //149 / 118 = 1
    16'b10010101_01110111 : OUT <= 1;  //149 / 119 = 1
    16'b10010101_01111000 : OUT <= 1;  //149 / 120 = 1
    16'b10010101_01111001 : OUT <= 1;  //149 / 121 = 1
    16'b10010101_01111010 : OUT <= 1;  //149 / 122 = 1
    16'b10010101_01111011 : OUT <= 1;  //149 / 123 = 1
    16'b10010101_01111100 : OUT <= 1;  //149 / 124 = 1
    16'b10010101_01111101 : OUT <= 1;  //149 / 125 = 1
    16'b10010101_01111110 : OUT <= 1;  //149 / 126 = 1
    16'b10010101_01111111 : OUT <= 1;  //149 / 127 = 1
    16'b10010101_10000000 : OUT <= 1;  //149 / 128 = 1
    16'b10010101_10000001 : OUT <= 1;  //149 / 129 = 1
    16'b10010101_10000010 : OUT <= 1;  //149 / 130 = 1
    16'b10010101_10000011 : OUT <= 1;  //149 / 131 = 1
    16'b10010101_10000100 : OUT <= 1;  //149 / 132 = 1
    16'b10010101_10000101 : OUT <= 1;  //149 / 133 = 1
    16'b10010101_10000110 : OUT <= 1;  //149 / 134 = 1
    16'b10010101_10000111 : OUT <= 1;  //149 / 135 = 1
    16'b10010101_10001000 : OUT <= 1;  //149 / 136 = 1
    16'b10010101_10001001 : OUT <= 1;  //149 / 137 = 1
    16'b10010101_10001010 : OUT <= 1;  //149 / 138 = 1
    16'b10010101_10001011 : OUT <= 1;  //149 / 139 = 1
    16'b10010101_10001100 : OUT <= 1;  //149 / 140 = 1
    16'b10010101_10001101 : OUT <= 1;  //149 / 141 = 1
    16'b10010101_10001110 : OUT <= 1;  //149 / 142 = 1
    16'b10010101_10001111 : OUT <= 1;  //149 / 143 = 1
    16'b10010101_10010000 : OUT <= 1;  //149 / 144 = 1
    16'b10010101_10010001 : OUT <= 1;  //149 / 145 = 1
    16'b10010101_10010010 : OUT <= 1;  //149 / 146 = 1
    16'b10010101_10010011 : OUT <= 1;  //149 / 147 = 1
    16'b10010101_10010100 : OUT <= 1;  //149 / 148 = 1
    16'b10010101_10010101 : OUT <= 1;  //149 / 149 = 1
    16'b10010101_10010110 : OUT <= 0;  //149 / 150 = 0
    16'b10010101_10010111 : OUT <= 0;  //149 / 151 = 0
    16'b10010101_10011000 : OUT <= 0;  //149 / 152 = 0
    16'b10010101_10011001 : OUT <= 0;  //149 / 153 = 0
    16'b10010101_10011010 : OUT <= 0;  //149 / 154 = 0
    16'b10010101_10011011 : OUT <= 0;  //149 / 155 = 0
    16'b10010101_10011100 : OUT <= 0;  //149 / 156 = 0
    16'b10010101_10011101 : OUT <= 0;  //149 / 157 = 0
    16'b10010101_10011110 : OUT <= 0;  //149 / 158 = 0
    16'b10010101_10011111 : OUT <= 0;  //149 / 159 = 0
    16'b10010101_10100000 : OUT <= 0;  //149 / 160 = 0
    16'b10010101_10100001 : OUT <= 0;  //149 / 161 = 0
    16'b10010101_10100010 : OUT <= 0;  //149 / 162 = 0
    16'b10010101_10100011 : OUT <= 0;  //149 / 163 = 0
    16'b10010101_10100100 : OUT <= 0;  //149 / 164 = 0
    16'b10010101_10100101 : OUT <= 0;  //149 / 165 = 0
    16'b10010101_10100110 : OUT <= 0;  //149 / 166 = 0
    16'b10010101_10100111 : OUT <= 0;  //149 / 167 = 0
    16'b10010101_10101000 : OUT <= 0;  //149 / 168 = 0
    16'b10010101_10101001 : OUT <= 0;  //149 / 169 = 0
    16'b10010101_10101010 : OUT <= 0;  //149 / 170 = 0
    16'b10010101_10101011 : OUT <= 0;  //149 / 171 = 0
    16'b10010101_10101100 : OUT <= 0;  //149 / 172 = 0
    16'b10010101_10101101 : OUT <= 0;  //149 / 173 = 0
    16'b10010101_10101110 : OUT <= 0;  //149 / 174 = 0
    16'b10010101_10101111 : OUT <= 0;  //149 / 175 = 0
    16'b10010101_10110000 : OUT <= 0;  //149 / 176 = 0
    16'b10010101_10110001 : OUT <= 0;  //149 / 177 = 0
    16'b10010101_10110010 : OUT <= 0;  //149 / 178 = 0
    16'b10010101_10110011 : OUT <= 0;  //149 / 179 = 0
    16'b10010101_10110100 : OUT <= 0;  //149 / 180 = 0
    16'b10010101_10110101 : OUT <= 0;  //149 / 181 = 0
    16'b10010101_10110110 : OUT <= 0;  //149 / 182 = 0
    16'b10010101_10110111 : OUT <= 0;  //149 / 183 = 0
    16'b10010101_10111000 : OUT <= 0;  //149 / 184 = 0
    16'b10010101_10111001 : OUT <= 0;  //149 / 185 = 0
    16'b10010101_10111010 : OUT <= 0;  //149 / 186 = 0
    16'b10010101_10111011 : OUT <= 0;  //149 / 187 = 0
    16'b10010101_10111100 : OUT <= 0;  //149 / 188 = 0
    16'b10010101_10111101 : OUT <= 0;  //149 / 189 = 0
    16'b10010101_10111110 : OUT <= 0;  //149 / 190 = 0
    16'b10010101_10111111 : OUT <= 0;  //149 / 191 = 0
    16'b10010101_11000000 : OUT <= 0;  //149 / 192 = 0
    16'b10010101_11000001 : OUT <= 0;  //149 / 193 = 0
    16'b10010101_11000010 : OUT <= 0;  //149 / 194 = 0
    16'b10010101_11000011 : OUT <= 0;  //149 / 195 = 0
    16'b10010101_11000100 : OUT <= 0;  //149 / 196 = 0
    16'b10010101_11000101 : OUT <= 0;  //149 / 197 = 0
    16'b10010101_11000110 : OUT <= 0;  //149 / 198 = 0
    16'b10010101_11000111 : OUT <= 0;  //149 / 199 = 0
    16'b10010101_11001000 : OUT <= 0;  //149 / 200 = 0
    16'b10010101_11001001 : OUT <= 0;  //149 / 201 = 0
    16'b10010101_11001010 : OUT <= 0;  //149 / 202 = 0
    16'b10010101_11001011 : OUT <= 0;  //149 / 203 = 0
    16'b10010101_11001100 : OUT <= 0;  //149 / 204 = 0
    16'b10010101_11001101 : OUT <= 0;  //149 / 205 = 0
    16'b10010101_11001110 : OUT <= 0;  //149 / 206 = 0
    16'b10010101_11001111 : OUT <= 0;  //149 / 207 = 0
    16'b10010101_11010000 : OUT <= 0;  //149 / 208 = 0
    16'b10010101_11010001 : OUT <= 0;  //149 / 209 = 0
    16'b10010101_11010010 : OUT <= 0;  //149 / 210 = 0
    16'b10010101_11010011 : OUT <= 0;  //149 / 211 = 0
    16'b10010101_11010100 : OUT <= 0;  //149 / 212 = 0
    16'b10010101_11010101 : OUT <= 0;  //149 / 213 = 0
    16'b10010101_11010110 : OUT <= 0;  //149 / 214 = 0
    16'b10010101_11010111 : OUT <= 0;  //149 / 215 = 0
    16'b10010101_11011000 : OUT <= 0;  //149 / 216 = 0
    16'b10010101_11011001 : OUT <= 0;  //149 / 217 = 0
    16'b10010101_11011010 : OUT <= 0;  //149 / 218 = 0
    16'b10010101_11011011 : OUT <= 0;  //149 / 219 = 0
    16'b10010101_11011100 : OUT <= 0;  //149 / 220 = 0
    16'b10010101_11011101 : OUT <= 0;  //149 / 221 = 0
    16'b10010101_11011110 : OUT <= 0;  //149 / 222 = 0
    16'b10010101_11011111 : OUT <= 0;  //149 / 223 = 0
    16'b10010101_11100000 : OUT <= 0;  //149 / 224 = 0
    16'b10010101_11100001 : OUT <= 0;  //149 / 225 = 0
    16'b10010101_11100010 : OUT <= 0;  //149 / 226 = 0
    16'b10010101_11100011 : OUT <= 0;  //149 / 227 = 0
    16'b10010101_11100100 : OUT <= 0;  //149 / 228 = 0
    16'b10010101_11100101 : OUT <= 0;  //149 / 229 = 0
    16'b10010101_11100110 : OUT <= 0;  //149 / 230 = 0
    16'b10010101_11100111 : OUT <= 0;  //149 / 231 = 0
    16'b10010101_11101000 : OUT <= 0;  //149 / 232 = 0
    16'b10010101_11101001 : OUT <= 0;  //149 / 233 = 0
    16'b10010101_11101010 : OUT <= 0;  //149 / 234 = 0
    16'b10010101_11101011 : OUT <= 0;  //149 / 235 = 0
    16'b10010101_11101100 : OUT <= 0;  //149 / 236 = 0
    16'b10010101_11101101 : OUT <= 0;  //149 / 237 = 0
    16'b10010101_11101110 : OUT <= 0;  //149 / 238 = 0
    16'b10010101_11101111 : OUT <= 0;  //149 / 239 = 0
    16'b10010101_11110000 : OUT <= 0;  //149 / 240 = 0
    16'b10010101_11110001 : OUT <= 0;  //149 / 241 = 0
    16'b10010101_11110010 : OUT <= 0;  //149 / 242 = 0
    16'b10010101_11110011 : OUT <= 0;  //149 / 243 = 0
    16'b10010101_11110100 : OUT <= 0;  //149 / 244 = 0
    16'b10010101_11110101 : OUT <= 0;  //149 / 245 = 0
    16'b10010101_11110110 : OUT <= 0;  //149 / 246 = 0
    16'b10010101_11110111 : OUT <= 0;  //149 / 247 = 0
    16'b10010101_11111000 : OUT <= 0;  //149 / 248 = 0
    16'b10010101_11111001 : OUT <= 0;  //149 / 249 = 0
    16'b10010101_11111010 : OUT <= 0;  //149 / 250 = 0
    16'b10010101_11111011 : OUT <= 0;  //149 / 251 = 0
    16'b10010101_11111100 : OUT <= 0;  //149 / 252 = 0
    16'b10010101_11111101 : OUT <= 0;  //149 / 253 = 0
    16'b10010101_11111110 : OUT <= 0;  //149 / 254 = 0
    16'b10010101_11111111 : OUT <= 0;  //149 / 255 = 0
    16'b10010110_00000000 : OUT <= 0;  //150 / 0 = 0
    16'b10010110_00000001 : OUT <= 150;  //150 / 1 = 150
    16'b10010110_00000010 : OUT <= 75;  //150 / 2 = 75
    16'b10010110_00000011 : OUT <= 50;  //150 / 3 = 50
    16'b10010110_00000100 : OUT <= 37;  //150 / 4 = 37
    16'b10010110_00000101 : OUT <= 30;  //150 / 5 = 30
    16'b10010110_00000110 : OUT <= 25;  //150 / 6 = 25
    16'b10010110_00000111 : OUT <= 21;  //150 / 7 = 21
    16'b10010110_00001000 : OUT <= 18;  //150 / 8 = 18
    16'b10010110_00001001 : OUT <= 16;  //150 / 9 = 16
    16'b10010110_00001010 : OUT <= 15;  //150 / 10 = 15
    16'b10010110_00001011 : OUT <= 13;  //150 / 11 = 13
    16'b10010110_00001100 : OUT <= 12;  //150 / 12 = 12
    16'b10010110_00001101 : OUT <= 11;  //150 / 13 = 11
    16'b10010110_00001110 : OUT <= 10;  //150 / 14 = 10
    16'b10010110_00001111 : OUT <= 10;  //150 / 15 = 10
    16'b10010110_00010000 : OUT <= 9;  //150 / 16 = 9
    16'b10010110_00010001 : OUT <= 8;  //150 / 17 = 8
    16'b10010110_00010010 : OUT <= 8;  //150 / 18 = 8
    16'b10010110_00010011 : OUT <= 7;  //150 / 19 = 7
    16'b10010110_00010100 : OUT <= 7;  //150 / 20 = 7
    16'b10010110_00010101 : OUT <= 7;  //150 / 21 = 7
    16'b10010110_00010110 : OUT <= 6;  //150 / 22 = 6
    16'b10010110_00010111 : OUT <= 6;  //150 / 23 = 6
    16'b10010110_00011000 : OUT <= 6;  //150 / 24 = 6
    16'b10010110_00011001 : OUT <= 6;  //150 / 25 = 6
    16'b10010110_00011010 : OUT <= 5;  //150 / 26 = 5
    16'b10010110_00011011 : OUT <= 5;  //150 / 27 = 5
    16'b10010110_00011100 : OUT <= 5;  //150 / 28 = 5
    16'b10010110_00011101 : OUT <= 5;  //150 / 29 = 5
    16'b10010110_00011110 : OUT <= 5;  //150 / 30 = 5
    16'b10010110_00011111 : OUT <= 4;  //150 / 31 = 4
    16'b10010110_00100000 : OUT <= 4;  //150 / 32 = 4
    16'b10010110_00100001 : OUT <= 4;  //150 / 33 = 4
    16'b10010110_00100010 : OUT <= 4;  //150 / 34 = 4
    16'b10010110_00100011 : OUT <= 4;  //150 / 35 = 4
    16'b10010110_00100100 : OUT <= 4;  //150 / 36 = 4
    16'b10010110_00100101 : OUT <= 4;  //150 / 37 = 4
    16'b10010110_00100110 : OUT <= 3;  //150 / 38 = 3
    16'b10010110_00100111 : OUT <= 3;  //150 / 39 = 3
    16'b10010110_00101000 : OUT <= 3;  //150 / 40 = 3
    16'b10010110_00101001 : OUT <= 3;  //150 / 41 = 3
    16'b10010110_00101010 : OUT <= 3;  //150 / 42 = 3
    16'b10010110_00101011 : OUT <= 3;  //150 / 43 = 3
    16'b10010110_00101100 : OUT <= 3;  //150 / 44 = 3
    16'b10010110_00101101 : OUT <= 3;  //150 / 45 = 3
    16'b10010110_00101110 : OUT <= 3;  //150 / 46 = 3
    16'b10010110_00101111 : OUT <= 3;  //150 / 47 = 3
    16'b10010110_00110000 : OUT <= 3;  //150 / 48 = 3
    16'b10010110_00110001 : OUT <= 3;  //150 / 49 = 3
    16'b10010110_00110010 : OUT <= 3;  //150 / 50 = 3
    16'b10010110_00110011 : OUT <= 2;  //150 / 51 = 2
    16'b10010110_00110100 : OUT <= 2;  //150 / 52 = 2
    16'b10010110_00110101 : OUT <= 2;  //150 / 53 = 2
    16'b10010110_00110110 : OUT <= 2;  //150 / 54 = 2
    16'b10010110_00110111 : OUT <= 2;  //150 / 55 = 2
    16'b10010110_00111000 : OUT <= 2;  //150 / 56 = 2
    16'b10010110_00111001 : OUT <= 2;  //150 / 57 = 2
    16'b10010110_00111010 : OUT <= 2;  //150 / 58 = 2
    16'b10010110_00111011 : OUT <= 2;  //150 / 59 = 2
    16'b10010110_00111100 : OUT <= 2;  //150 / 60 = 2
    16'b10010110_00111101 : OUT <= 2;  //150 / 61 = 2
    16'b10010110_00111110 : OUT <= 2;  //150 / 62 = 2
    16'b10010110_00111111 : OUT <= 2;  //150 / 63 = 2
    16'b10010110_01000000 : OUT <= 2;  //150 / 64 = 2
    16'b10010110_01000001 : OUT <= 2;  //150 / 65 = 2
    16'b10010110_01000010 : OUT <= 2;  //150 / 66 = 2
    16'b10010110_01000011 : OUT <= 2;  //150 / 67 = 2
    16'b10010110_01000100 : OUT <= 2;  //150 / 68 = 2
    16'b10010110_01000101 : OUT <= 2;  //150 / 69 = 2
    16'b10010110_01000110 : OUT <= 2;  //150 / 70 = 2
    16'b10010110_01000111 : OUT <= 2;  //150 / 71 = 2
    16'b10010110_01001000 : OUT <= 2;  //150 / 72 = 2
    16'b10010110_01001001 : OUT <= 2;  //150 / 73 = 2
    16'b10010110_01001010 : OUT <= 2;  //150 / 74 = 2
    16'b10010110_01001011 : OUT <= 2;  //150 / 75 = 2
    16'b10010110_01001100 : OUT <= 1;  //150 / 76 = 1
    16'b10010110_01001101 : OUT <= 1;  //150 / 77 = 1
    16'b10010110_01001110 : OUT <= 1;  //150 / 78 = 1
    16'b10010110_01001111 : OUT <= 1;  //150 / 79 = 1
    16'b10010110_01010000 : OUT <= 1;  //150 / 80 = 1
    16'b10010110_01010001 : OUT <= 1;  //150 / 81 = 1
    16'b10010110_01010010 : OUT <= 1;  //150 / 82 = 1
    16'b10010110_01010011 : OUT <= 1;  //150 / 83 = 1
    16'b10010110_01010100 : OUT <= 1;  //150 / 84 = 1
    16'b10010110_01010101 : OUT <= 1;  //150 / 85 = 1
    16'b10010110_01010110 : OUT <= 1;  //150 / 86 = 1
    16'b10010110_01010111 : OUT <= 1;  //150 / 87 = 1
    16'b10010110_01011000 : OUT <= 1;  //150 / 88 = 1
    16'b10010110_01011001 : OUT <= 1;  //150 / 89 = 1
    16'b10010110_01011010 : OUT <= 1;  //150 / 90 = 1
    16'b10010110_01011011 : OUT <= 1;  //150 / 91 = 1
    16'b10010110_01011100 : OUT <= 1;  //150 / 92 = 1
    16'b10010110_01011101 : OUT <= 1;  //150 / 93 = 1
    16'b10010110_01011110 : OUT <= 1;  //150 / 94 = 1
    16'b10010110_01011111 : OUT <= 1;  //150 / 95 = 1
    16'b10010110_01100000 : OUT <= 1;  //150 / 96 = 1
    16'b10010110_01100001 : OUT <= 1;  //150 / 97 = 1
    16'b10010110_01100010 : OUT <= 1;  //150 / 98 = 1
    16'b10010110_01100011 : OUT <= 1;  //150 / 99 = 1
    16'b10010110_01100100 : OUT <= 1;  //150 / 100 = 1
    16'b10010110_01100101 : OUT <= 1;  //150 / 101 = 1
    16'b10010110_01100110 : OUT <= 1;  //150 / 102 = 1
    16'b10010110_01100111 : OUT <= 1;  //150 / 103 = 1
    16'b10010110_01101000 : OUT <= 1;  //150 / 104 = 1
    16'b10010110_01101001 : OUT <= 1;  //150 / 105 = 1
    16'b10010110_01101010 : OUT <= 1;  //150 / 106 = 1
    16'b10010110_01101011 : OUT <= 1;  //150 / 107 = 1
    16'b10010110_01101100 : OUT <= 1;  //150 / 108 = 1
    16'b10010110_01101101 : OUT <= 1;  //150 / 109 = 1
    16'b10010110_01101110 : OUT <= 1;  //150 / 110 = 1
    16'b10010110_01101111 : OUT <= 1;  //150 / 111 = 1
    16'b10010110_01110000 : OUT <= 1;  //150 / 112 = 1
    16'b10010110_01110001 : OUT <= 1;  //150 / 113 = 1
    16'b10010110_01110010 : OUT <= 1;  //150 / 114 = 1
    16'b10010110_01110011 : OUT <= 1;  //150 / 115 = 1
    16'b10010110_01110100 : OUT <= 1;  //150 / 116 = 1
    16'b10010110_01110101 : OUT <= 1;  //150 / 117 = 1
    16'b10010110_01110110 : OUT <= 1;  //150 / 118 = 1
    16'b10010110_01110111 : OUT <= 1;  //150 / 119 = 1
    16'b10010110_01111000 : OUT <= 1;  //150 / 120 = 1
    16'b10010110_01111001 : OUT <= 1;  //150 / 121 = 1
    16'b10010110_01111010 : OUT <= 1;  //150 / 122 = 1
    16'b10010110_01111011 : OUT <= 1;  //150 / 123 = 1
    16'b10010110_01111100 : OUT <= 1;  //150 / 124 = 1
    16'b10010110_01111101 : OUT <= 1;  //150 / 125 = 1
    16'b10010110_01111110 : OUT <= 1;  //150 / 126 = 1
    16'b10010110_01111111 : OUT <= 1;  //150 / 127 = 1
    16'b10010110_10000000 : OUT <= 1;  //150 / 128 = 1
    16'b10010110_10000001 : OUT <= 1;  //150 / 129 = 1
    16'b10010110_10000010 : OUT <= 1;  //150 / 130 = 1
    16'b10010110_10000011 : OUT <= 1;  //150 / 131 = 1
    16'b10010110_10000100 : OUT <= 1;  //150 / 132 = 1
    16'b10010110_10000101 : OUT <= 1;  //150 / 133 = 1
    16'b10010110_10000110 : OUT <= 1;  //150 / 134 = 1
    16'b10010110_10000111 : OUT <= 1;  //150 / 135 = 1
    16'b10010110_10001000 : OUT <= 1;  //150 / 136 = 1
    16'b10010110_10001001 : OUT <= 1;  //150 / 137 = 1
    16'b10010110_10001010 : OUT <= 1;  //150 / 138 = 1
    16'b10010110_10001011 : OUT <= 1;  //150 / 139 = 1
    16'b10010110_10001100 : OUT <= 1;  //150 / 140 = 1
    16'b10010110_10001101 : OUT <= 1;  //150 / 141 = 1
    16'b10010110_10001110 : OUT <= 1;  //150 / 142 = 1
    16'b10010110_10001111 : OUT <= 1;  //150 / 143 = 1
    16'b10010110_10010000 : OUT <= 1;  //150 / 144 = 1
    16'b10010110_10010001 : OUT <= 1;  //150 / 145 = 1
    16'b10010110_10010010 : OUT <= 1;  //150 / 146 = 1
    16'b10010110_10010011 : OUT <= 1;  //150 / 147 = 1
    16'b10010110_10010100 : OUT <= 1;  //150 / 148 = 1
    16'b10010110_10010101 : OUT <= 1;  //150 / 149 = 1
    16'b10010110_10010110 : OUT <= 1;  //150 / 150 = 1
    16'b10010110_10010111 : OUT <= 0;  //150 / 151 = 0
    16'b10010110_10011000 : OUT <= 0;  //150 / 152 = 0
    16'b10010110_10011001 : OUT <= 0;  //150 / 153 = 0
    16'b10010110_10011010 : OUT <= 0;  //150 / 154 = 0
    16'b10010110_10011011 : OUT <= 0;  //150 / 155 = 0
    16'b10010110_10011100 : OUT <= 0;  //150 / 156 = 0
    16'b10010110_10011101 : OUT <= 0;  //150 / 157 = 0
    16'b10010110_10011110 : OUT <= 0;  //150 / 158 = 0
    16'b10010110_10011111 : OUT <= 0;  //150 / 159 = 0
    16'b10010110_10100000 : OUT <= 0;  //150 / 160 = 0
    16'b10010110_10100001 : OUT <= 0;  //150 / 161 = 0
    16'b10010110_10100010 : OUT <= 0;  //150 / 162 = 0
    16'b10010110_10100011 : OUT <= 0;  //150 / 163 = 0
    16'b10010110_10100100 : OUT <= 0;  //150 / 164 = 0
    16'b10010110_10100101 : OUT <= 0;  //150 / 165 = 0
    16'b10010110_10100110 : OUT <= 0;  //150 / 166 = 0
    16'b10010110_10100111 : OUT <= 0;  //150 / 167 = 0
    16'b10010110_10101000 : OUT <= 0;  //150 / 168 = 0
    16'b10010110_10101001 : OUT <= 0;  //150 / 169 = 0
    16'b10010110_10101010 : OUT <= 0;  //150 / 170 = 0
    16'b10010110_10101011 : OUT <= 0;  //150 / 171 = 0
    16'b10010110_10101100 : OUT <= 0;  //150 / 172 = 0
    16'b10010110_10101101 : OUT <= 0;  //150 / 173 = 0
    16'b10010110_10101110 : OUT <= 0;  //150 / 174 = 0
    16'b10010110_10101111 : OUT <= 0;  //150 / 175 = 0
    16'b10010110_10110000 : OUT <= 0;  //150 / 176 = 0
    16'b10010110_10110001 : OUT <= 0;  //150 / 177 = 0
    16'b10010110_10110010 : OUT <= 0;  //150 / 178 = 0
    16'b10010110_10110011 : OUT <= 0;  //150 / 179 = 0
    16'b10010110_10110100 : OUT <= 0;  //150 / 180 = 0
    16'b10010110_10110101 : OUT <= 0;  //150 / 181 = 0
    16'b10010110_10110110 : OUT <= 0;  //150 / 182 = 0
    16'b10010110_10110111 : OUT <= 0;  //150 / 183 = 0
    16'b10010110_10111000 : OUT <= 0;  //150 / 184 = 0
    16'b10010110_10111001 : OUT <= 0;  //150 / 185 = 0
    16'b10010110_10111010 : OUT <= 0;  //150 / 186 = 0
    16'b10010110_10111011 : OUT <= 0;  //150 / 187 = 0
    16'b10010110_10111100 : OUT <= 0;  //150 / 188 = 0
    16'b10010110_10111101 : OUT <= 0;  //150 / 189 = 0
    16'b10010110_10111110 : OUT <= 0;  //150 / 190 = 0
    16'b10010110_10111111 : OUT <= 0;  //150 / 191 = 0
    16'b10010110_11000000 : OUT <= 0;  //150 / 192 = 0
    16'b10010110_11000001 : OUT <= 0;  //150 / 193 = 0
    16'b10010110_11000010 : OUT <= 0;  //150 / 194 = 0
    16'b10010110_11000011 : OUT <= 0;  //150 / 195 = 0
    16'b10010110_11000100 : OUT <= 0;  //150 / 196 = 0
    16'b10010110_11000101 : OUT <= 0;  //150 / 197 = 0
    16'b10010110_11000110 : OUT <= 0;  //150 / 198 = 0
    16'b10010110_11000111 : OUT <= 0;  //150 / 199 = 0
    16'b10010110_11001000 : OUT <= 0;  //150 / 200 = 0
    16'b10010110_11001001 : OUT <= 0;  //150 / 201 = 0
    16'b10010110_11001010 : OUT <= 0;  //150 / 202 = 0
    16'b10010110_11001011 : OUT <= 0;  //150 / 203 = 0
    16'b10010110_11001100 : OUT <= 0;  //150 / 204 = 0
    16'b10010110_11001101 : OUT <= 0;  //150 / 205 = 0
    16'b10010110_11001110 : OUT <= 0;  //150 / 206 = 0
    16'b10010110_11001111 : OUT <= 0;  //150 / 207 = 0
    16'b10010110_11010000 : OUT <= 0;  //150 / 208 = 0
    16'b10010110_11010001 : OUT <= 0;  //150 / 209 = 0
    16'b10010110_11010010 : OUT <= 0;  //150 / 210 = 0
    16'b10010110_11010011 : OUT <= 0;  //150 / 211 = 0
    16'b10010110_11010100 : OUT <= 0;  //150 / 212 = 0
    16'b10010110_11010101 : OUT <= 0;  //150 / 213 = 0
    16'b10010110_11010110 : OUT <= 0;  //150 / 214 = 0
    16'b10010110_11010111 : OUT <= 0;  //150 / 215 = 0
    16'b10010110_11011000 : OUT <= 0;  //150 / 216 = 0
    16'b10010110_11011001 : OUT <= 0;  //150 / 217 = 0
    16'b10010110_11011010 : OUT <= 0;  //150 / 218 = 0
    16'b10010110_11011011 : OUT <= 0;  //150 / 219 = 0
    16'b10010110_11011100 : OUT <= 0;  //150 / 220 = 0
    16'b10010110_11011101 : OUT <= 0;  //150 / 221 = 0
    16'b10010110_11011110 : OUT <= 0;  //150 / 222 = 0
    16'b10010110_11011111 : OUT <= 0;  //150 / 223 = 0
    16'b10010110_11100000 : OUT <= 0;  //150 / 224 = 0
    16'b10010110_11100001 : OUT <= 0;  //150 / 225 = 0
    16'b10010110_11100010 : OUT <= 0;  //150 / 226 = 0
    16'b10010110_11100011 : OUT <= 0;  //150 / 227 = 0
    16'b10010110_11100100 : OUT <= 0;  //150 / 228 = 0
    16'b10010110_11100101 : OUT <= 0;  //150 / 229 = 0
    16'b10010110_11100110 : OUT <= 0;  //150 / 230 = 0
    16'b10010110_11100111 : OUT <= 0;  //150 / 231 = 0
    16'b10010110_11101000 : OUT <= 0;  //150 / 232 = 0
    16'b10010110_11101001 : OUT <= 0;  //150 / 233 = 0
    16'b10010110_11101010 : OUT <= 0;  //150 / 234 = 0
    16'b10010110_11101011 : OUT <= 0;  //150 / 235 = 0
    16'b10010110_11101100 : OUT <= 0;  //150 / 236 = 0
    16'b10010110_11101101 : OUT <= 0;  //150 / 237 = 0
    16'b10010110_11101110 : OUT <= 0;  //150 / 238 = 0
    16'b10010110_11101111 : OUT <= 0;  //150 / 239 = 0
    16'b10010110_11110000 : OUT <= 0;  //150 / 240 = 0
    16'b10010110_11110001 : OUT <= 0;  //150 / 241 = 0
    16'b10010110_11110010 : OUT <= 0;  //150 / 242 = 0
    16'b10010110_11110011 : OUT <= 0;  //150 / 243 = 0
    16'b10010110_11110100 : OUT <= 0;  //150 / 244 = 0
    16'b10010110_11110101 : OUT <= 0;  //150 / 245 = 0
    16'b10010110_11110110 : OUT <= 0;  //150 / 246 = 0
    16'b10010110_11110111 : OUT <= 0;  //150 / 247 = 0
    16'b10010110_11111000 : OUT <= 0;  //150 / 248 = 0
    16'b10010110_11111001 : OUT <= 0;  //150 / 249 = 0
    16'b10010110_11111010 : OUT <= 0;  //150 / 250 = 0
    16'b10010110_11111011 : OUT <= 0;  //150 / 251 = 0
    16'b10010110_11111100 : OUT <= 0;  //150 / 252 = 0
    16'b10010110_11111101 : OUT <= 0;  //150 / 253 = 0
    16'b10010110_11111110 : OUT <= 0;  //150 / 254 = 0
    16'b10010110_11111111 : OUT <= 0;  //150 / 255 = 0
    16'b10010111_00000000 : OUT <= 0;  //151 / 0 = 0
    16'b10010111_00000001 : OUT <= 151;  //151 / 1 = 151
    16'b10010111_00000010 : OUT <= 75;  //151 / 2 = 75
    16'b10010111_00000011 : OUT <= 50;  //151 / 3 = 50
    16'b10010111_00000100 : OUT <= 37;  //151 / 4 = 37
    16'b10010111_00000101 : OUT <= 30;  //151 / 5 = 30
    16'b10010111_00000110 : OUT <= 25;  //151 / 6 = 25
    16'b10010111_00000111 : OUT <= 21;  //151 / 7 = 21
    16'b10010111_00001000 : OUT <= 18;  //151 / 8 = 18
    16'b10010111_00001001 : OUT <= 16;  //151 / 9 = 16
    16'b10010111_00001010 : OUT <= 15;  //151 / 10 = 15
    16'b10010111_00001011 : OUT <= 13;  //151 / 11 = 13
    16'b10010111_00001100 : OUT <= 12;  //151 / 12 = 12
    16'b10010111_00001101 : OUT <= 11;  //151 / 13 = 11
    16'b10010111_00001110 : OUT <= 10;  //151 / 14 = 10
    16'b10010111_00001111 : OUT <= 10;  //151 / 15 = 10
    16'b10010111_00010000 : OUT <= 9;  //151 / 16 = 9
    16'b10010111_00010001 : OUT <= 8;  //151 / 17 = 8
    16'b10010111_00010010 : OUT <= 8;  //151 / 18 = 8
    16'b10010111_00010011 : OUT <= 7;  //151 / 19 = 7
    16'b10010111_00010100 : OUT <= 7;  //151 / 20 = 7
    16'b10010111_00010101 : OUT <= 7;  //151 / 21 = 7
    16'b10010111_00010110 : OUT <= 6;  //151 / 22 = 6
    16'b10010111_00010111 : OUT <= 6;  //151 / 23 = 6
    16'b10010111_00011000 : OUT <= 6;  //151 / 24 = 6
    16'b10010111_00011001 : OUT <= 6;  //151 / 25 = 6
    16'b10010111_00011010 : OUT <= 5;  //151 / 26 = 5
    16'b10010111_00011011 : OUT <= 5;  //151 / 27 = 5
    16'b10010111_00011100 : OUT <= 5;  //151 / 28 = 5
    16'b10010111_00011101 : OUT <= 5;  //151 / 29 = 5
    16'b10010111_00011110 : OUT <= 5;  //151 / 30 = 5
    16'b10010111_00011111 : OUT <= 4;  //151 / 31 = 4
    16'b10010111_00100000 : OUT <= 4;  //151 / 32 = 4
    16'b10010111_00100001 : OUT <= 4;  //151 / 33 = 4
    16'b10010111_00100010 : OUT <= 4;  //151 / 34 = 4
    16'b10010111_00100011 : OUT <= 4;  //151 / 35 = 4
    16'b10010111_00100100 : OUT <= 4;  //151 / 36 = 4
    16'b10010111_00100101 : OUT <= 4;  //151 / 37 = 4
    16'b10010111_00100110 : OUT <= 3;  //151 / 38 = 3
    16'b10010111_00100111 : OUT <= 3;  //151 / 39 = 3
    16'b10010111_00101000 : OUT <= 3;  //151 / 40 = 3
    16'b10010111_00101001 : OUT <= 3;  //151 / 41 = 3
    16'b10010111_00101010 : OUT <= 3;  //151 / 42 = 3
    16'b10010111_00101011 : OUT <= 3;  //151 / 43 = 3
    16'b10010111_00101100 : OUT <= 3;  //151 / 44 = 3
    16'b10010111_00101101 : OUT <= 3;  //151 / 45 = 3
    16'b10010111_00101110 : OUT <= 3;  //151 / 46 = 3
    16'b10010111_00101111 : OUT <= 3;  //151 / 47 = 3
    16'b10010111_00110000 : OUT <= 3;  //151 / 48 = 3
    16'b10010111_00110001 : OUT <= 3;  //151 / 49 = 3
    16'b10010111_00110010 : OUT <= 3;  //151 / 50 = 3
    16'b10010111_00110011 : OUT <= 2;  //151 / 51 = 2
    16'b10010111_00110100 : OUT <= 2;  //151 / 52 = 2
    16'b10010111_00110101 : OUT <= 2;  //151 / 53 = 2
    16'b10010111_00110110 : OUT <= 2;  //151 / 54 = 2
    16'b10010111_00110111 : OUT <= 2;  //151 / 55 = 2
    16'b10010111_00111000 : OUT <= 2;  //151 / 56 = 2
    16'b10010111_00111001 : OUT <= 2;  //151 / 57 = 2
    16'b10010111_00111010 : OUT <= 2;  //151 / 58 = 2
    16'b10010111_00111011 : OUT <= 2;  //151 / 59 = 2
    16'b10010111_00111100 : OUT <= 2;  //151 / 60 = 2
    16'b10010111_00111101 : OUT <= 2;  //151 / 61 = 2
    16'b10010111_00111110 : OUT <= 2;  //151 / 62 = 2
    16'b10010111_00111111 : OUT <= 2;  //151 / 63 = 2
    16'b10010111_01000000 : OUT <= 2;  //151 / 64 = 2
    16'b10010111_01000001 : OUT <= 2;  //151 / 65 = 2
    16'b10010111_01000010 : OUT <= 2;  //151 / 66 = 2
    16'b10010111_01000011 : OUT <= 2;  //151 / 67 = 2
    16'b10010111_01000100 : OUT <= 2;  //151 / 68 = 2
    16'b10010111_01000101 : OUT <= 2;  //151 / 69 = 2
    16'b10010111_01000110 : OUT <= 2;  //151 / 70 = 2
    16'b10010111_01000111 : OUT <= 2;  //151 / 71 = 2
    16'b10010111_01001000 : OUT <= 2;  //151 / 72 = 2
    16'b10010111_01001001 : OUT <= 2;  //151 / 73 = 2
    16'b10010111_01001010 : OUT <= 2;  //151 / 74 = 2
    16'b10010111_01001011 : OUT <= 2;  //151 / 75 = 2
    16'b10010111_01001100 : OUT <= 1;  //151 / 76 = 1
    16'b10010111_01001101 : OUT <= 1;  //151 / 77 = 1
    16'b10010111_01001110 : OUT <= 1;  //151 / 78 = 1
    16'b10010111_01001111 : OUT <= 1;  //151 / 79 = 1
    16'b10010111_01010000 : OUT <= 1;  //151 / 80 = 1
    16'b10010111_01010001 : OUT <= 1;  //151 / 81 = 1
    16'b10010111_01010010 : OUT <= 1;  //151 / 82 = 1
    16'b10010111_01010011 : OUT <= 1;  //151 / 83 = 1
    16'b10010111_01010100 : OUT <= 1;  //151 / 84 = 1
    16'b10010111_01010101 : OUT <= 1;  //151 / 85 = 1
    16'b10010111_01010110 : OUT <= 1;  //151 / 86 = 1
    16'b10010111_01010111 : OUT <= 1;  //151 / 87 = 1
    16'b10010111_01011000 : OUT <= 1;  //151 / 88 = 1
    16'b10010111_01011001 : OUT <= 1;  //151 / 89 = 1
    16'b10010111_01011010 : OUT <= 1;  //151 / 90 = 1
    16'b10010111_01011011 : OUT <= 1;  //151 / 91 = 1
    16'b10010111_01011100 : OUT <= 1;  //151 / 92 = 1
    16'b10010111_01011101 : OUT <= 1;  //151 / 93 = 1
    16'b10010111_01011110 : OUT <= 1;  //151 / 94 = 1
    16'b10010111_01011111 : OUT <= 1;  //151 / 95 = 1
    16'b10010111_01100000 : OUT <= 1;  //151 / 96 = 1
    16'b10010111_01100001 : OUT <= 1;  //151 / 97 = 1
    16'b10010111_01100010 : OUT <= 1;  //151 / 98 = 1
    16'b10010111_01100011 : OUT <= 1;  //151 / 99 = 1
    16'b10010111_01100100 : OUT <= 1;  //151 / 100 = 1
    16'b10010111_01100101 : OUT <= 1;  //151 / 101 = 1
    16'b10010111_01100110 : OUT <= 1;  //151 / 102 = 1
    16'b10010111_01100111 : OUT <= 1;  //151 / 103 = 1
    16'b10010111_01101000 : OUT <= 1;  //151 / 104 = 1
    16'b10010111_01101001 : OUT <= 1;  //151 / 105 = 1
    16'b10010111_01101010 : OUT <= 1;  //151 / 106 = 1
    16'b10010111_01101011 : OUT <= 1;  //151 / 107 = 1
    16'b10010111_01101100 : OUT <= 1;  //151 / 108 = 1
    16'b10010111_01101101 : OUT <= 1;  //151 / 109 = 1
    16'b10010111_01101110 : OUT <= 1;  //151 / 110 = 1
    16'b10010111_01101111 : OUT <= 1;  //151 / 111 = 1
    16'b10010111_01110000 : OUT <= 1;  //151 / 112 = 1
    16'b10010111_01110001 : OUT <= 1;  //151 / 113 = 1
    16'b10010111_01110010 : OUT <= 1;  //151 / 114 = 1
    16'b10010111_01110011 : OUT <= 1;  //151 / 115 = 1
    16'b10010111_01110100 : OUT <= 1;  //151 / 116 = 1
    16'b10010111_01110101 : OUT <= 1;  //151 / 117 = 1
    16'b10010111_01110110 : OUT <= 1;  //151 / 118 = 1
    16'b10010111_01110111 : OUT <= 1;  //151 / 119 = 1
    16'b10010111_01111000 : OUT <= 1;  //151 / 120 = 1
    16'b10010111_01111001 : OUT <= 1;  //151 / 121 = 1
    16'b10010111_01111010 : OUT <= 1;  //151 / 122 = 1
    16'b10010111_01111011 : OUT <= 1;  //151 / 123 = 1
    16'b10010111_01111100 : OUT <= 1;  //151 / 124 = 1
    16'b10010111_01111101 : OUT <= 1;  //151 / 125 = 1
    16'b10010111_01111110 : OUT <= 1;  //151 / 126 = 1
    16'b10010111_01111111 : OUT <= 1;  //151 / 127 = 1
    16'b10010111_10000000 : OUT <= 1;  //151 / 128 = 1
    16'b10010111_10000001 : OUT <= 1;  //151 / 129 = 1
    16'b10010111_10000010 : OUT <= 1;  //151 / 130 = 1
    16'b10010111_10000011 : OUT <= 1;  //151 / 131 = 1
    16'b10010111_10000100 : OUT <= 1;  //151 / 132 = 1
    16'b10010111_10000101 : OUT <= 1;  //151 / 133 = 1
    16'b10010111_10000110 : OUT <= 1;  //151 / 134 = 1
    16'b10010111_10000111 : OUT <= 1;  //151 / 135 = 1
    16'b10010111_10001000 : OUT <= 1;  //151 / 136 = 1
    16'b10010111_10001001 : OUT <= 1;  //151 / 137 = 1
    16'b10010111_10001010 : OUT <= 1;  //151 / 138 = 1
    16'b10010111_10001011 : OUT <= 1;  //151 / 139 = 1
    16'b10010111_10001100 : OUT <= 1;  //151 / 140 = 1
    16'b10010111_10001101 : OUT <= 1;  //151 / 141 = 1
    16'b10010111_10001110 : OUT <= 1;  //151 / 142 = 1
    16'b10010111_10001111 : OUT <= 1;  //151 / 143 = 1
    16'b10010111_10010000 : OUT <= 1;  //151 / 144 = 1
    16'b10010111_10010001 : OUT <= 1;  //151 / 145 = 1
    16'b10010111_10010010 : OUT <= 1;  //151 / 146 = 1
    16'b10010111_10010011 : OUT <= 1;  //151 / 147 = 1
    16'b10010111_10010100 : OUT <= 1;  //151 / 148 = 1
    16'b10010111_10010101 : OUT <= 1;  //151 / 149 = 1
    16'b10010111_10010110 : OUT <= 1;  //151 / 150 = 1
    16'b10010111_10010111 : OUT <= 1;  //151 / 151 = 1
    16'b10010111_10011000 : OUT <= 0;  //151 / 152 = 0
    16'b10010111_10011001 : OUT <= 0;  //151 / 153 = 0
    16'b10010111_10011010 : OUT <= 0;  //151 / 154 = 0
    16'b10010111_10011011 : OUT <= 0;  //151 / 155 = 0
    16'b10010111_10011100 : OUT <= 0;  //151 / 156 = 0
    16'b10010111_10011101 : OUT <= 0;  //151 / 157 = 0
    16'b10010111_10011110 : OUT <= 0;  //151 / 158 = 0
    16'b10010111_10011111 : OUT <= 0;  //151 / 159 = 0
    16'b10010111_10100000 : OUT <= 0;  //151 / 160 = 0
    16'b10010111_10100001 : OUT <= 0;  //151 / 161 = 0
    16'b10010111_10100010 : OUT <= 0;  //151 / 162 = 0
    16'b10010111_10100011 : OUT <= 0;  //151 / 163 = 0
    16'b10010111_10100100 : OUT <= 0;  //151 / 164 = 0
    16'b10010111_10100101 : OUT <= 0;  //151 / 165 = 0
    16'b10010111_10100110 : OUT <= 0;  //151 / 166 = 0
    16'b10010111_10100111 : OUT <= 0;  //151 / 167 = 0
    16'b10010111_10101000 : OUT <= 0;  //151 / 168 = 0
    16'b10010111_10101001 : OUT <= 0;  //151 / 169 = 0
    16'b10010111_10101010 : OUT <= 0;  //151 / 170 = 0
    16'b10010111_10101011 : OUT <= 0;  //151 / 171 = 0
    16'b10010111_10101100 : OUT <= 0;  //151 / 172 = 0
    16'b10010111_10101101 : OUT <= 0;  //151 / 173 = 0
    16'b10010111_10101110 : OUT <= 0;  //151 / 174 = 0
    16'b10010111_10101111 : OUT <= 0;  //151 / 175 = 0
    16'b10010111_10110000 : OUT <= 0;  //151 / 176 = 0
    16'b10010111_10110001 : OUT <= 0;  //151 / 177 = 0
    16'b10010111_10110010 : OUT <= 0;  //151 / 178 = 0
    16'b10010111_10110011 : OUT <= 0;  //151 / 179 = 0
    16'b10010111_10110100 : OUT <= 0;  //151 / 180 = 0
    16'b10010111_10110101 : OUT <= 0;  //151 / 181 = 0
    16'b10010111_10110110 : OUT <= 0;  //151 / 182 = 0
    16'b10010111_10110111 : OUT <= 0;  //151 / 183 = 0
    16'b10010111_10111000 : OUT <= 0;  //151 / 184 = 0
    16'b10010111_10111001 : OUT <= 0;  //151 / 185 = 0
    16'b10010111_10111010 : OUT <= 0;  //151 / 186 = 0
    16'b10010111_10111011 : OUT <= 0;  //151 / 187 = 0
    16'b10010111_10111100 : OUT <= 0;  //151 / 188 = 0
    16'b10010111_10111101 : OUT <= 0;  //151 / 189 = 0
    16'b10010111_10111110 : OUT <= 0;  //151 / 190 = 0
    16'b10010111_10111111 : OUT <= 0;  //151 / 191 = 0
    16'b10010111_11000000 : OUT <= 0;  //151 / 192 = 0
    16'b10010111_11000001 : OUT <= 0;  //151 / 193 = 0
    16'b10010111_11000010 : OUT <= 0;  //151 / 194 = 0
    16'b10010111_11000011 : OUT <= 0;  //151 / 195 = 0
    16'b10010111_11000100 : OUT <= 0;  //151 / 196 = 0
    16'b10010111_11000101 : OUT <= 0;  //151 / 197 = 0
    16'b10010111_11000110 : OUT <= 0;  //151 / 198 = 0
    16'b10010111_11000111 : OUT <= 0;  //151 / 199 = 0
    16'b10010111_11001000 : OUT <= 0;  //151 / 200 = 0
    16'b10010111_11001001 : OUT <= 0;  //151 / 201 = 0
    16'b10010111_11001010 : OUT <= 0;  //151 / 202 = 0
    16'b10010111_11001011 : OUT <= 0;  //151 / 203 = 0
    16'b10010111_11001100 : OUT <= 0;  //151 / 204 = 0
    16'b10010111_11001101 : OUT <= 0;  //151 / 205 = 0
    16'b10010111_11001110 : OUT <= 0;  //151 / 206 = 0
    16'b10010111_11001111 : OUT <= 0;  //151 / 207 = 0
    16'b10010111_11010000 : OUT <= 0;  //151 / 208 = 0
    16'b10010111_11010001 : OUT <= 0;  //151 / 209 = 0
    16'b10010111_11010010 : OUT <= 0;  //151 / 210 = 0
    16'b10010111_11010011 : OUT <= 0;  //151 / 211 = 0
    16'b10010111_11010100 : OUT <= 0;  //151 / 212 = 0
    16'b10010111_11010101 : OUT <= 0;  //151 / 213 = 0
    16'b10010111_11010110 : OUT <= 0;  //151 / 214 = 0
    16'b10010111_11010111 : OUT <= 0;  //151 / 215 = 0
    16'b10010111_11011000 : OUT <= 0;  //151 / 216 = 0
    16'b10010111_11011001 : OUT <= 0;  //151 / 217 = 0
    16'b10010111_11011010 : OUT <= 0;  //151 / 218 = 0
    16'b10010111_11011011 : OUT <= 0;  //151 / 219 = 0
    16'b10010111_11011100 : OUT <= 0;  //151 / 220 = 0
    16'b10010111_11011101 : OUT <= 0;  //151 / 221 = 0
    16'b10010111_11011110 : OUT <= 0;  //151 / 222 = 0
    16'b10010111_11011111 : OUT <= 0;  //151 / 223 = 0
    16'b10010111_11100000 : OUT <= 0;  //151 / 224 = 0
    16'b10010111_11100001 : OUT <= 0;  //151 / 225 = 0
    16'b10010111_11100010 : OUT <= 0;  //151 / 226 = 0
    16'b10010111_11100011 : OUT <= 0;  //151 / 227 = 0
    16'b10010111_11100100 : OUT <= 0;  //151 / 228 = 0
    16'b10010111_11100101 : OUT <= 0;  //151 / 229 = 0
    16'b10010111_11100110 : OUT <= 0;  //151 / 230 = 0
    16'b10010111_11100111 : OUT <= 0;  //151 / 231 = 0
    16'b10010111_11101000 : OUT <= 0;  //151 / 232 = 0
    16'b10010111_11101001 : OUT <= 0;  //151 / 233 = 0
    16'b10010111_11101010 : OUT <= 0;  //151 / 234 = 0
    16'b10010111_11101011 : OUT <= 0;  //151 / 235 = 0
    16'b10010111_11101100 : OUT <= 0;  //151 / 236 = 0
    16'b10010111_11101101 : OUT <= 0;  //151 / 237 = 0
    16'b10010111_11101110 : OUT <= 0;  //151 / 238 = 0
    16'b10010111_11101111 : OUT <= 0;  //151 / 239 = 0
    16'b10010111_11110000 : OUT <= 0;  //151 / 240 = 0
    16'b10010111_11110001 : OUT <= 0;  //151 / 241 = 0
    16'b10010111_11110010 : OUT <= 0;  //151 / 242 = 0
    16'b10010111_11110011 : OUT <= 0;  //151 / 243 = 0
    16'b10010111_11110100 : OUT <= 0;  //151 / 244 = 0
    16'b10010111_11110101 : OUT <= 0;  //151 / 245 = 0
    16'b10010111_11110110 : OUT <= 0;  //151 / 246 = 0
    16'b10010111_11110111 : OUT <= 0;  //151 / 247 = 0
    16'b10010111_11111000 : OUT <= 0;  //151 / 248 = 0
    16'b10010111_11111001 : OUT <= 0;  //151 / 249 = 0
    16'b10010111_11111010 : OUT <= 0;  //151 / 250 = 0
    16'b10010111_11111011 : OUT <= 0;  //151 / 251 = 0
    16'b10010111_11111100 : OUT <= 0;  //151 / 252 = 0
    16'b10010111_11111101 : OUT <= 0;  //151 / 253 = 0
    16'b10010111_11111110 : OUT <= 0;  //151 / 254 = 0
    16'b10010111_11111111 : OUT <= 0;  //151 / 255 = 0
    16'b10011000_00000000 : OUT <= 0;  //152 / 0 = 0
    16'b10011000_00000001 : OUT <= 152;  //152 / 1 = 152
    16'b10011000_00000010 : OUT <= 76;  //152 / 2 = 76
    16'b10011000_00000011 : OUT <= 50;  //152 / 3 = 50
    16'b10011000_00000100 : OUT <= 38;  //152 / 4 = 38
    16'b10011000_00000101 : OUT <= 30;  //152 / 5 = 30
    16'b10011000_00000110 : OUT <= 25;  //152 / 6 = 25
    16'b10011000_00000111 : OUT <= 21;  //152 / 7 = 21
    16'b10011000_00001000 : OUT <= 19;  //152 / 8 = 19
    16'b10011000_00001001 : OUT <= 16;  //152 / 9 = 16
    16'b10011000_00001010 : OUT <= 15;  //152 / 10 = 15
    16'b10011000_00001011 : OUT <= 13;  //152 / 11 = 13
    16'b10011000_00001100 : OUT <= 12;  //152 / 12 = 12
    16'b10011000_00001101 : OUT <= 11;  //152 / 13 = 11
    16'b10011000_00001110 : OUT <= 10;  //152 / 14 = 10
    16'b10011000_00001111 : OUT <= 10;  //152 / 15 = 10
    16'b10011000_00010000 : OUT <= 9;  //152 / 16 = 9
    16'b10011000_00010001 : OUT <= 8;  //152 / 17 = 8
    16'b10011000_00010010 : OUT <= 8;  //152 / 18 = 8
    16'b10011000_00010011 : OUT <= 8;  //152 / 19 = 8
    16'b10011000_00010100 : OUT <= 7;  //152 / 20 = 7
    16'b10011000_00010101 : OUT <= 7;  //152 / 21 = 7
    16'b10011000_00010110 : OUT <= 6;  //152 / 22 = 6
    16'b10011000_00010111 : OUT <= 6;  //152 / 23 = 6
    16'b10011000_00011000 : OUT <= 6;  //152 / 24 = 6
    16'b10011000_00011001 : OUT <= 6;  //152 / 25 = 6
    16'b10011000_00011010 : OUT <= 5;  //152 / 26 = 5
    16'b10011000_00011011 : OUT <= 5;  //152 / 27 = 5
    16'b10011000_00011100 : OUT <= 5;  //152 / 28 = 5
    16'b10011000_00011101 : OUT <= 5;  //152 / 29 = 5
    16'b10011000_00011110 : OUT <= 5;  //152 / 30 = 5
    16'b10011000_00011111 : OUT <= 4;  //152 / 31 = 4
    16'b10011000_00100000 : OUT <= 4;  //152 / 32 = 4
    16'b10011000_00100001 : OUT <= 4;  //152 / 33 = 4
    16'b10011000_00100010 : OUT <= 4;  //152 / 34 = 4
    16'b10011000_00100011 : OUT <= 4;  //152 / 35 = 4
    16'b10011000_00100100 : OUT <= 4;  //152 / 36 = 4
    16'b10011000_00100101 : OUT <= 4;  //152 / 37 = 4
    16'b10011000_00100110 : OUT <= 4;  //152 / 38 = 4
    16'b10011000_00100111 : OUT <= 3;  //152 / 39 = 3
    16'b10011000_00101000 : OUT <= 3;  //152 / 40 = 3
    16'b10011000_00101001 : OUT <= 3;  //152 / 41 = 3
    16'b10011000_00101010 : OUT <= 3;  //152 / 42 = 3
    16'b10011000_00101011 : OUT <= 3;  //152 / 43 = 3
    16'b10011000_00101100 : OUT <= 3;  //152 / 44 = 3
    16'b10011000_00101101 : OUT <= 3;  //152 / 45 = 3
    16'b10011000_00101110 : OUT <= 3;  //152 / 46 = 3
    16'b10011000_00101111 : OUT <= 3;  //152 / 47 = 3
    16'b10011000_00110000 : OUT <= 3;  //152 / 48 = 3
    16'b10011000_00110001 : OUT <= 3;  //152 / 49 = 3
    16'b10011000_00110010 : OUT <= 3;  //152 / 50 = 3
    16'b10011000_00110011 : OUT <= 2;  //152 / 51 = 2
    16'b10011000_00110100 : OUT <= 2;  //152 / 52 = 2
    16'b10011000_00110101 : OUT <= 2;  //152 / 53 = 2
    16'b10011000_00110110 : OUT <= 2;  //152 / 54 = 2
    16'b10011000_00110111 : OUT <= 2;  //152 / 55 = 2
    16'b10011000_00111000 : OUT <= 2;  //152 / 56 = 2
    16'b10011000_00111001 : OUT <= 2;  //152 / 57 = 2
    16'b10011000_00111010 : OUT <= 2;  //152 / 58 = 2
    16'b10011000_00111011 : OUT <= 2;  //152 / 59 = 2
    16'b10011000_00111100 : OUT <= 2;  //152 / 60 = 2
    16'b10011000_00111101 : OUT <= 2;  //152 / 61 = 2
    16'b10011000_00111110 : OUT <= 2;  //152 / 62 = 2
    16'b10011000_00111111 : OUT <= 2;  //152 / 63 = 2
    16'b10011000_01000000 : OUT <= 2;  //152 / 64 = 2
    16'b10011000_01000001 : OUT <= 2;  //152 / 65 = 2
    16'b10011000_01000010 : OUT <= 2;  //152 / 66 = 2
    16'b10011000_01000011 : OUT <= 2;  //152 / 67 = 2
    16'b10011000_01000100 : OUT <= 2;  //152 / 68 = 2
    16'b10011000_01000101 : OUT <= 2;  //152 / 69 = 2
    16'b10011000_01000110 : OUT <= 2;  //152 / 70 = 2
    16'b10011000_01000111 : OUT <= 2;  //152 / 71 = 2
    16'b10011000_01001000 : OUT <= 2;  //152 / 72 = 2
    16'b10011000_01001001 : OUT <= 2;  //152 / 73 = 2
    16'b10011000_01001010 : OUT <= 2;  //152 / 74 = 2
    16'b10011000_01001011 : OUT <= 2;  //152 / 75 = 2
    16'b10011000_01001100 : OUT <= 2;  //152 / 76 = 2
    16'b10011000_01001101 : OUT <= 1;  //152 / 77 = 1
    16'b10011000_01001110 : OUT <= 1;  //152 / 78 = 1
    16'b10011000_01001111 : OUT <= 1;  //152 / 79 = 1
    16'b10011000_01010000 : OUT <= 1;  //152 / 80 = 1
    16'b10011000_01010001 : OUT <= 1;  //152 / 81 = 1
    16'b10011000_01010010 : OUT <= 1;  //152 / 82 = 1
    16'b10011000_01010011 : OUT <= 1;  //152 / 83 = 1
    16'b10011000_01010100 : OUT <= 1;  //152 / 84 = 1
    16'b10011000_01010101 : OUT <= 1;  //152 / 85 = 1
    16'b10011000_01010110 : OUT <= 1;  //152 / 86 = 1
    16'b10011000_01010111 : OUT <= 1;  //152 / 87 = 1
    16'b10011000_01011000 : OUT <= 1;  //152 / 88 = 1
    16'b10011000_01011001 : OUT <= 1;  //152 / 89 = 1
    16'b10011000_01011010 : OUT <= 1;  //152 / 90 = 1
    16'b10011000_01011011 : OUT <= 1;  //152 / 91 = 1
    16'b10011000_01011100 : OUT <= 1;  //152 / 92 = 1
    16'b10011000_01011101 : OUT <= 1;  //152 / 93 = 1
    16'b10011000_01011110 : OUT <= 1;  //152 / 94 = 1
    16'b10011000_01011111 : OUT <= 1;  //152 / 95 = 1
    16'b10011000_01100000 : OUT <= 1;  //152 / 96 = 1
    16'b10011000_01100001 : OUT <= 1;  //152 / 97 = 1
    16'b10011000_01100010 : OUT <= 1;  //152 / 98 = 1
    16'b10011000_01100011 : OUT <= 1;  //152 / 99 = 1
    16'b10011000_01100100 : OUT <= 1;  //152 / 100 = 1
    16'b10011000_01100101 : OUT <= 1;  //152 / 101 = 1
    16'b10011000_01100110 : OUT <= 1;  //152 / 102 = 1
    16'b10011000_01100111 : OUT <= 1;  //152 / 103 = 1
    16'b10011000_01101000 : OUT <= 1;  //152 / 104 = 1
    16'b10011000_01101001 : OUT <= 1;  //152 / 105 = 1
    16'b10011000_01101010 : OUT <= 1;  //152 / 106 = 1
    16'b10011000_01101011 : OUT <= 1;  //152 / 107 = 1
    16'b10011000_01101100 : OUT <= 1;  //152 / 108 = 1
    16'b10011000_01101101 : OUT <= 1;  //152 / 109 = 1
    16'b10011000_01101110 : OUT <= 1;  //152 / 110 = 1
    16'b10011000_01101111 : OUT <= 1;  //152 / 111 = 1
    16'b10011000_01110000 : OUT <= 1;  //152 / 112 = 1
    16'b10011000_01110001 : OUT <= 1;  //152 / 113 = 1
    16'b10011000_01110010 : OUT <= 1;  //152 / 114 = 1
    16'b10011000_01110011 : OUT <= 1;  //152 / 115 = 1
    16'b10011000_01110100 : OUT <= 1;  //152 / 116 = 1
    16'b10011000_01110101 : OUT <= 1;  //152 / 117 = 1
    16'b10011000_01110110 : OUT <= 1;  //152 / 118 = 1
    16'b10011000_01110111 : OUT <= 1;  //152 / 119 = 1
    16'b10011000_01111000 : OUT <= 1;  //152 / 120 = 1
    16'b10011000_01111001 : OUT <= 1;  //152 / 121 = 1
    16'b10011000_01111010 : OUT <= 1;  //152 / 122 = 1
    16'b10011000_01111011 : OUT <= 1;  //152 / 123 = 1
    16'b10011000_01111100 : OUT <= 1;  //152 / 124 = 1
    16'b10011000_01111101 : OUT <= 1;  //152 / 125 = 1
    16'b10011000_01111110 : OUT <= 1;  //152 / 126 = 1
    16'b10011000_01111111 : OUT <= 1;  //152 / 127 = 1
    16'b10011000_10000000 : OUT <= 1;  //152 / 128 = 1
    16'b10011000_10000001 : OUT <= 1;  //152 / 129 = 1
    16'b10011000_10000010 : OUT <= 1;  //152 / 130 = 1
    16'b10011000_10000011 : OUT <= 1;  //152 / 131 = 1
    16'b10011000_10000100 : OUT <= 1;  //152 / 132 = 1
    16'b10011000_10000101 : OUT <= 1;  //152 / 133 = 1
    16'b10011000_10000110 : OUT <= 1;  //152 / 134 = 1
    16'b10011000_10000111 : OUT <= 1;  //152 / 135 = 1
    16'b10011000_10001000 : OUT <= 1;  //152 / 136 = 1
    16'b10011000_10001001 : OUT <= 1;  //152 / 137 = 1
    16'b10011000_10001010 : OUT <= 1;  //152 / 138 = 1
    16'b10011000_10001011 : OUT <= 1;  //152 / 139 = 1
    16'b10011000_10001100 : OUT <= 1;  //152 / 140 = 1
    16'b10011000_10001101 : OUT <= 1;  //152 / 141 = 1
    16'b10011000_10001110 : OUT <= 1;  //152 / 142 = 1
    16'b10011000_10001111 : OUT <= 1;  //152 / 143 = 1
    16'b10011000_10010000 : OUT <= 1;  //152 / 144 = 1
    16'b10011000_10010001 : OUT <= 1;  //152 / 145 = 1
    16'b10011000_10010010 : OUT <= 1;  //152 / 146 = 1
    16'b10011000_10010011 : OUT <= 1;  //152 / 147 = 1
    16'b10011000_10010100 : OUT <= 1;  //152 / 148 = 1
    16'b10011000_10010101 : OUT <= 1;  //152 / 149 = 1
    16'b10011000_10010110 : OUT <= 1;  //152 / 150 = 1
    16'b10011000_10010111 : OUT <= 1;  //152 / 151 = 1
    16'b10011000_10011000 : OUT <= 1;  //152 / 152 = 1
    16'b10011000_10011001 : OUT <= 0;  //152 / 153 = 0
    16'b10011000_10011010 : OUT <= 0;  //152 / 154 = 0
    16'b10011000_10011011 : OUT <= 0;  //152 / 155 = 0
    16'b10011000_10011100 : OUT <= 0;  //152 / 156 = 0
    16'b10011000_10011101 : OUT <= 0;  //152 / 157 = 0
    16'b10011000_10011110 : OUT <= 0;  //152 / 158 = 0
    16'b10011000_10011111 : OUT <= 0;  //152 / 159 = 0
    16'b10011000_10100000 : OUT <= 0;  //152 / 160 = 0
    16'b10011000_10100001 : OUT <= 0;  //152 / 161 = 0
    16'b10011000_10100010 : OUT <= 0;  //152 / 162 = 0
    16'b10011000_10100011 : OUT <= 0;  //152 / 163 = 0
    16'b10011000_10100100 : OUT <= 0;  //152 / 164 = 0
    16'b10011000_10100101 : OUT <= 0;  //152 / 165 = 0
    16'b10011000_10100110 : OUT <= 0;  //152 / 166 = 0
    16'b10011000_10100111 : OUT <= 0;  //152 / 167 = 0
    16'b10011000_10101000 : OUT <= 0;  //152 / 168 = 0
    16'b10011000_10101001 : OUT <= 0;  //152 / 169 = 0
    16'b10011000_10101010 : OUT <= 0;  //152 / 170 = 0
    16'b10011000_10101011 : OUT <= 0;  //152 / 171 = 0
    16'b10011000_10101100 : OUT <= 0;  //152 / 172 = 0
    16'b10011000_10101101 : OUT <= 0;  //152 / 173 = 0
    16'b10011000_10101110 : OUT <= 0;  //152 / 174 = 0
    16'b10011000_10101111 : OUT <= 0;  //152 / 175 = 0
    16'b10011000_10110000 : OUT <= 0;  //152 / 176 = 0
    16'b10011000_10110001 : OUT <= 0;  //152 / 177 = 0
    16'b10011000_10110010 : OUT <= 0;  //152 / 178 = 0
    16'b10011000_10110011 : OUT <= 0;  //152 / 179 = 0
    16'b10011000_10110100 : OUT <= 0;  //152 / 180 = 0
    16'b10011000_10110101 : OUT <= 0;  //152 / 181 = 0
    16'b10011000_10110110 : OUT <= 0;  //152 / 182 = 0
    16'b10011000_10110111 : OUT <= 0;  //152 / 183 = 0
    16'b10011000_10111000 : OUT <= 0;  //152 / 184 = 0
    16'b10011000_10111001 : OUT <= 0;  //152 / 185 = 0
    16'b10011000_10111010 : OUT <= 0;  //152 / 186 = 0
    16'b10011000_10111011 : OUT <= 0;  //152 / 187 = 0
    16'b10011000_10111100 : OUT <= 0;  //152 / 188 = 0
    16'b10011000_10111101 : OUT <= 0;  //152 / 189 = 0
    16'b10011000_10111110 : OUT <= 0;  //152 / 190 = 0
    16'b10011000_10111111 : OUT <= 0;  //152 / 191 = 0
    16'b10011000_11000000 : OUT <= 0;  //152 / 192 = 0
    16'b10011000_11000001 : OUT <= 0;  //152 / 193 = 0
    16'b10011000_11000010 : OUT <= 0;  //152 / 194 = 0
    16'b10011000_11000011 : OUT <= 0;  //152 / 195 = 0
    16'b10011000_11000100 : OUT <= 0;  //152 / 196 = 0
    16'b10011000_11000101 : OUT <= 0;  //152 / 197 = 0
    16'b10011000_11000110 : OUT <= 0;  //152 / 198 = 0
    16'b10011000_11000111 : OUT <= 0;  //152 / 199 = 0
    16'b10011000_11001000 : OUT <= 0;  //152 / 200 = 0
    16'b10011000_11001001 : OUT <= 0;  //152 / 201 = 0
    16'b10011000_11001010 : OUT <= 0;  //152 / 202 = 0
    16'b10011000_11001011 : OUT <= 0;  //152 / 203 = 0
    16'b10011000_11001100 : OUT <= 0;  //152 / 204 = 0
    16'b10011000_11001101 : OUT <= 0;  //152 / 205 = 0
    16'b10011000_11001110 : OUT <= 0;  //152 / 206 = 0
    16'b10011000_11001111 : OUT <= 0;  //152 / 207 = 0
    16'b10011000_11010000 : OUT <= 0;  //152 / 208 = 0
    16'b10011000_11010001 : OUT <= 0;  //152 / 209 = 0
    16'b10011000_11010010 : OUT <= 0;  //152 / 210 = 0
    16'b10011000_11010011 : OUT <= 0;  //152 / 211 = 0
    16'b10011000_11010100 : OUT <= 0;  //152 / 212 = 0
    16'b10011000_11010101 : OUT <= 0;  //152 / 213 = 0
    16'b10011000_11010110 : OUT <= 0;  //152 / 214 = 0
    16'b10011000_11010111 : OUT <= 0;  //152 / 215 = 0
    16'b10011000_11011000 : OUT <= 0;  //152 / 216 = 0
    16'b10011000_11011001 : OUT <= 0;  //152 / 217 = 0
    16'b10011000_11011010 : OUT <= 0;  //152 / 218 = 0
    16'b10011000_11011011 : OUT <= 0;  //152 / 219 = 0
    16'b10011000_11011100 : OUT <= 0;  //152 / 220 = 0
    16'b10011000_11011101 : OUT <= 0;  //152 / 221 = 0
    16'b10011000_11011110 : OUT <= 0;  //152 / 222 = 0
    16'b10011000_11011111 : OUT <= 0;  //152 / 223 = 0
    16'b10011000_11100000 : OUT <= 0;  //152 / 224 = 0
    16'b10011000_11100001 : OUT <= 0;  //152 / 225 = 0
    16'b10011000_11100010 : OUT <= 0;  //152 / 226 = 0
    16'b10011000_11100011 : OUT <= 0;  //152 / 227 = 0
    16'b10011000_11100100 : OUT <= 0;  //152 / 228 = 0
    16'b10011000_11100101 : OUT <= 0;  //152 / 229 = 0
    16'b10011000_11100110 : OUT <= 0;  //152 / 230 = 0
    16'b10011000_11100111 : OUT <= 0;  //152 / 231 = 0
    16'b10011000_11101000 : OUT <= 0;  //152 / 232 = 0
    16'b10011000_11101001 : OUT <= 0;  //152 / 233 = 0
    16'b10011000_11101010 : OUT <= 0;  //152 / 234 = 0
    16'b10011000_11101011 : OUT <= 0;  //152 / 235 = 0
    16'b10011000_11101100 : OUT <= 0;  //152 / 236 = 0
    16'b10011000_11101101 : OUT <= 0;  //152 / 237 = 0
    16'b10011000_11101110 : OUT <= 0;  //152 / 238 = 0
    16'b10011000_11101111 : OUT <= 0;  //152 / 239 = 0
    16'b10011000_11110000 : OUT <= 0;  //152 / 240 = 0
    16'b10011000_11110001 : OUT <= 0;  //152 / 241 = 0
    16'b10011000_11110010 : OUT <= 0;  //152 / 242 = 0
    16'b10011000_11110011 : OUT <= 0;  //152 / 243 = 0
    16'b10011000_11110100 : OUT <= 0;  //152 / 244 = 0
    16'b10011000_11110101 : OUT <= 0;  //152 / 245 = 0
    16'b10011000_11110110 : OUT <= 0;  //152 / 246 = 0
    16'b10011000_11110111 : OUT <= 0;  //152 / 247 = 0
    16'b10011000_11111000 : OUT <= 0;  //152 / 248 = 0
    16'b10011000_11111001 : OUT <= 0;  //152 / 249 = 0
    16'b10011000_11111010 : OUT <= 0;  //152 / 250 = 0
    16'b10011000_11111011 : OUT <= 0;  //152 / 251 = 0
    16'b10011000_11111100 : OUT <= 0;  //152 / 252 = 0
    16'b10011000_11111101 : OUT <= 0;  //152 / 253 = 0
    16'b10011000_11111110 : OUT <= 0;  //152 / 254 = 0
    16'b10011000_11111111 : OUT <= 0;  //152 / 255 = 0
    16'b10011001_00000000 : OUT <= 0;  //153 / 0 = 0
    16'b10011001_00000001 : OUT <= 153;  //153 / 1 = 153
    16'b10011001_00000010 : OUT <= 76;  //153 / 2 = 76
    16'b10011001_00000011 : OUT <= 51;  //153 / 3 = 51
    16'b10011001_00000100 : OUT <= 38;  //153 / 4 = 38
    16'b10011001_00000101 : OUT <= 30;  //153 / 5 = 30
    16'b10011001_00000110 : OUT <= 25;  //153 / 6 = 25
    16'b10011001_00000111 : OUT <= 21;  //153 / 7 = 21
    16'b10011001_00001000 : OUT <= 19;  //153 / 8 = 19
    16'b10011001_00001001 : OUT <= 17;  //153 / 9 = 17
    16'b10011001_00001010 : OUT <= 15;  //153 / 10 = 15
    16'b10011001_00001011 : OUT <= 13;  //153 / 11 = 13
    16'b10011001_00001100 : OUT <= 12;  //153 / 12 = 12
    16'b10011001_00001101 : OUT <= 11;  //153 / 13 = 11
    16'b10011001_00001110 : OUT <= 10;  //153 / 14 = 10
    16'b10011001_00001111 : OUT <= 10;  //153 / 15 = 10
    16'b10011001_00010000 : OUT <= 9;  //153 / 16 = 9
    16'b10011001_00010001 : OUT <= 9;  //153 / 17 = 9
    16'b10011001_00010010 : OUT <= 8;  //153 / 18 = 8
    16'b10011001_00010011 : OUT <= 8;  //153 / 19 = 8
    16'b10011001_00010100 : OUT <= 7;  //153 / 20 = 7
    16'b10011001_00010101 : OUT <= 7;  //153 / 21 = 7
    16'b10011001_00010110 : OUT <= 6;  //153 / 22 = 6
    16'b10011001_00010111 : OUT <= 6;  //153 / 23 = 6
    16'b10011001_00011000 : OUT <= 6;  //153 / 24 = 6
    16'b10011001_00011001 : OUT <= 6;  //153 / 25 = 6
    16'b10011001_00011010 : OUT <= 5;  //153 / 26 = 5
    16'b10011001_00011011 : OUT <= 5;  //153 / 27 = 5
    16'b10011001_00011100 : OUT <= 5;  //153 / 28 = 5
    16'b10011001_00011101 : OUT <= 5;  //153 / 29 = 5
    16'b10011001_00011110 : OUT <= 5;  //153 / 30 = 5
    16'b10011001_00011111 : OUT <= 4;  //153 / 31 = 4
    16'b10011001_00100000 : OUT <= 4;  //153 / 32 = 4
    16'b10011001_00100001 : OUT <= 4;  //153 / 33 = 4
    16'b10011001_00100010 : OUT <= 4;  //153 / 34 = 4
    16'b10011001_00100011 : OUT <= 4;  //153 / 35 = 4
    16'b10011001_00100100 : OUT <= 4;  //153 / 36 = 4
    16'b10011001_00100101 : OUT <= 4;  //153 / 37 = 4
    16'b10011001_00100110 : OUT <= 4;  //153 / 38 = 4
    16'b10011001_00100111 : OUT <= 3;  //153 / 39 = 3
    16'b10011001_00101000 : OUT <= 3;  //153 / 40 = 3
    16'b10011001_00101001 : OUT <= 3;  //153 / 41 = 3
    16'b10011001_00101010 : OUT <= 3;  //153 / 42 = 3
    16'b10011001_00101011 : OUT <= 3;  //153 / 43 = 3
    16'b10011001_00101100 : OUT <= 3;  //153 / 44 = 3
    16'b10011001_00101101 : OUT <= 3;  //153 / 45 = 3
    16'b10011001_00101110 : OUT <= 3;  //153 / 46 = 3
    16'b10011001_00101111 : OUT <= 3;  //153 / 47 = 3
    16'b10011001_00110000 : OUT <= 3;  //153 / 48 = 3
    16'b10011001_00110001 : OUT <= 3;  //153 / 49 = 3
    16'b10011001_00110010 : OUT <= 3;  //153 / 50 = 3
    16'b10011001_00110011 : OUT <= 3;  //153 / 51 = 3
    16'b10011001_00110100 : OUT <= 2;  //153 / 52 = 2
    16'b10011001_00110101 : OUT <= 2;  //153 / 53 = 2
    16'b10011001_00110110 : OUT <= 2;  //153 / 54 = 2
    16'b10011001_00110111 : OUT <= 2;  //153 / 55 = 2
    16'b10011001_00111000 : OUT <= 2;  //153 / 56 = 2
    16'b10011001_00111001 : OUT <= 2;  //153 / 57 = 2
    16'b10011001_00111010 : OUT <= 2;  //153 / 58 = 2
    16'b10011001_00111011 : OUT <= 2;  //153 / 59 = 2
    16'b10011001_00111100 : OUT <= 2;  //153 / 60 = 2
    16'b10011001_00111101 : OUT <= 2;  //153 / 61 = 2
    16'b10011001_00111110 : OUT <= 2;  //153 / 62 = 2
    16'b10011001_00111111 : OUT <= 2;  //153 / 63 = 2
    16'b10011001_01000000 : OUT <= 2;  //153 / 64 = 2
    16'b10011001_01000001 : OUT <= 2;  //153 / 65 = 2
    16'b10011001_01000010 : OUT <= 2;  //153 / 66 = 2
    16'b10011001_01000011 : OUT <= 2;  //153 / 67 = 2
    16'b10011001_01000100 : OUT <= 2;  //153 / 68 = 2
    16'b10011001_01000101 : OUT <= 2;  //153 / 69 = 2
    16'b10011001_01000110 : OUT <= 2;  //153 / 70 = 2
    16'b10011001_01000111 : OUT <= 2;  //153 / 71 = 2
    16'b10011001_01001000 : OUT <= 2;  //153 / 72 = 2
    16'b10011001_01001001 : OUT <= 2;  //153 / 73 = 2
    16'b10011001_01001010 : OUT <= 2;  //153 / 74 = 2
    16'b10011001_01001011 : OUT <= 2;  //153 / 75 = 2
    16'b10011001_01001100 : OUT <= 2;  //153 / 76 = 2
    16'b10011001_01001101 : OUT <= 1;  //153 / 77 = 1
    16'b10011001_01001110 : OUT <= 1;  //153 / 78 = 1
    16'b10011001_01001111 : OUT <= 1;  //153 / 79 = 1
    16'b10011001_01010000 : OUT <= 1;  //153 / 80 = 1
    16'b10011001_01010001 : OUT <= 1;  //153 / 81 = 1
    16'b10011001_01010010 : OUT <= 1;  //153 / 82 = 1
    16'b10011001_01010011 : OUT <= 1;  //153 / 83 = 1
    16'b10011001_01010100 : OUT <= 1;  //153 / 84 = 1
    16'b10011001_01010101 : OUT <= 1;  //153 / 85 = 1
    16'b10011001_01010110 : OUT <= 1;  //153 / 86 = 1
    16'b10011001_01010111 : OUT <= 1;  //153 / 87 = 1
    16'b10011001_01011000 : OUT <= 1;  //153 / 88 = 1
    16'b10011001_01011001 : OUT <= 1;  //153 / 89 = 1
    16'b10011001_01011010 : OUT <= 1;  //153 / 90 = 1
    16'b10011001_01011011 : OUT <= 1;  //153 / 91 = 1
    16'b10011001_01011100 : OUT <= 1;  //153 / 92 = 1
    16'b10011001_01011101 : OUT <= 1;  //153 / 93 = 1
    16'b10011001_01011110 : OUT <= 1;  //153 / 94 = 1
    16'b10011001_01011111 : OUT <= 1;  //153 / 95 = 1
    16'b10011001_01100000 : OUT <= 1;  //153 / 96 = 1
    16'b10011001_01100001 : OUT <= 1;  //153 / 97 = 1
    16'b10011001_01100010 : OUT <= 1;  //153 / 98 = 1
    16'b10011001_01100011 : OUT <= 1;  //153 / 99 = 1
    16'b10011001_01100100 : OUT <= 1;  //153 / 100 = 1
    16'b10011001_01100101 : OUT <= 1;  //153 / 101 = 1
    16'b10011001_01100110 : OUT <= 1;  //153 / 102 = 1
    16'b10011001_01100111 : OUT <= 1;  //153 / 103 = 1
    16'b10011001_01101000 : OUT <= 1;  //153 / 104 = 1
    16'b10011001_01101001 : OUT <= 1;  //153 / 105 = 1
    16'b10011001_01101010 : OUT <= 1;  //153 / 106 = 1
    16'b10011001_01101011 : OUT <= 1;  //153 / 107 = 1
    16'b10011001_01101100 : OUT <= 1;  //153 / 108 = 1
    16'b10011001_01101101 : OUT <= 1;  //153 / 109 = 1
    16'b10011001_01101110 : OUT <= 1;  //153 / 110 = 1
    16'b10011001_01101111 : OUT <= 1;  //153 / 111 = 1
    16'b10011001_01110000 : OUT <= 1;  //153 / 112 = 1
    16'b10011001_01110001 : OUT <= 1;  //153 / 113 = 1
    16'b10011001_01110010 : OUT <= 1;  //153 / 114 = 1
    16'b10011001_01110011 : OUT <= 1;  //153 / 115 = 1
    16'b10011001_01110100 : OUT <= 1;  //153 / 116 = 1
    16'b10011001_01110101 : OUT <= 1;  //153 / 117 = 1
    16'b10011001_01110110 : OUT <= 1;  //153 / 118 = 1
    16'b10011001_01110111 : OUT <= 1;  //153 / 119 = 1
    16'b10011001_01111000 : OUT <= 1;  //153 / 120 = 1
    16'b10011001_01111001 : OUT <= 1;  //153 / 121 = 1
    16'b10011001_01111010 : OUT <= 1;  //153 / 122 = 1
    16'b10011001_01111011 : OUT <= 1;  //153 / 123 = 1
    16'b10011001_01111100 : OUT <= 1;  //153 / 124 = 1
    16'b10011001_01111101 : OUT <= 1;  //153 / 125 = 1
    16'b10011001_01111110 : OUT <= 1;  //153 / 126 = 1
    16'b10011001_01111111 : OUT <= 1;  //153 / 127 = 1
    16'b10011001_10000000 : OUT <= 1;  //153 / 128 = 1
    16'b10011001_10000001 : OUT <= 1;  //153 / 129 = 1
    16'b10011001_10000010 : OUT <= 1;  //153 / 130 = 1
    16'b10011001_10000011 : OUT <= 1;  //153 / 131 = 1
    16'b10011001_10000100 : OUT <= 1;  //153 / 132 = 1
    16'b10011001_10000101 : OUT <= 1;  //153 / 133 = 1
    16'b10011001_10000110 : OUT <= 1;  //153 / 134 = 1
    16'b10011001_10000111 : OUT <= 1;  //153 / 135 = 1
    16'b10011001_10001000 : OUT <= 1;  //153 / 136 = 1
    16'b10011001_10001001 : OUT <= 1;  //153 / 137 = 1
    16'b10011001_10001010 : OUT <= 1;  //153 / 138 = 1
    16'b10011001_10001011 : OUT <= 1;  //153 / 139 = 1
    16'b10011001_10001100 : OUT <= 1;  //153 / 140 = 1
    16'b10011001_10001101 : OUT <= 1;  //153 / 141 = 1
    16'b10011001_10001110 : OUT <= 1;  //153 / 142 = 1
    16'b10011001_10001111 : OUT <= 1;  //153 / 143 = 1
    16'b10011001_10010000 : OUT <= 1;  //153 / 144 = 1
    16'b10011001_10010001 : OUT <= 1;  //153 / 145 = 1
    16'b10011001_10010010 : OUT <= 1;  //153 / 146 = 1
    16'b10011001_10010011 : OUT <= 1;  //153 / 147 = 1
    16'b10011001_10010100 : OUT <= 1;  //153 / 148 = 1
    16'b10011001_10010101 : OUT <= 1;  //153 / 149 = 1
    16'b10011001_10010110 : OUT <= 1;  //153 / 150 = 1
    16'b10011001_10010111 : OUT <= 1;  //153 / 151 = 1
    16'b10011001_10011000 : OUT <= 1;  //153 / 152 = 1
    16'b10011001_10011001 : OUT <= 1;  //153 / 153 = 1
    16'b10011001_10011010 : OUT <= 0;  //153 / 154 = 0
    16'b10011001_10011011 : OUT <= 0;  //153 / 155 = 0
    16'b10011001_10011100 : OUT <= 0;  //153 / 156 = 0
    16'b10011001_10011101 : OUT <= 0;  //153 / 157 = 0
    16'b10011001_10011110 : OUT <= 0;  //153 / 158 = 0
    16'b10011001_10011111 : OUT <= 0;  //153 / 159 = 0
    16'b10011001_10100000 : OUT <= 0;  //153 / 160 = 0
    16'b10011001_10100001 : OUT <= 0;  //153 / 161 = 0
    16'b10011001_10100010 : OUT <= 0;  //153 / 162 = 0
    16'b10011001_10100011 : OUT <= 0;  //153 / 163 = 0
    16'b10011001_10100100 : OUT <= 0;  //153 / 164 = 0
    16'b10011001_10100101 : OUT <= 0;  //153 / 165 = 0
    16'b10011001_10100110 : OUT <= 0;  //153 / 166 = 0
    16'b10011001_10100111 : OUT <= 0;  //153 / 167 = 0
    16'b10011001_10101000 : OUT <= 0;  //153 / 168 = 0
    16'b10011001_10101001 : OUT <= 0;  //153 / 169 = 0
    16'b10011001_10101010 : OUT <= 0;  //153 / 170 = 0
    16'b10011001_10101011 : OUT <= 0;  //153 / 171 = 0
    16'b10011001_10101100 : OUT <= 0;  //153 / 172 = 0
    16'b10011001_10101101 : OUT <= 0;  //153 / 173 = 0
    16'b10011001_10101110 : OUT <= 0;  //153 / 174 = 0
    16'b10011001_10101111 : OUT <= 0;  //153 / 175 = 0
    16'b10011001_10110000 : OUT <= 0;  //153 / 176 = 0
    16'b10011001_10110001 : OUT <= 0;  //153 / 177 = 0
    16'b10011001_10110010 : OUT <= 0;  //153 / 178 = 0
    16'b10011001_10110011 : OUT <= 0;  //153 / 179 = 0
    16'b10011001_10110100 : OUT <= 0;  //153 / 180 = 0
    16'b10011001_10110101 : OUT <= 0;  //153 / 181 = 0
    16'b10011001_10110110 : OUT <= 0;  //153 / 182 = 0
    16'b10011001_10110111 : OUT <= 0;  //153 / 183 = 0
    16'b10011001_10111000 : OUT <= 0;  //153 / 184 = 0
    16'b10011001_10111001 : OUT <= 0;  //153 / 185 = 0
    16'b10011001_10111010 : OUT <= 0;  //153 / 186 = 0
    16'b10011001_10111011 : OUT <= 0;  //153 / 187 = 0
    16'b10011001_10111100 : OUT <= 0;  //153 / 188 = 0
    16'b10011001_10111101 : OUT <= 0;  //153 / 189 = 0
    16'b10011001_10111110 : OUT <= 0;  //153 / 190 = 0
    16'b10011001_10111111 : OUT <= 0;  //153 / 191 = 0
    16'b10011001_11000000 : OUT <= 0;  //153 / 192 = 0
    16'b10011001_11000001 : OUT <= 0;  //153 / 193 = 0
    16'b10011001_11000010 : OUT <= 0;  //153 / 194 = 0
    16'b10011001_11000011 : OUT <= 0;  //153 / 195 = 0
    16'b10011001_11000100 : OUT <= 0;  //153 / 196 = 0
    16'b10011001_11000101 : OUT <= 0;  //153 / 197 = 0
    16'b10011001_11000110 : OUT <= 0;  //153 / 198 = 0
    16'b10011001_11000111 : OUT <= 0;  //153 / 199 = 0
    16'b10011001_11001000 : OUT <= 0;  //153 / 200 = 0
    16'b10011001_11001001 : OUT <= 0;  //153 / 201 = 0
    16'b10011001_11001010 : OUT <= 0;  //153 / 202 = 0
    16'b10011001_11001011 : OUT <= 0;  //153 / 203 = 0
    16'b10011001_11001100 : OUT <= 0;  //153 / 204 = 0
    16'b10011001_11001101 : OUT <= 0;  //153 / 205 = 0
    16'b10011001_11001110 : OUT <= 0;  //153 / 206 = 0
    16'b10011001_11001111 : OUT <= 0;  //153 / 207 = 0
    16'b10011001_11010000 : OUT <= 0;  //153 / 208 = 0
    16'b10011001_11010001 : OUT <= 0;  //153 / 209 = 0
    16'b10011001_11010010 : OUT <= 0;  //153 / 210 = 0
    16'b10011001_11010011 : OUT <= 0;  //153 / 211 = 0
    16'b10011001_11010100 : OUT <= 0;  //153 / 212 = 0
    16'b10011001_11010101 : OUT <= 0;  //153 / 213 = 0
    16'b10011001_11010110 : OUT <= 0;  //153 / 214 = 0
    16'b10011001_11010111 : OUT <= 0;  //153 / 215 = 0
    16'b10011001_11011000 : OUT <= 0;  //153 / 216 = 0
    16'b10011001_11011001 : OUT <= 0;  //153 / 217 = 0
    16'b10011001_11011010 : OUT <= 0;  //153 / 218 = 0
    16'b10011001_11011011 : OUT <= 0;  //153 / 219 = 0
    16'b10011001_11011100 : OUT <= 0;  //153 / 220 = 0
    16'b10011001_11011101 : OUT <= 0;  //153 / 221 = 0
    16'b10011001_11011110 : OUT <= 0;  //153 / 222 = 0
    16'b10011001_11011111 : OUT <= 0;  //153 / 223 = 0
    16'b10011001_11100000 : OUT <= 0;  //153 / 224 = 0
    16'b10011001_11100001 : OUT <= 0;  //153 / 225 = 0
    16'b10011001_11100010 : OUT <= 0;  //153 / 226 = 0
    16'b10011001_11100011 : OUT <= 0;  //153 / 227 = 0
    16'b10011001_11100100 : OUT <= 0;  //153 / 228 = 0
    16'b10011001_11100101 : OUT <= 0;  //153 / 229 = 0
    16'b10011001_11100110 : OUT <= 0;  //153 / 230 = 0
    16'b10011001_11100111 : OUT <= 0;  //153 / 231 = 0
    16'b10011001_11101000 : OUT <= 0;  //153 / 232 = 0
    16'b10011001_11101001 : OUT <= 0;  //153 / 233 = 0
    16'b10011001_11101010 : OUT <= 0;  //153 / 234 = 0
    16'b10011001_11101011 : OUT <= 0;  //153 / 235 = 0
    16'b10011001_11101100 : OUT <= 0;  //153 / 236 = 0
    16'b10011001_11101101 : OUT <= 0;  //153 / 237 = 0
    16'b10011001_11101110 : OUT <= 0;  //153 / 238 = 0
    16'b10011001_11101111 : OUT <= 0;  //153 / 239 = 0
    16'b10011001_11110000 : OUT <= 0;  //153 / 240 = 0
    16'b10011001_11110001 : OUT <= 0;  //153 / 241 = 0
    16'b10011001_11110010 : OUT <= 0;  //153 / 242 = 0
    16'b10011001_11110011 : OUT <= 0;  //153 / 243 = 0
    16'b10011001_11110100 : OUT <= 0;  //153 / 244 = 0
    16'b10011001_11110101 : OUT <= 0;  //153 / 245 = 0
    16'b10011001_11110110 : OUT <= 0;  //153 / 246 = 0
    16'b10011001_11110111 : OUT <= 0;  //153 / 247 = 0
    16'b10011001_11111000 : OUT <= 0;  //153 / 248 = 0
    16'b10011001_11111001 : OUT <= 0;  //153 / 249 = 0
    16'b10011001_11111010 : OUT <= 0;  //153 / 250 = 0
    16'b10011001_11111011 : OUT <= 0;  //153 / 251 = 0
    16'b10011001_11111100 : OUT <= 0;  //153 / 252 = 0
    16'b10011001_11111101 : OUT <= 0;  //153 / 253 = 0
    16'b10011001_11111110 : OUT <= 0;  //153 / 254 = 0
    16'b10011001_11111111 : OUT <= 0;  //153 / 255 = 0
    16'b10011010_00000000 : OUT <= 0;  //154 / 0 = 0
    16'b10011010_00000001 : OUT <= 154;  //154 / 1 = 154
    16'b10011010_00000010 : OUT <= 77;  //154 / 2 = 77
    16'b10011010_00000011 : OUT <= 51;  //154 / 3 = 51
    16'b10011010_00000100 : OUT <= 38;  //154 / 4 = 38
    16'b10011010_00000101 : OUT <= 30;  //154 / 5 = 30
    16'b10011010_00000110 : OUT <= 25;  //154 / 6 = 25
    16'b10011010_00000111 : OUT <= 22;  //154 / 7 = 22
    16'b10011010_00001000 : OUT <= 19;  //154 / 8 = 19
    16'b10011010_00001001 : OUT <= 17;  //154 / 9 = 17
    16'b10011010_00001010 : OUT <= 15;  //154 / 10 = 15
    16'b10011010_00001011 : OUT <= 14;  //154 / 11 = 14
    16'b10011010_00001100 : OUT <= 12;  //154 / 12 = 12
    16'b10011010_00001101 : OUT <= 11;  //154 / 13 = 11
    16'b10011010_00001110 : OUT <= 11;  //154 / 14 = 11
    16'b10011010_00001111 : OUT <= 10;  //154 / 15 = 10
    16'b10011010_00010000 : OUT <= 9;  //154 / 16 = 9
    16'b10011010_00010001 : OUT <= 9;  //154 / 17 = 9
    16'b10011010_00010010 : OUT <= 8;  //154 / 18 = 8
    16'b10011010_00010011 : OUT <= 8;  //154 / 19 = 8
    16'b10011010_00010100 : OUT <= 7;  //154 / 20 = 7
    16'b10011010_00010101 : OUT <= 7;  //154 / 21 = 7
    16'b10011010_00010110 : OUT <= 7;  //154 / 22 = 7
    16'b10011010_00010111 : OUT <= 6;  //154 / 23 = 6
    16'b10011010_00011000 : OUT <= 6;  //154 / 24 = 6
    16'b10011010_00011001 : OUT <= 6;  //154 / 25 = 6
    16'b10011010_00011010 : OUT <= 5;  //154 / 26 = 5
    16'b10011010_00011011 : OUT <= 5;  //154 / 27 = 5
    16'b10011010_00011100 : OUT <= 5;  //154 / 28 = 5
    16'b10011010_00011101 : OUT <= 5;  //154 / 29 = 5
    16'b10011010_00011110 : OUT <= 5;  //154 / 30 = 5
    16'b10011010_00011111 : OUT <= 4;  //154 / 31 = 4
    16'b10011010_00100000 : OUT <= 4;  //154 / 32 = 4
    16'b10011010_00100001 : OUT <= 4;  //154 / 33 = 4
    16'b10011010_00100010 : OUT <= 4;  //154 / 34 = 4
    16'b10011010_00100011 : OUT <= 4;  //154 / 35 = 4
    16'b10011010_00100100 : OUT <= 4;  //154 / 36 = 4
    16'b10011010_00100101 : OUT <= 4;  //154 / 37 = 4
    16'b10011010_00100110 : OUT <= 4;  //154 / 38 = 4
    16'b10011010_00100111 : OUT <= 3;  //154 / 39 = 3
    16'b10011010_00101000 : OUT <= 3;  //154 / 40 = 3
    16'b10011010_00101001 : OUT <= 3;  //154 / 41 = 3
    16'b10011010_00101010 : OUT <= 3;  //154 / 42 = 3
    16'b10011010_00101011 : OUT <= 3;  //154 / 43 = 3
    16'b10011010_00101100 : OUT <= 3;  //154 / 44 = 3
    16'b10011010_00101101 : OUT <= 3;  //154 / 45 = 3
    16'b10011010_00101110 : OUT <= 3;  //154 / 46 = 3
    16'b10011010_00101111 : OUT <= 3;  //154 / 47 = 3
    16'b10011010_00110000 : OUT <= 3;  //154 / 48 = 3
    16'b10011010_00110001 : OUT <= 3;  //154 / 49 = 3
    16'b10011010_00110010 : OUT <= 3;  //154 / 50 = 3
    16'b10011010_00110011 : OUT <= 3;  //154 / 51 = 3
    16'b10011010_00110100 : OUT <= 2;  //154 / 52 = 2
    16'b10011010_00110101 : OUT <= 2;  //154 / 53 = 2
    16'b10011010_00110110 : OUT <= 2;  //154 / 54 = 2
    16'b10011010_00110111 : OUT <= 2;  //154 / 55 = 2
    16'b10011010_00111000 : OUT <= 2;  //154 / 56 = 2
    16'b10011010_00111001 : OUT <= 2;  //154 / 57 = 2
    16'b10011010_00111010 : OUT <= 2;  //154 / 58 = 2
    16'b10011010_00111011 : OUT <= 2;  //154 / 59 = 2
    16'b10011010_00111100 : OUT <= 2;  //154 / 60 = 2
    16'b10011010_00111101 : OUT <= 2;  //154 / 61 = 2
    16'b10011010_00111110 : OUT <= 2;  //154 / 62 = 2
    16'b10011010_00111111 : OUT <= 2;  //154 / 63 = 2
    16'b10011010_01000000 : OUT <= 2;  //154 / 64 = 2
    16'b10011010_01000001 : OUT <= 2;  //154 / 65 = 2
    16'b10011010_01000010 : OUT <= 2;  //154 / 66 = 2
    16'b10011010_01000011 : OUT <= 2;  //154 / 67 = 2
    16'b10011010_01000100 : OUT <= 2;  //154 / 68 = 2
    16'b10011010_01000101 : OUT <= 2;  //154 / 69 = 2
    16'b10011010_01000110 : OUT <= 2;  //154 / 70 = 2
    16'b10011010_01000111 : OUT <= 2;  //154 / 71 = 2
    16'b10011010_01001000 : OUT <= 2;  //154 / 72 = 2
    16'b10011010_01001001 : OUT <= 2;  //154 / 73 = 2
    16'b10011010_01001010 : OUT <= 2;  //154 / 74 = 2
    16'b10011010_01001011 : OUT <= 2;  //154 / 75 = 2
    16'b10011010_01001100 : OUT <= 2;  //154 / 76 = 2
    16'b10011010_01001101 : OUT <= 2;  //154 / 77 = 2
    16'b10011010_01001110 : OUT <= 1;  //154 / 78 = 1
    16'b10011010_01001111 : OUT <= 1;  //154 / 79 = 1
    16'b10011010_01010000 : OUT <= 1;  //154 / 80 = 1
    16'b10011010_01010001 : OUT <= 1;  //154 / 81 = 1
    16'b10011010_01010010 : OUT <= 1;  //154 / 82 = 1
    16'b10011010_01010011 : OUT <= 1;  //154 / 83 = 1
    16'b10011010_01010100 : OUT <= 1;  //154 / 84 = 1
    16'b10011010_01010101 : OUT <= 1;  //154 / 85 = 1
    16'b10011010_01010110 : OUT <= 1;  //154 / 86 = 1
    16'b10011010_01010111 : OUT <= 1;  //154 / 87 = 1
    16'b10011010_01011000 : OUT <= 1;  //154 / 88 = 1
    16'b10011010_01011001 : OUT <= 1;  //154 / 89 = 1
    16'b10011010_01011010 : OUT <= 1;  //154 / 90 = 1
    16'b10011010_01011011 : OUT <= 1;  //154 / 91 = 1
    16'b10011010_01011100 : OUT <= 1;  //154 / 92 = 1
    16'b10011010_01011101 : OUT <= 1;  //154 / 93 = 1
    16'b10011010_01011110 : OUT <= 1;  //154 / 94 = 1
    16'b10011010_01011111 : OUT <= 1;  //154 / 95 = 1
    16'b10011010_01100000 : OUT <= 1;  //154 / 96 = 1
    16'b10011010_01100001 : OUT <= 1;  //154 / 97 = 1
    16'b10011010_01100010 : OUT <= 1;  //154 / 98 = 1
    16'b10011010_01100011 : OUT <= 1;  //154 / 99 = 1
    16'b10011010_01100100 : OUT <= 1;  //154 / 100 = 1
    16'b10011010_01100101 : OUT <= 1;  //154 / 101 = 1
    16'b10011010_01100110 : OUT <= 1;  //154 / 102 = 1
    16'b10011010_01100111 : OUT <= 1;  //154 / 103 = 1
    16'b10011010_01101000 : OUT <= 1;  //154 / 104 = 1
    16'b10011010_01101001 : OUT <= 1;  //154 / 105 = 1
    16'b10011010_01101010 : OUT <= 1;  //154 / 106 = 1
    16'b10011010_01101011 : OUT <= 1;  //154 / 107 = 1
    16'b10011010_01101100 : OUT <= 1;  //154 / 108 = 1
    16'b10011010_01101101 : OUT <= 1;  //154 / 109 = 1
    16'b10011010_01101110 : OUT <= 1;  //154 / 110 = 1
    16'b10011010_01101111 : OUT <= 1;  //154 / 111 = 1
    16'b10011010_01110000 : OUT <= 1;  //154 / 112 = 1
    16'b10011010_01110001 : OUT <= 1;  //154 / 113 = 1
    16'b10011010_01110010 : OUT <= 1;  //154 / 114 = 1
    16'b10011010_01110011 : OUT <= 1;  //154 / 115 = 1
    16'b10011010_01110100 : OUT <= 1;  //154 / 116 = 1
    16'b10011010_01110101 : OUT <= 1;  //154 / 117 = 1
    16'b10011010_01110110 : OUT <= 1;  //154 / 118 = 1
    16'b10011010_01110111 : OUT <= 1;  //154 / 119 = 1
    16'b10011010_01111000 : OUT <= 1;  //154 / 120 = 1
    16'b10011010_01111001 : OUT <= 1;  //154 / 121 = 1
    16'b10011010_01111010 : OUT <= 1;  //154 / 122 = 1
    16'b10011010_01111011 : OUT <= 1;  //154 / 123 = 1
    16'b10011010_01111100 : OUT <= 1;  //154 / 124 = 1
    16'b10011010_01111101 : OUT <= 1;  //154 / 125 = 1
    16'b10011010_01111110 : OUT <= 1;  //154 / 126 = 1
    16'b10011010_01111111 : OUT <= 1;  //154 / 127 = 1
    16'b10011010_10000000 : OUT <= 1;  //154 / 128 = 1
    16'b10011010_10000001 : OUT <= 1;  //154 / 129 = 1
    16'b10011010_10000010 : OUT <= 1;  //154 / 130 = 1
    16'b10011010_10000011 : OUT <= 1;  //154 / 131 = 1
    16'b10011010_10000100 : OUT <= 1;  //154 / 132 = 1
    16'b10011010_10000101 : OUT <= 1;  //154 / 133 = 1
    16'b10011010_10000110 : OUT <= 1;  //154 / 134 = 1
    16'b10011010_10000111 : OUT <= 1;  //154 / 135 = 1
    16'b10011010_10001000 : OUT <= 1;  //154 / 136 = 1
    16'b10011010_10001001 : OUT <= 1;  //154 / 137 = 1
    16'b10011010_10001010 : OUT <= 1;  //154 / 138 = 1
    16'b10011010_10001011 : OUT <= 1;  //154 / 139 = 1
    16'b10011010_10001100 : OUT <= 1;  //154 / 140 = 1
    16'b10011010_10001101 : OUT <= 1;  //154 / 141 = 1
    16'b10011010_10001110 : OUT <= 1;  //154 / 142 = 1
    16'b10011010_10001111 : OUT <= 1;  //154 / 143 = 1
    16'b10011010_10010000 : OUT <= 1;  //154 / 144 = 1
    16'b10011010_10010001 : OUT <= 1;  //154 / 145 = 1
    16'b10011010_10010010 : OUT <= 1;  //154 / 146 = 1
    16'b10011010_10010011 : OUT <= 1;  //154 / 147 = 1
    16'b10011010_10010100 : OUT <= 1;  //154 / 148 = 1
    16'b10011010_10010101 : OUT <= 1;  //154 / 149 = 1
    16'b10011010_10010110 : OUT <= 1;  //154 / 150 = 1
    16'b10011010_10010111 : OUT <= 1;  //154 / 151 = 1
    16'b10011010_10011000 : OUT <= 1;  //154 / 152 = 1
    16'b10011010_10011001 : OUT <= 1;  //154 / 153 = 1
    16'b10011010_10011010 : OUT <= 1;  //154 / 154 = 1
    16'b10011010_10011011 : OUT <= 0;  //154 / 155 = 0
    16'b10011010_10011100 : OUT <= 0;  //154 / 156 = 0
    16'b10011010_10011101 : OUT <= 0;  //154 / 157 = 0
    16'b10011010_10011110 : OUT <= 0;  //154 / 158 = 0
    16'b10011010_10011111 : OUT <= 0;  //154 / 159 = 0
    16'b10011010_10100000 : OUT <= 0;  //154 / 160 = 0
    16'b10011010_10100001 : OUT <= 0;  //154 / 161 = 0
    16'b10011010_10100010 : OUT <= 0;  //154 / 162 = 0
    16'b10011010_10100011 : OUT <= 0;  //154 / 163 = 0
    16'b10011010_10100100 : OUT <= 0;  //154 / 164 = 0
    16'b10011010_10100101 : OUT <= 0;  //154 / 165 = 0
    16'b10011010_10100110 : OUT <= 0;  //154 / 166 = 0
    16'b10011010_10100111 : OUT <= 0;  //154 / 167 = 0
    16'b10011010_10101000 : OUT <= 0;  //154 / 168 = 0
    16'b10011010_10101001 : OUT <= 0;  //154 / 169 = 0
    16'b10011010_10101010 : OUT <= 0;  //154 / 170 = 0
    16'b10011010_10101011 : OUT <= 0;  //154 / 171 = 0
    16'b10011010_10101100 : OUT <= 0;  //154 / 172 = 0
    16'b10011010_10101101 : OUT <= 0;  //154 / 173 = 0
    16'b10011010_10101110 : OUT <= 0;  //154 / 174 = 0
    16'b10011010_10101111 : OUT <= 0;  //154 / 175 = 0
    16'b10011010_10110000 : OUT <= 0;  //154 / 176 = 0
    16'b10011010_10110001 : OUT <= 0;  //154 / 177 = 0
    16'b10011010_10110010 : OUT <= 0;  //154 / 178 = 0
    16'b10011010_10110011 : OUT <= 0;  //154 / 179 = 0
    16'b10011010_10110100 : OUT <= 0;  //154 / 180 = 0
    16'b10011010_10110101 : OUT <= 0;  //154 / 181 = 0
    16'b10011010_10110110 : OUT <= 0;  //154 / 182 = 0
    16'b10011010_10110111 : OUT <= 0;  //154 / 183 = 0
    16'b10011010_10111000 : OUT <= 0;  //154 / 184 = 0
    16'b10011010_10111001 : OUT <= 0;  //154 / 185 = 0
    16'b10011010_10111010 : OUT <= 0;  //154 / 186 = 0
    16'b10011010_10111011 : OUT <= 0;  //154 / 187 = 0
    16'b10011010_10111100 : OUT <= 0;  //154 / 188 = 0
    16'b10011010_10111101 : OUT <= 0;  //154 / 189 = 0
    16'b10011010_10111110 : OUT <= 0;  //154 / 190 = 0
    16'b10011010_10111111 : OUT <= 0;  //154 / 191 = 0
    16'b10011010_11000000 : OUT <= 0;  //154 / 192 = 0
    16'b10011010_11000001 : OUT <= 0;  //154 / 193 = 0
    16'b10011010_11000010 : OUT <= 0;  //154 / 194 = 0
    16'b10011010_11000011 : OUT <= 0;  //154 / 195 = 0
    16'b10011010_11000100 : OUT <= 0;  //154 / 196 = 0
    16'b10011010_11000101 : OUT <= 0;  //154 / 197 = 0
    16'b10011010_11000110 : OUT <= 0;  //154 / 198 = 0
    16'b10011010_11000111 : OUT <= 0;  //154 / 199 = 0
    16'b10011010_11001000 : OUT <= 0;  //154 / 200 = 0
    16'b10011010_11001001 : OUT <= 0;  //154 / 201 = 0
    16'b10011010_11001010 : OUT <= 0;  //154 / 202 = 0
    16'b10011010_11001011 : OUT <= 0;  //154 / 203 = 0
    16'b10011010_11001100 : OUT <= 0;  //154 / 204 = 0
    16'b10011010_11001101 : OUT <= 0;  //154 / 205 = 0
    16'b10011010_11001110 : OUT <= 0;  //154 / 206 = 0
    16'b10011010_11001111 : OUT <= 0;  //154 / 207 = 0
    16'b10011010_11010000 : OUT <= 0;  //154 / 208 = 0
    16'b10011010_11010001 : OUT <= 0;  //154 / 209 = 0
    16'b10011010_11010010 : OUT <= 0;  //154 / 210 = 0
    16'b10011010_11010011 : OUT <= 0;  //154 / 211 = 0
    16'b10011010_11010100 : OUT <= 0;  //154 / 212 = 0
    16'b10011010_11010101 : OUT <= 0;  //154 / 213 = 0
    16'b10011010_11010110 : OUT <= 0;  //154 / 214 = 0
    16'b10011010_11010111 : OUT <= 0;  //154 / 215 = 0
    16'b10011010_11011000 : OUT <= 0;  //154 / 216 = 0
    16'b10011010_11011001 : OUT <= 0;  //154 / 217 = 0
    16'b10011010_11011010 : OUT <= 0;  //154 / 218 = 0
    16'b10011010_11011011 : OUT <= 0;  //154 / 219 = 0
    16'b10011010_11011100 : OUT <= 0;  //154 / 220 = 0
    16'b10011010_11011101 : OUT <= 0;  //154 / 221 = 0
    16'b10011010_11011110 : OUT <= 0;  //154 / 222 = 0
    16'b10011010_11011111 : OUT <= 0;  //154 / 223 = 0
    16'b10011010_11100000 : OUT <= 0;  //154 / 224 = 0
    16'b10011010_11100001 : OUT <= 0;  //154 / 225 = 0
    16'b10011010_11100010 : OUT <= 0;  //154 / 226 = 0
    16'b10011010_11100011 : OUT <= 0;  //154 / 227 = 0
    16'b10011010_11100100 : OUT <= 0;  //154 / 228 = 0
    16'b10011010_11100101 : OUT <= 0;  //154 / 229 = 0
    16'b10011010_11100110 : OUT <= 0;  //154 / 230 = 0
    16'b10011010_11100111 : OUT <= 0;  //154 / 231 = 0
    16'b10011010_11101000 : OUT <= 0;  //154 / 232 = 0
    16'b10011010_11101001 : OUT <= 0;  //154 / 233 = 0
    16'b10011010_11101010 : OUT <= 0;  //154 / 234 = 0
    16'b10011010_11101011 : OUT <= 0;  //154 / 235 = 0
    16'b10011010_11101100 : OUT <= 0;  //154 / 236 = 0
    16'b10011010_11101101 : OUT <= 0;  //154 / 237 = 0
    16'b10011010_11101110 : OUT <= 0;  //154 / 238 = 0
    16'b10011010_11101111 : OUT <= 0;  //154 / 239 = 0
    16'b10011010_11110000 : OUT <= 0;  //154 / 240 = 0
    16'b10011010_11110001 : OUT <= 0;  //154 / 241 = 0
    16'b10011010_11110010 : OUT <= 0;  //154 / 242 = 0
    16'b10011010_11110011 : OUT <= 0;  //154 / 243 = 0
    16'b10011010_11110100 : OUT <= 0;  //154 / 244 = 0
    16'b10011010_11110101 : OUT <= 0;  //154 / 245 = 0
    16'b10011010_11110110 : OUT <= 0;  //154 / 246 = 0
    16'b10011010_11110111 : OUT <= 0;  //154 / 247 = 0
    16'b10011010_11111000 : OUT <= 0;  //154 / 248 = 0
    16'b10011010_11111001 : OUT <= 0;  //154 / 249 = 0
    16'b10011010_11111010 : OUT <= 0;  //154 / 250 = 0
    16'b10011010_11111011 : OUT <= 0;  //154 / 251 = 0
    16'b10011010_11111100 : OUT <= 0;  //154 / 252 = 0
    16'b10011010_11111101 : OUT <= 0;  //154 / 253 = 0
    16'b10011010_11111110 : OUT <= 0;  //154 / 254 = 0
    16'b10011010_11111111 : OUT <= 0;  //154 / 255 = 0
    16'b10011011_00000000 : OUT <= 0;  //155 / 0 = 0
    16'b10011011_00000001 : OUT <= 155;  //155 / 1 = 155
    16'b10011011_00000010 : OUT <= 77;  //155 / 2 = 77
    16'b10011011_00000011 : OUT <= 51;  //155 / 3 = 51
    16'b10011011_00000100 : OUT <= 38;  //155 / 4 = 38
    16'b10011011_00000101 : OUT <= 31;  //155 / 5 = 31
    16'b10011011_00000110 : OUT <= 25;  //155 / 6 = 25
    16'b10011011_00000111 : OUT <= 22;  //155 / 7 = 22
    16'b10011011_00001000 : OUT <= 19;  //155 / 8 = 19
    16'b10011011_00001001 : OUT <= 17;  //155 / 9 = 17
    16'b10011011_00001010 : OUT <= 15;  //155 / 10 = 15
    16'b10011011_00001011 : OUT <= 14;  //155 / 11 = 14
    16'b10011011_00001100 : OUT <= 12;  //155 / 12 = 12
    16'b10011011_00001101 : OUT <= 11;  //155 / 13 = 11
    16'b10011011_00001110 : OUT <= 11;  //155 / 14 = 11
    16'b10011011_00001111 : OUT <= 10;  //155 / 15 = 10
    16'b10011011_00010000 : OUT <= 9;  //155 / 16 = 9
    16'b10011011_00010001 : OUT <= 9;  //155 / 17 = 9
    16'b10011011_00010010 : OUT <= 8;  //155 / 18 = 8
    16'b10011011_00010011 : OUT <= 8;  //155 / 19 = 8
    16'b10011011_00010100 : OUT <= 7;  //155 / 20 = 7
    16'b10011011_00010101 : OUT <= 7;  //155 / 21 = 7
    16'b10011011_00010110 : OUT <= 7;  //155 / 22 = 7
    16'b10011011_00010111 : OUT <= 6;  //155 / 23 = 6
    16'b10011011_00011000 : OUT <= 6;  //155 / 24 = 6
    16'b10011011_00011001 : OUT <= 6;  //155 / 25 = 6
    16'b10011011_00011010 : OUT <= 5;  //155 / 26 = 5
    16'b10011011_00011011 : OUT <= 5;  //155 / 27 = 5
    16'b10011011_00011100 : OUT <= 5;  //155 / 28 = 5
    16'b10011011_00011101 : OUT <= 5;  //155 / 29 = 5
    16'b10011011_00011110 : OUT <= 5;  //155 / 30 = 5
    16'b10011011_00011111 : OUT <= 5;  //155 / 31 = 5
    16'b10011011_00100000 : OUT <= 4;  //155 / 32 = 4
    16'b10011011_00100001 : OUT <= 4;  //155 / 33 = 4
    16'b10011011_00100010 : OUT <= 4;  //155 / 34 = 4
    16'b10011011_00100011 : OUT <= 4;  //155 / 35 = 4
    16'b10011011_00100100 : OUT <= 4;  //155 / 36 = 4
    16'b10011011_00100101 : OUT <= 4;  //155 / 37 = 4
    16'b10011011_00100110 : OUT <= 4;  //155 / 38 = 4
    16'b10011011_00100111 : OUT <= 3;  //155 / 39 = 3
    16'b10011011_00101000 : OUT <= 3;  //155 / 40 = 3
    16'b10011011_00101001 : OUT <= 3;  //155 / 41 = 3
    16'b10011011_00101010 : OUT <= 3;  //155 / 42 = 3
    16'b10011011_00101011 : OUT <= 3;  //155 / 43 = 3
    16'b10011011_00101100 : OUT <= 3;  //155 / 44 = 3
    16'b10011011_00101101 : OUT <= 3;  //155 / 45 = 3
    16'b10011011_00101110 : OUT <= 3;  //155 / 46 = 3
    16'b10011011_00101111 : OUT <= 3;  //155 / 47 = 3
    16'b10011011_00110000 : OUT <= 3;  //155 / 48 = 3
    16'b10011011_00110001 : OUT <= 3;  //155 / 49 = 3
    16'b10011011_00110010 : OUT <= 3;  //155 / 50 = 3
    16'b10011011_00110011 : OUT <= 3;  //155 / 51 = 3
    16'b10011011_00110100 : OUT <= 2;  //155 / 52 = 2
    16'b10011011_00110101 : OUT <= 2;  //155 / 53 = 2
    16'b10011011_00110110 : OUT <= 2;  //155 / 54 = 2
    16'b10011011_00110111 : OUT <= 2;  //155 / 55 = 2
    16'b10011011_00111000 : OUT <= 2;  //155 / 56 = 2
    16'b10011011_00111001 : OUT <= 2;  //155 / 57 = 2
    16'b10011011_00111010 : OUT <= 2;  //155 / 58 = 2
    16'b10011011_00111011 : OUT <= 2;  //155 / 59 = 2
    16'b10011011_00111100 : OUT <= 2;  //155 / 60 = 2
    16'b10011011_00111101 : OUT <= 2;  //155 / 61 = 2
    16'b10011011_00111110 : OUT <= 2;  //155 / 62 = 2
    16'b10011011_00111111 : OUT <= 2;  //155 / 63 = 2
    16'b10011011_01000000 : OUT <= 2;  //155 / 64 = 2
    16'b10011011_01000001 : OUT <= 2;  //155 / 65 = 2
    16'b10011011_01000010 : OUT <= 2;  //155 / 66 = 2
    16'b10011011_01000011 : OUT <= 2;  //155 / 67 = 2
    16'b10011011_01000100 : OUT <= 2;  //155 / 68 = 2
    16'b10011011_01000101 : OUT <= 2;  //155 / 69 = 2
    16'b10011011_01000110 : OUT <= 2;  //155 / 70 = 2
    16'b10011011_01000111 : OUT <= 2;  //155 / 71 = 2
    16'b10011011_01001000 : OUT <= 2;  //155 / 72 = 2
    16'b10011011_01001001 : OUT <= 2;  //155 / 73 = 2
    16'b10011011_01001010 : OUT <= 2;  //155 / 74 = 2
    16'b10011011_01001011 : OUT <= 2;  //155 / 75 = 2
    16'b10011011_01001100 : OUT <= 2;  //155 / 76 = 2
    16'b10011011_01001101 : OUT <= 2;  //155 / 77 = 2
    16'b10011011_01001110 : OUT <= 1;  //155 / 78 = 1
    16'b10011011_01001111 : OUT <= 1;  //155 / 79 = 1
    16'b10011011_01010000 : OUT <= 1;  //155 / 80 = 1
    16'b10011011_01010001 : OUT <= 1;  //155 / 81 = 1
    16'b10011011_01010010 : OUT <= 1;  //155 / 82 = 1
    16'b10011011_01010011 : OUT <= 1;  //155 / 83 = 1
    16'b10011011_01010100 : OUT <= 1;  //155 / 84 = 1
    16'b10011011_01010101 : OUT <= 1;  //155 / 85 = 1
    16'b10011011_01010110 : OUT <= 1;  //155 / 86 = 1
    16'b10011011_01010111 : OUT <= 1;  //155 / 87 = 1
    16'b10011011_01011000 : OUT <= 1;  //155 / 88 = 1
    16'b10011011_01011001 : OUT <= 1;  //155 / 89 = 1
    16'b10011011_01011010 : OUT <= 1;  //155 / 90 = 1
    16'b10011011_01011011 : OUT <= 1;  //155 / 91 = 1
    16'b10011011_01011100 : OUT <= 1;  //155 / 92 = 1
    16'b10011011_01011101 : OUT <= 1;  //155 / 93 = 1
    16'b10011011_01011110 : OUT <= 1;  //155 / 94 = 1
    16'b10011011_01011111 : OUT <= 1;  //155 / 95 = 1
    16'b10011011_01100000 : OUT <= 1;  //155 / 96 = 1
    16'b10011011_01100001 : OUT <= 1;  //155 / 97 = 1
    16'b10011011_01100010 : OUT <= 1;  //155 / 98 = 1
    16'b10011011_01100011 : OUT <= 1;  //155 / 99 = 1
    16'b10011011_01100100 : OUT <= 1;  //155 / 100 = 1
    16'b10011011_01100101 : OUT <= 1;  //155 / 101 = 1
    16'b10011011_01100110 : OUT <= 1;  //155 / 102 = 1
    16'b10011011_01100111 : OUT <= 1;  //155 / 103 = 1
    16'b10011011_01101000 : OUT <= 1;  //155 / 104 = 1
    16'b10011011_01101001 : OUT <= 1;  //155 / 105 = 1
    16'b10011011_01101010 : OUT <= 1;  //155 / 106 = 1
    16'b10011011_01101011 : OUT <= 1;  //155 / 107 = 1
    16'b10011011_01101100 : OUT <= 1;  //155 / 108 = 1
    16'b10011011_01101101 : OUT <= 1;  //155 / 109 = 1
    16'b10011011_01101110 : OUT <= 1;  //155 / 110 = 1
    16'b10011011_01101111 : OUT <= 1;  //155 / 111 = 1
    16'b10011011_01110000 : OUT <= 1;  //155 / 112 = 1
    16'b10011011_01110001 : OUT <= 1;  //155 / 113 = 1
    16'b10011011_01110010 : OUT <= 1;  //155 / 114 = 1
    16'b10011011_01110011 : OUT <= 1;  //155 / 115 = 1
    16'b10011011_01110100 : OUT <= 1;  //155 / 116 = 1
    16'b10011011_01110101 : OUT <= 1;  //155 / 117 = 1
    16'b10011011_01110110 : OUT <= 1;  //155 / 118 = 1
    16'b10011011_01110111 : OUT <= 1;  //155 / 119 = 1
    16'b10011011_01111000 : OUT <= 1;  //155 / 120 = 1
    16'b10011011_01111001 : OUT <= 1;  //155 / 121 = 1
    16'b10011011_01111010 : OUT <= 1;  //155 / 122 = 1
    16'b10011011_01111011 : OUT <= 1;  //155 / 123 = 1
    16'b10011011_01111100 : OUT <= 1;  //155 / 124 = 1
    16'b10011011_01111101 : OUT <= 1;  //155 / 125 = 1
    16'b10011011_01111110 : OUT <= 1;  //155 / 126 = 1
    16'b10011011_01111111 : OUT <= 1;  //155 / 127 = 1
    16'b10011011_10000000 : OUT <= 1;  //155 / 128 = 1
    16'b10011011_10000001 : OUT <= 1;  //155 / 129 = 1
    16'b10011011_10000010 : OUT <= 1;  //155 / 130 = 1
    16'b10011011_10000011 : OUT <= 1;  //155 / 131 = 1
    16'b10011011_10000100 : OUT <= 1;  //155 / 132 = 1
    16'b10011011_10000101 : OUT <= 1;  //155 / 133 = 1
    16'b10011011_10000110 : OUT <= 1;  //155 / 134 = 1
    16'b10011011_10000111 : OUT <= 1;  //155 / 135 = 1
    16'b10011011_10001000 : OUT <= 1;  //155 / 136 = 1
    16'b10011011_10001001 : OUT <= 1;  //155 / 137 = 1
    16'b10011011_10001010 : OUT <= 1;  //155 / 138 = 1
    16'b10011011_10001011 : OUT <= 1;  //155 / 139 = 1
    16'b10011011_10001100 : OUT <= 1;  //155 / 140 = 1
    16'b10011011_10001101 : OUT <= 1;  //155 / 141 = 1
    16'b10011011_10001110 : OUT <= 1;  //155 / 142 = 1
    16'b10011011_10001111 : OUT <= 1;  //155 / 143 = 1
    16'b10011011_10010000 : OUT <= 1;  //155 / 144 = 1
    16'b10011011_10010001 : OUT <= 1;  //155 / 145 = 1
    16'b10011011_10010010 : OUT <= 1;  //155 / 146 = 1
    16'b10011011_10010011 : OUT <= 1;  //155 / 147 = 1
    16'b10011011_10010100 : OUT <= 1;  //155 / 148 = 1
    16'b10011011_10010101 : OUT <= 1;  //155 / 149 = 1
    16'b10011011_10010110 : OUT <= 1;  //155 / 150 = 1
    16'b10011011_10010111 : OUT <= 1;  //155 / 151 = 1
    16'b10011011_10011000 : OUT <= 1;  //155 / 152 = 1
    16'b10011011_10011001 : OUT <= 1;  //155 / 153 = 1
    16'b10011011_10011010 : OUT <= 1;  //155 / 154 = 1
    16'b10011011_10011011 : OUT <= 1;  //155 / 155 = 1
    16'b10011011_10011100 : OUT <= 0;  //155 / 156 = 0
    16'b10011011_10011101 : OUT <= 0;  //155 / 157 = 0
    16'b10011011_10011110 : OUT <= 0;  //155 / 158 = 0
    16'b10011011_10011111 : OUT <= 0;  //155 / 159 = 0
    16'b10011011_10100000 : OUT <= 0;  //155 / 160 = 0
    16'b10011011_10100001 : OUT <= 0;  //155 / 161 = 0
    16'b10011011_10100010 : OUT <= 0;  //155 / 162 = 0
    16'b10011011_10100011 : OUT <= 0;  //155 / 163 = 0
    16'b10011011_10100100 : OUT <= 0;  //155 / 164 = 0
    16'b10011011_10100101 : OUT <= 0;  //155 / 165 = 0
    16'b10011011_10100110 : OUT <= 0;  //155 / 166 = 0
    16'b10011011_10100111 : OUT <= 0;  //155 / 167 = 0
    16'b10011011_10101000 : OUT <= 0;  //155 / 168 = 0
    16'b10011011_10101001 : OUT <= 0;  //155 / 169 = 0
    16'b10011011_10101010 : OUT <= 0;  //155 / 170 = 0
    16'b10011011_10101011 : OUT <= 0;  //155 / 171 = 0
    16'b10011011_10101100 : OUT <= 0;  //155 / 172 = 0
    16'b10011011_10101101 : OUT <= 0;  //155 / 173 = 0
    16'b10011011_10101110 : OUT <= 0;  //155 / 174 = 0
    16'b10011011_10101111 : OUT <= 0;  //155 / 175 = 0
    16'b10011011_10110000 : OUT <= 0;  //155 / 176 = 0
    16'b10011011_10110001 : OUT <= 0;  //155 / 177 = 0
    16'b10011011_10110010 : OUT <= 0;  //155 / 178 = 0
    16'b10011011_10110011 : OUT <= 0;  //155 / 179 = 0
    16'b10011011_10110100 : OUT <= 0;  //155 / 180 = 0
    16'b10011011_10110101 : OUT <= 0;  //155 / 181 = 0
    16'b10011011_10110110 : OUT <= 0;  //155 / 182 = 0
    16'b10011011_10110111 : OUT <= 0;  //155 / 183 = 0
    16'b10011011_10111000 : OUT <= 0;  //155 / 184 = 0
    16'b10011011_10111001 : OUT <= 0;  //155 / 185 = 0
    16'b10011011_10111010 : OUT <= 0;  //155 / 186 = 0
    16'b10011011_10111011 : OUT <= 0;  //155 / 187 = 0
    16'b10011011_10111100 : OUT <= 0;  //155 / 188 = 0
    16'b10011011_10111101 : OUT <= 0;  //155 / 189 = 0
    16'b10011011_10111110 : OUT <= 0;  //155 / 190 = 0
    16'b10011011_10111111 : OUT <= 0;  //155 / 191 = 0
    16'b10011011_11000000 : OUT <= 0;  //155 / 192 = 0
    16'b10011011_11000001 : OUT <= 0;  //155 / 193 = 0
    16'b10011011_11000010 : OUT <= 0;  //155 / 194 = 0
    16'b10011011_11000011 : OUT <= 0;  //155 / 195 = 0
    16'b10011011_11000100 : OUT <= 0;  //155 / 196 = 0
    16'b10011011_11000101 : OUT <= 0;  //155 / 197 = 0
    16'b10011011_11000110 : OUT <= 0;  //155 / 198 = 0
    16'b10011011_11000111 : OUT <= 0;  //155 / 199 = 0
    16'b10011011_11001000 : OUT <= 0;  //155 / 200 = 0
    16'b10011011_11001001 : OUT <= 0;  //155 / 201 = 0
    16'b10011011_11001010 : OUT <= 0;  //155 / 202 = 0
    16'b10011011_11001011 : OUT <= 0;  //155 / 203 = 0
    16'b10011011_11001100 : OUT <= 0;  //155 / 204 = 0
    16'b10011011_11001101 : OUT <= 0;  //155 / 205 = 0
    16'b10011011_11001110 : OUT <= 0;  //155 / 206 = 0
    16'b10011011_11001111 : OUT <= 0;  //155 / 207 = 0
    16'b10011011_11010000 : OUT <= 0;  //155 / 208 = 0
    16'b10011011_11010001 : OUT <= 0;  //155 / 209 = 0
    16'b10011011_11010010 : OUT <= 0;  //155 / 210 = 0
    16'b10011011_11010011 : OUT <= 0;  //155 / 211 = 0
    16'b10011011_11010100 : OUT <= 0;  //155 / 212 = 0
    16'b10011011_11010101 : OUT <= 0;  //155 / 213 = 0
    16'b10011011_11010110 : OUT <= 0;  //155 / 214 = 0
    16'b10011011_11010111 : OUT <= 0;  //155 / 215 = 0
    16'b10011011_11011000 : OUT <= 0;  //155 / 216 = 0
    16'b10011011_11011001 : OUT <= 0;  //155 / 217 = 0
    16'b10011011_11011010 : OUT <= 0;  //155 / 218 = 0
    16'b10011011_11011011 : OUT <= 0;  //155 / 219 = 0
    16'b10011011_11011100 : OUT <= 0;  //155 / 220 = 0
    16'b10011011_11011101 : OUT <= 0;  //155 / 221 = 0
    16'b10011011_11011110 : OUT <= 0;  //155 / 222 = 0
    16'b10011011_11011111 : OUT <= 0;  //155 / 223 = 0
    16'b10011011_11100000 : OUT <= 0;  //155 / 224 = 0
    16'b10011011_11100001 : OUT <= 0;  //155 / 225 = 0
    16'b10011011_11100010 : OUT <= 0;  //155 / 226 = 0
    16'b10011011_11100011 : OUT <= 0;  //155 / 227 = 0
    16'b10011011_11100100 : OUT <= 0;  //155 / 228 = 0
    16'b10011011_11100101 : OUT <= 0;  //155 / 229 = 0
    16'b10011011_11100110 : OUT <= 0;  //155 / 230 = 0
    16'b10011011_11100111 : OUT <= 0;  //155 / 231 = 0
    16'b10011011_11101000 : OUT <= 0;  //155 / 232 = 0
    16'b10011011_11101001 : OUT <= 0;  //155 / 233 = 0
    16'b10011011_11101010 : OUT <= 0;  //155 / 234 = 0
    16'b10011011_11101011 : OUT <= 0;  //155 / 235 = 0
    16'b10011011_11101100 : OUT <= 0;  //155 / 236 = 0
    16'b10011011_11101101 : OUT <= 0;  //155 / 237 = 0
    16'b10011011_11101110 : OUT <= 0;  //155 / 238 = 0
    16'b10011011_11101111 : OUT <= 0;  //155 / 239 = 0
    16'b10011011_11110000 : OUT <= 0;  //155 / 240 = 0
    16'b10011011_11110001 : OUT <= 0;  //155 / 241 = 0
    16'b10011011_11110010 : OUT <= 0;  //155 / 242 = 0
    16'b10011011_11110011 : OUT <= 0;  //155 / 243 = 0
    16'b10011011_11110100 : OUT <= 0;  //155 / 244 = 0
    16'b10011011_11110101 : OUT <= 0;  //155 / 245 = 0
    16'b10011011_11110110 : OUT <= 0;  //155 / 246 = 0
    16'b10011011_11110111 : OUT <= 0;  //155 / 247 = 0
    16'b10011011_11111000 : OUT <= 0;  //155 / 248 = 0
    16'b10011011_11111001 : OUT <= 0;  //155 / 249 = 0
    16'b10011011_11111010 : OUT <= 0;  //155 / 250 = 0
    16'b10011011_11111011 : OUT <= 0;  //155 / 251 = 0
    16'b10011011_11111100 : OUT <= 0;  //155 / 252 = 0
    16'b10011011_11111101 : OUT <= 0;  //155 / 253 = 0
    16'b10011011_11111110 : OUT <= 0;  //155 / 254 = 0
    16'b10011011_11111111 : OUT <= 0;  //155 / 255 = 0
    16'b10011100_00000000 : OUT <= 0;  //156 / 0 = 0
    16'b10011100_00000001 : OUT <= 156;  //156 / 1 = 156
    16'b10011100_00000010 : OUT <= 78;  //156 / 2 = 78
    16'b10011100_00000011 : OUT <= 52;  //156 / 3 = 52
    16'b10011100_00000100 : OUT <= 39;  //156 / 4 = 39
    16'b10011100_00000101 : OUT <= 31;  //156 / 5 = 31
    16'b10011100_00000110 : OUT <= 26;  //156 / 6 = 26
    16'b10011100_00000111 : OUT <= 22;  //156 / 7 = 22
    16'b10011100_00001000 : OUT <= 19;  //156 / 8 = 19
    16'b10011100_00001001 : OUT <= 17;  //156 / 9 = 17
    16'b10011100_00001010 : OUT <= 15;  //156 / 10 = 15
    16'b10011100_00001011 : OUT <= 14;  //156 / 11 = 14
    16'b10011100_00001100 : OUT <= 13;  //156 / 12 = 13
    16'b10011100_00001101 : OUT <= 12;  //156 / 13 = 12
    16'b10011100_00001110 : OUT <= 11;  //156 / 14 = 11
    16'b10011100_00001111 : OUT <= 10;  //156 / 15 = 10
    16'b10011100_00010000 : OUT <= 9;  //156 / 16 = 9
    16'b10011100_00010001 : OUT <= 9;  //156 / 17 = 9
    16'b10011100_00010010 : OUT <= 8;  //156 / 18 = 8
    16'b10011100_00010011 : OUT <= 8;  //156 / 19 = 8
    16'b10011100_00010100 : OUT <= 7;  //156 / 20 = 7
    16'b10011100_00010101 : OUT <= 7;  //156 / 21 = 7
    16'b10011100_00010110 : OUT <= 7;  //156 / 22 = 7
    16'b10011100_00010111 : OUT <= 6;  //156 / 23 = 6
    16'b10011100_00011000 : OUT <= 6;  //156 / 24 = 6
    16'b10011100_00011001 : OUT <= 6;  //156 / 25 = 6
    16'b10011100_00011010 : OUT <= 6;  //156 / 26 = 6
    16'b10011100_00011011 : OUT <= 5;  //156 / 27 = 5
    16'b10011100_00011100 : OUT <= 5;  //156 / 28 = 5
    16'b10011100_00011101 : OUT <= 5;  //156 / 29 = 5
    16'b10011100_00011110 : OUT <= 5;  //156 / 30 = 5
    16'b10011100_00011111 : OUT <= 5;  //156 / 31 = 5
    16'b10011100_00100000 : OUT <= 4;  //156 / 32 = 4
    16'b10011100_00100001 : OUT <= 4;  //156 / 33 = 4
    16'b10011100_00100010 : OUT <= 4;  //156 / 34 = 4
    16'b10011100_00100011 : OUT <= 4;  //156 / 35 = 4
    16'b10011100_00100100 : OUT <= 4;  //156 / 36 = 4
    16'b10011100_00100101 : OUT <= 4;  //156 / 37 = 4
    16'b10011100_00100110 : OUT <= 4;  //156 / 38 = 4
    16'b10011100_00100111 : OUT <= 4;  //156 / 39 = 4
    16'b10011100_00101000 : OUT <= 3;  //156 / 40 = 3
    16'b10011100_00101001 : OUT <= 3;  //156 / 41 = 3
    16'b10011100_00101010 : OUT <= 3;  //156 / 42 = 3
    16'b10011100_00101011 : OUT <= 3;  //156 / 43 = 3
    16'b10011100_00101100 : OUT <= 3;  //156 / 44 = 3
    16'b10011100_00101101 : OUT <= 3;  //156 / 45 = 3
    16'b10011100_00101110 : OUT <= 3;  //156 / 46 = 3
    16'b10011100_00101111 : OUT <= 3;  //156 / 47 = 3
    16'b10011100_00110000 : OUT <= 3;  //156 / 48 = 3
    16'b10011100_00110001 : OUT <= 3;  //156 / 49 = 3
    16'b10011100_00110010 : OUT <= 3;  //156 / 50 = 3
    16'b10011100_00110011 : OUT <= 3;  //156 / 51 = 3
    16'b10011100_00110100 : OUT <= 3;  //156 / 52 = 3
    16'b10011100_00110101 : OUT <= 2;  //156 / 53 = 2
    16'b10011100_00110110 : OUT <= 2;  //156 / 54 = 2
    16'b10011100_00110111 : OUT <= 2;  //156 / 55 = 2
    16'b10011100_00111000 : OUT <= 2;  //156 / 56 = 2
    16'b10011100_00111001 : OUT <= 2;  //156 / 57 = 2
    16'b10011100_00111010 : OUT <= 2;  //156 / 58 = 2
    16'b10011100_00111011 : OUT <= 2;  //156 / 59 = 2
    16'b10011100_00111100 : OUT <= 2;  //156 / 60 = 2
    16'b10011100_00111101 : OUT <= 2;  //156 / 61 = 2
    16'b10011100_00111110 : OUT <= 2;  //156 / 62 = 2
    16'b10011100_00111111 : OUT <= 2;  //156 / 63 = 2
    16'b10011100_01000000 : OUT <= 2;  //156 / 64 = 2
    16'b10011100_01000001 : OUT <= 2;  //156 / 65 = 2
    16'b10011100_01000010 : OUT <= 2;  //156 / 66 = 2
    16'b10011100_01000011 : OUT <= 2;  //156 / 67 = 2
    16'b10011100_01000100 : OUT <= 2;  //156 / 68 = 2
    16'b10011100_01000101 : OUT <= 2;  //156 / 69 = 2
    16'b10011100_01000110 : OUT <= 2;  //156 / 70 = 2
    16'b10011100_01000111 : OUT <= 2;  //156 / 71 = 2
    16'b10011100_01001000 : OUT <= 2;  //156 / 72 = 2
    16'b10011100_01001001 : OUT <= 2;  //156 / 73 = 2
    16'b10011100_01001010 : OUT <= 2;  //156 / 74 = 2
    16'b10011100_01001011 : OUT <= 2;  //156 / 75 = 2
    16'b10011100_01001100 : OUT <= 2;  //156 / 76 = 2
    16'b10011100_01001101 : OUT <= 2;  //156 / 77 = 2
    16'b10011100_01001110 : OUT <= 2;  //156 / 78 = 2
    16'b10011100_01001111 : OUT <= 1;  //156 / 79 = 1
    16'b10011100_01010000 : OUT <= 1;  //156 / 80 = 1
    16'b10011100_01010001 : OUT <= 1;  //156 / 81 = 1
    16'b10011100_01010010 : OUT <= 1;  //156 / 82 = 1
    16'b10011100_01010011 : OUT <= 1;  //156 / 83 = 1
    16'b10011100_01010100 : OUT <= 1;  //156 / 84 = 1
    16'b10011100_01010101 : OUT <= 1;  //156 / 85 = 1
    16'b10011100_01010110 : OUT <= 1;  //156 / 86 = 1
    16'b10011100_01010111 : OUT <= 1;  //156 / 87 = 1
    16'b10011100_01011000 : OUT <= 1;  //156 / 88 = 1
    16'b10011100_01011001 : OUT <= 1;  //156 / 89 = 1
    16'b10011100_01011010 : OUT <= 1;  //156 / 90 = 1
    16'b10011100_01011011 : OUT <= 1;  //156 / 91 = 1
    16'b10011100_01011100 : OUT <= 1;  //156 / 92 = 1
    16'b10011100_01011101 : OUT <= 1;  //156 / 93 = 1
    16'b10011100_01011110 : OUT <= 1;  //156 / 94 = 1
    16'b10011100_01011111 : OUT <= 1;  //156 / 95 = 1
    16'b10011100_01100000 : OUT <= 1;  //156 / 96 = 1
    16'b10011100_01100001 : OUT <= 1;  //156 / 97 = 1
    16'b10011100_01100010 : OUT <= 1;  //156 / 98 = 1
    16'b10011100_01100011 : OUT <= 1;  //156 / 99 = 1
    16'b10011100_01100100 : OUT <= 1;  //156 / 100 = 1
    16'b10011100_01100101 : OUT <= 1;  //156 / 101 = 1
    16'b10011100_01100110 : OUT <= 1;  //156 / 102 = 1
    16'b10011100_01100111 : OUT <= 1;  //156 / 103 = 1
    16'b10011100_01101000 : OUT <= 1;  //156 / 104 = 1
    16'b10011100_01101001 : OUT <= 1;  //156 / 105 = 1
    16'b10011100_01101010 : OUT <= 1;  //156 / 106 = 1
    16'b10011100_01101011 : OUT <= 1;  //156 / 107 = 1
    16'b10011100_01101100 : OUT <= 1;  //156 / 108 = 1
    16'b10011100_01101101 : OUT <= 1;  //156 / 109 = 1
    16'b10011100_01101110 : OUT <= 1;  //156 / 110 = 1
    16'b10011100_01101111 : OUT <= 1;  //156 / 111 = 1
    16'b10011100_01110000 : OUT <= 1;  //156 / 112 = 1
    16'b10011100_01110001 : OUT <= 1;  //156 / 113 = 1
    16'b10011100_01110010 : OUT <= 1;  //156 / 114 = 1
    16'b10011100_01110011 : OUT <= 1;  //156 / 115 = 1
    16'b10011100_01110100 : OUT <= 1;  //156 / 116 = 1
    16'b10011100_01110101 : OUT <= 1;  //156 / 117 = 1
    16'b10011100_01110110 : OUT <= 1;  //156 / 118 = 1
    16'b10011100_01110111 : OUT <= 1;  //156 / 119 = 1
    16'b10011100_01111000 : OUT <= 1;  //156 / 120 = 1
    16'b10011100_01111001 : OUT <= 1;  //156 / 121 = 1
    16'b10011100_01111010 : OUT <= 1;  //156 / 122 = 1
    16'b10011100_01111011 : OUT <= 1;  //156 / 123 = 1
    16'b10011100_01111100 : OUT <= 1;  //156 / 124 = 1
    16'b10011100_01111101 : OUT <= 1;  //156 / 125 = 1
    16'b10011100_01111110 : OUT <= 1;  //156 / 126 = 1
    16'b10011100_01111111 : OUT <= 1;  //156 / 127 = 1
    16'b10011100_10000000 : OUT <= 1;  //156 / 128 = 1
    16'b10011100_10000001 : OUT <= 1;  //156 / 129 = 1
    16'b10011100_10000010 : OUT <= 1;  //156 / 130 = 1
    16'b10011100_10000011 : OUT <= 1;  //156 / 131 = 1
    16'b10011100_10000100 : OUT <= 1;  //156 / 132 = 1
    16'b10011100_10000101 : OUT <= 1;  //156 / 133 = 1
    16'b10011100_10000110 : OUT <= 1;  //156 / 134 = 1
    16'b10011100_10000111 : OUT <= 1;  //156 / 135 = 1
    16'b10011100_10001000 : OUT <= 1;  //156 / 136 = 1
    16'b10011100_10001001 : OUT <= 1;  //156 / 137 = 1
    16'b10011100_10001010 : OUT <= 1;  //156 / 138 = 1
    16'b10011100_10001011 : OUT <= 1;  //156 / 139 = 1
    16'b10011100_10001100 : OUT <= 1;  //156 / 140 = 1
    16'b10011100_10001101 : OUT <= 1;  //156 / 141 = 1
    16'b10011100_10001110 : OUT <= 1;  //156 / 142 = 1
    16'b10011100_10001111 : OUT <= 1;  //156 / 143 = 1
    16'b10011100_10010000 : OUT <= 1;  //156 / 144 = 1
    16'b10011100_10010001 : OUT <= 1;  //156 / 145 = 1
    16'b10011100_10010010 : OUT <= 1;  //156 / 146 = 1
    16'b10011100_10010011 : OUT <= 1;  //156 / 147 = 1
    16'b10011100_10010100 : OUT <= 1;  //156 / 148 = 1
    16'b10011100_10010101 : OUT <= 1;  //156 / 149 = 1
    16'b10011100_10010110 : OUT <= 1;  //156 / 150 = 1
    16'b10011100_10010111 : OUT <= 1;  //156 / 151 = 1
    16'b10011100_10011000 : OUT <= 1;  //156 / 152 = 1
    16'b10011100_10011001 : OUT <= 1;  //156 / 153 = 1
    16'b10011100_10011010 : OUT <= 1;  //156 / 154 = 1
    16'b10011100_10011011 : OUT <= 1;  //156 / 155 = 1
    16'b10011100_10011100 : OUT <= 1;  //156 / 156 = 1
    16'b10011100_10011101 : OUT <= 0;  //156 / 157 = 0
    16'b10011100_10011110 : OUT <= 0;  //156 / 158 = 0
    16'b10011100_10011111 : OUT <= 0;  //156 / 159 = 0
    16'b10011100_10100000 : OUT <= 0;  //156 / 160 = 0
    16'b10011100_10100001 : OUT <= 0;  //156 / 161 = 0
    16'b10011100_10100010 : OUT <= 0;  //156 / 162 = 0
    16'b10011100_10100011 : OUT <= 0;  //156 / 163 = 0
    16'b10011100_10100100 : OUT <= 0;  //156 / 164 = 0
    16'b10011100_10100101 : OUT <= 0;  //156 / 165 = 0
    16'b10011100_10100110 : OUT <= 0;  //156 / 166 = 0
    16'b10011100_10100111 : OUT <= 0;  //156 / 167 = 0
    16'b10011100_10101000 : OUT <= 0;  //156 / 168 = 0
    16'b10011100_10101001 : OUT <= 0;  //156 / 169 = 0
    16'b10011100_10101010 : OUT <= 0;  //156 / 170 = 0
    16'b10011100_10101011 : OUT <= 0;  //156 / 171 = 0
    16'b10011100_10101100 : OUT <= 0;  //156 / 172 = 0
    16'b10011100_10101101 : OUT <= 0;  //156 / 173 = 0
    16'b10011100_10101110 : OUT <= 0;  //156 / 174 = 0
    16'b10011100_10101111 : OUT <= 0;  //156 / 175 = 0
    16'b10011100_10110000 : OUT <= 0;  //156 / 176 = 0
    16'b10011100_10110001 : OUT <= 0;  //156 / 177 = 0
    16'b10011100_10110010 : OUT <= 0;  //156 / 178 = 0
    16'b10011100_10110011 : OUT <= 0;  //156 / 179 = 0
    16'b10011100_10110100 : OUT <= 0;  //156 / 180 = 0
    16'b10011100_10110101 : OUT <= 0;  //156 / 181 = 0
    16'b10011100_10110110 : OUT <= 0;  //156 / 182 = 0
    16'b10011100_10110111 : OUT <= 0;  //156 / 183 = 0
    16'b10011100_10111000 : OUT <= 0;  //156 / 184 = 0
    16'b10011100_10111001 : OUT <= 0;  //156 / 185 = 0
    16'b10011100_10111010 : OUT <= 0;  //156 / 186 = 0
    16'b10011100_10111011 : OUT <= 0;  //156 / 187 = 0
    16'b10011100_10111100 : OUT <= 0;  //156 / 188 = 0
    16'b10011100_10111101 : OUT <= 0;  //156 / 189 = 0
    16'b10011100_10111110 : OUT <= 0;  //156 / 190 = 0
    16'b10011100_10111111 : OUT <= 0;  //156 / 191 = 0
    16'b10011100_11000000 : OUT <= 0;  //156 / 192 = 0
    16'b10011100_11000001 : OUT <= 0;  //156 / 193 = 0
    16'b10011100_11000010 : OUT <= 0;  //156 / 194 = 0
    16'b10011100_11000011 : OUT <= 0;  //156 / 195 = 0
    16'b10011100_11000100 : OUT <= 0;  //156 / 196 = 0
    16'b10011100_11000101 : OUT <= 0;  //156 / 197 = 0
    16'b10011100_11000110 : OUT <= 0;  //156 / 198 = 0
    16'b10011100_11000111 : OUT <= 0;  //156 / 199 = 0
    16'b10011100_11001000 : OUT <= 0;  //156 / 200 = 0
    16'b10011100_11001001 : OUT <= 0;  //156 / 201 = 0
    16'b10011100_11001010 : OUT <= 0;  //156 / 202 = 0
    16'b10011100_11001011 : OUT <= 0;  //156 / 203 = 0
    16'b10011100_11001100 : OUT <= 0;  //156 / 204 = 0
    16'b10011100_11001101 : OUT <= 0;  //156 / 205 = 0
    16'b10011100_11001110 : OUT <= 0;  //156 / 206 = 0
    16'b10011100_11001111 : OUT <= 0;  //156 / 207 = 0
    16'b10011100_11010000 : OUT <= 0;  //156 / 208 = 0
    16'b10011100_11010001 : OUT <= 0;  //156 / 209 = 0
    16'b10011100_11010010 : OUT <= 0;  //156 / 210 = 0
    16'b10011100_11010011 : OUT <= 0;  //156 / 211 = 0
    16'b10011100_11010100 : OUT <= 0;  //156 / 212 = 0
    16'b10011100_11010101 : OUT <= 0;  //156 / 213 = 0
    16'b10011100_11010110 : OUT <= 0;  //156 / 214 = 0
    16'b10011100_11010111 : OUT <= 0;  //156 / 215 = 0
    16'b10011100_11011000 : OUT <= 0;  //156 / 216 = 0
    16'b10011100_11011001 : OUT <= 0;  //156 / 217 = 0
    16'b10011100_11011010 : OUT <= 0;  //156 / 218 = 0
    16'b10011100_11011011 : OUT <= 0;  //156 / 219 = 0
    16'b10011100_11011100 : OUT <= 0;  //156 / 220 = 0
    16'b10011100_11011101 : OUT <= 0;  //156 / 221 = 0
    16'b10011100_11011110 : OUT <= 0;  //156 / 222 = 0
    16'b10011100_11011111 : OUT <= 0;  //156 / 223 = 0
    16'b10011100_11100000 : OUT <= 0;  //156 / 224 = 0
    16'b10011100_11100001 : OUT <= 0;  //156 / 225 = 0
    16'b10011100_11100010 : OUT <= 0;  //156 / 226 = 0
    16'b10011100_11100011 : OUT <= 0;  //156 / 227 = 0
    16'b10011100_11100100 : OUT <= 0;  //156 / 228 = 0
    16'b10011100_11100101 : OUT <= 0;  //156 / 229 = 0
    16'b10011100_11100110 : OUT <= 0;  //156 / 230 = 0
    16'b10011100_11100111 : OUT <= 0;  //156 / 231 = 0
    16'b10011100_11101000 : OUT <= 0;  //156 / 232 = 0
    16'b10011100_11101001 : OUT <= 0;  //156 / 233 = 0
    16'b10011100_11101010 : OUT <= 0;  //156 / 234 = 0
    16'b10011100_11101011 : OUT <= 0;  //156 / 235 = 0
    16'b10011100_11101100 : OUT <= 0;  //156 / 236 = 0
    16'b10011100_11101101 : OUT <= 0;  //156 / 237 = 0
    16'b10011100_11101110 : OUT <= 0;  //156 / 238 = 0
    16'b10011100_11101111 : OUT <= 0;  //156 / 239 = 0
    16'b10011100_11110000 : OUT <= 0;  //156 / 240 = 0
    16'b10011100_11110001 : OUT <= 0;  //156 / 241 = 0
    16'b10011100_11110010 : OUT <= 0;  //156 / 242 = 0
    16'b10011100_11110011 : OUT <= 0;  //156 / 243 = 0
    16'b10011100_11110100 : OUT <= 0;  //156 / 244 = 0
    16'b10011100_11110101 : OUT <= 0;  //156 / 245 = 0
    16'b10011100_11110110 : OUT <= 0;  //156 / 246 = 0
    16'b10011100_11110111 : OUT <= 0;  //156 / 247 = 0
    16'b10011100_11111000 : OUT <= 0;  //156 / 248 = 0
    16'b10011100_11111001 : OUT <= 0;  //156 / 249 = 0
    16'b10011100_11111010 : OUT <= 0;  //156 / 250 = 0
    16'b10011100_11111011 : OUT <= 0;  //156 / 251 = 0
    16'b10011100_11111100 : OUT <= 0;  //156 / 252 = 0
    16'b10011100_11111101 : OUT <= 0;  //156 / 253 = 0
    16'b10011100_11111110 : OUT <= 0;  //156 / 254 = 0
    16'b10011100_11111111 : OUT <= 0;  //156 / 255 = 0
    16'b10011101_00000000 : OUT <= 0;  //157 / 0 = 0
    16'b10011101_00000001 : OUT <= 157;  //157 / 1 = 157
    16'b10011101_00000010 : OUT <= 78;  //157 / 2 = 78
    16'b10011101_00000011 : OUT <= 52;  //157 / 3 = 52
    16'b10011101_00000100 : OUT <= 39;  //157 / 4 = 39
    16'b10011101_00000101 : OUT <= 31;  //157 / 5 = 31
    16'b10011101_00000110 : OUT <= 26;  //157 / 6 = 26
    16'b10011101_00000111 : OUT <= 22;  //157 / 7 = 22
    16'b10011101_00001000 : OUT <= 19;  //157 / 8 = 19
    16'b10011101_00001001 : OUT <= 17;  //157 / 9 = 17
    16'b10011101_00001010 : OUT <= 15;  //157 / 10 = 15
    16'b10011101_00001011 : OUT <= 14;  //157 / 11 = 14
    16'b10011101_00001100 : OUT <= 13;  //157 / 12 = 13
    16'b10011101_00001101 : OUT <= 12;  //157 / 13 = 12
    16'b10011101_00001110 : OUT <= 11;  //157 / 14 = 11
    16'b10011101_00001111 : OUT <= 10;  //157 / 15 = 10
    16'b10011101_00010000 : OUT <= 9;  //157 / 16 = 9
    16'b10011101_00010001 : OUT <= 9;  //157 / 17 = 9
    16'b10011101_00010010 : OUT <= 8;  //157 / 18 = 8
    16'b10011101_00010011 : OUT <= 8;  //157 / 19 = 8
    16'b10011101_00010100 : OUT <= 7;  //157 / 20 = 7
    16'b10011101_00010101 : OUT <= 7;  //157 / 21 = 7
    16'b10011101_00010110 : OUT <= 7;  //157 / 22 = 7
    16'b10011101_00010111 : OUT <= 6;  //157 / 23 = 6
    16'b10011101_00011000 : OUT <= 6;  //157 / 24 = 6
    16'b10011101_00011001 : OUT <= 6;  //157 / 25 = 6
    16'b10011101_00011010 : OUT <= 6;  //157 / 26 = 6
    16'b10011101_00011011 : OUT <= 5;  //157 / 27 = 5
    16'b10011101_00011100 : OUT <= 5;  //157 / 28 = 5
    16'b10011101_00011101 : OUT <= 5;  //157 / 29 = 5
    16'b10011101_00011110 : OUT <= 5;  //157 / 30 = 5
    16'b10011101_00011111 : OUT <= 5;  //157 / 31 = 5
    16'b10011101_00100000 : OUT <= 4;  //157 / 32 = 4
    16'b10011101_00100001 : OUT <= 4;  //157 / 33 = 4
    16'b10011101_00100010 : OUT <= 4;  //157 / 34 = 4
    16'b10011101_00100011 : OUT <= 4;  //157 / 35 = 4
    16'b10011101_00100100 : OUT <= 4;  //157 / 36 = 4
    16'b10011101_00100101 : OUT <= 4;  //157 / 37 = 4
    16'b10011101_00100110 : OUT <= 4;  //157 / 38 = 4
    16'b10011101_00100111 : OUT <= 4;  //157 / 39 = 4
    16'b10011101_00101000 : OUT <= 3;  //157 / 40 = 3
    16'b10011101_00101001 : OUT <= 3;  //157 / 41 = 3
    16'b10011101_00101010 : OUT <= 3;  //157 / 42 = 3
    16'b10011101_00101011 : OUT <= 3;  //157 / 43 = 3
    16'b10011101_00101100 : OUT <= 3;  //157 / 44 = 3
    16'b10011101_00101101 : OUT <= 3;  //157 / 45 = 3
    16'b10011101_00101110 : OUT <= 3;  //157 / 46 = 3
    16'b10011101_00101111 : OUT <= 3;  //157 / 47 = 3
    16'b10011101_00110000 : OUT <= 3;  //157 / 48 = 3
    16'b10011101_00110001 : OUT <= 3;  //157 / 49 = 3
    16'b10011101_00110010 : OUT <= 3;  //157 / 50 = 3
    16'b10011101_00110011 : OUT <= 3;  //157 / 51 = 3
    16'b10011101_00110100 : OUT <= 3;  //157 / 52 = 3
    16'b10011101_00110101 : OUT <= 2;  //157 / 53 = 2
    16'b10011101_00110110 : OUT <= 2;  //157 / 54 = 2
    16'b10011101_00110111 : OUT <= 2;  //157 / 55 = 2
    16'b10011101_00111000 : OUT <= 2;  //157 / 56 = 2
    16'b10011101_00111001 : OUT <= 2;  //157 / 57 = 2
    16'b10011101_00111010 : OUT <= 2;  //157 / 58 = 2
    16'b10011101_00111011 : OUT <= 2;  //157 / 59 = 2
    16'b10011101_00111100 : OUT <= 2;  //157 / 60 = 2
    16'b10011101_00111101 : OUT <= 2;  //157 / 61 = 2
    16'b10011101_00111110 : OUT <= 2;  //157 / 62 = 2
    16'b10011101_00111111 : OUT <= 2;  //157 / 63 = 2
    16'b10011101_01000000 : OUT <= 2;  //157 / 64 = 2
    16'b10011101_01000001 : OUT <= 2;  //157 / 65 = 2
    16'b10011101_01000010 : OUT <= 2;  //157 / 66 = 2
    16'b10011101_01000011 : OUT <= 2;  //157 / 67 = 2
    16'b10011101_01000100 : OUT <= 2;  //157 / 68 = 2
    16'b10011101_01000101 : OUT <= 2;  //157 / 69 = 2
    16'b10011101_01000110 : OUT <= 2;  //157 / 70 = 2
    16'b10011101_01000111 : OUT <= 2;  //157 / 71 = 2
    16'b10011101_01001000 : OUT <= 2;  //157 / 72 = 2
    16'b10011101_01001001 : OUT <= 2;  //157 / 73 = 2
    16'b10011101_01001010 : OUT <= 2;  //157 / 74 = 2
    16'b10011101_01001011 : OUT <= 2;  //157 / 75 = 2
    16'b10011101_01001100 : OUT <= 2;  //157 / 76 = 2
    16'b10011101_01001101 : OUT <= 2;  //157 / 77 = 2
    16'b10011101_01001110 : OUT <= 2;  //157 / 78 = 2
    16'b10011101_01001111 : OUT <= 1;  //157 / 79 = 1
    16'b10011101_01010000 : OUT <= 1;  //157 / 80 = 1
    16'b10011101_01010001 : OUT <= 1;  //157 / 81 = 1
    16'b10011101_01010010 : OUT <= 1;  //157 / 82 = 1
    16'b10011101_01010011 : OUT <= 1;  //157 / 83 = 1
    16'b10011101_01010100 : OUT <= 1;  //157 / 84 = 1
    16'b10011101_01010101 : OUT <= 1;  //157 / 85 = 1
    16'b10011101_01010110 : OUT <= 1;  //157 / 86 = 1
    16'b10011101_01010111 : OUT <= 1;  //157 / 87 = 1
    16'b10011101_01011000 : OUT <= 1;  //157 / 88 = 1
    16'b10011101_01011001 : OUT <= 1;  //157 / 89 = 1
    16'b10011101_01011010 : OUT <= 1;  //157 / 90 = 1
    16'b10011101_01011011 : OUT <= 1;  //157 / 91 = 1
    16'b10011101_01011100 : OUT <= 1;  //157 / 92 = 1
    16'b10011101_01011101 : OUT <= 1;  //157 / 93 = 1
    16'b10011101_01011110 : OUT <= 1;  //157 / 94 = 1
    16'b10011101_01011111 : OUT <= 1;  //157 / 95 = 1
    16'b10011101_01100000 : OUT <= 1;  //157 / 96 = 1
    16'b10011101_01100001 : OUT <= 1;  //157 / 97 = 1
    16'b10011101_01100010 : OUT <= 1;  //157 / 98 = 1
    16'b10011101_01100011 : OUT <= 1;  //157 / 99 = 1
    16'b10011101_01100100 : OUT <= 1;  //157 / 100 = 1
    16'b10011101_01100101 : OUT <= 1;  //157 / 101 = 1
    16'b10011101_01100110 : OUT <= 1;  //157 / 102 = 1
    16'b10011101_01100111 : OUT <= 1;  //157 / 103 = 1
    16'b10011101_01101000 : OUT <= 1;  //157 / 104 = 1
    16'b10011101_01101001 : OUT <= 1;  //157 / 105 = 1
    16'b10011101_01101010 : OUT <= 1;  //157 / 106 = 1
    16'b10011101_01101011 : OUT <= 1;  //157 / 107 = 1
    16'b10011101_01101100 : OUT <= 1;  //157 / 108 = 1
    16'b10011101_01101101 : OUT <= 1;  //157 / 109 = 1
    16'b10011101_01101110 : OUT <= 1;  //157 / 110 = 1
    16'b10011101_01101111 : OUT <= 1;  //157 / 111 = 1
    16'b10011101_01110000 : OUT <= 1;  //157 / 112 = 1
    16'b10011101_01110001 : OUT <= 1;  //157 / 113 = 1
    16'b10011101_01110010 : OUT <= 1;  //157 / 114 = 1
    16'b10011101_01110011 : OUT <= 1;  //157 / 115 = 1
    16'b10011101_01110100 : OUT <= 1;  //157 / 116 = 1
    16'b10011101_01110101 : OUT <= 1;  //157 / 117 = 1
    16'b10011101_01110110 : OUT <= 1;  //157 / 118 = 1
    16'b10011101_01110111 : OUT <= 1;  //157 / 119 = 1
    16'b10011101_01111000 : OUT <= 1;  //157 / 120 = 1
    16'b10011101_01111001 : OUT <= 1;  //157 / 121 = 1
    16'b10011101_01111010 : OUT <= 1;  //157 / 122 = 1
    16'b10011101_01111011 : OUT <= 1;  //157 / 123 = 1
    16'b10011101_01111100 : OUT <= 1;  //157 / 124 = 1
    16'b10011101_01111101 : OUT <= 1;  //157 / 125 = 1
    16'b10011101_01111110 : OUT <= 1;  //157 / 126 = 1
    16'b10011101_01111111 : OUT <= 1;  //157 / 127 = 1
    16'b10011101_10000000 : OUT <= 1;  //157 / 128 = 1
    16'b10011101_10000001 : OUT <= 1;  //157 / 129 = 1
    16'b10011101_10000010 : OUT <= 1;  //157 / 130 = 1
    16'b10011101_10000011 : OUT <= 1;  //157 / 131 = 1
    16'b10011101_10000100 : OUT <= 1;  //157 / 132 = 1
    16'b10011101_10000101 : OUT <= 1;  //157 / 133 = 1
    16'b10011101_10000110 : OUT <= 1;  //157 / 134 = 1
    16'b10011101_10000111 : OUT <= 1;  //157 / 135 = 1
    16'b10011101_10001000 : OUT <= 1;  //157 / 136 = 1
    16'b10011101_10001001 : OUT <= 1;  //157 / 137 = 1
    16'b10011101_10001010 : OUT <= 1;  //157 / 138 = 1
    16'b10011101_10001011 : OUT <= 1;  //157 / 139 = 1
    16'b10011101_10001100 : OUT <= 1;  //157 / 140 = 1
    16'b10011101_10001101 : OUT <= 1;  //157 / 141 = 1
    16'b10011101_10001110 : OUT <= 1;  //157 / 142 = 1
    16'b10011101_10001111 : OUT <= 1;  //157 / 143 = 1
    16'b10011101_10010000 : OUT <= 1;  //157 / 144 = 1
    16'b10011101_10010001 : OUT <= 1;  //157 / 145 = 1
    16'b10011101_10010010 : OUT <= 1;  //157 / 146 = 1
    16'b10011101_10010011 : OUT <= 1;  //157 / 147 = 1
    16'b10011101_10010100 : OUT <= 1;  //157 / 148 = 1
    16'b10011101_10010101 : OUT <= 1;  //157 / 149 = 1
    16'b10011101_10010110 : OUT <= 1;  //157 / 150 = 1
    16'b10011101_10010111 : OUT <= 1;  //157 / 151 = 1
    16'b10011101_10011000 : OUT <= 1;  //157 / 152 = 1
    16'b10011101_10011001 : OUT <= 1;  //157 / 153 = 1
    16'b10011101_10011010 : OUT <= 1;  //157 / 154 = 1
    16'b10011101_10011011 : OUT <= 1;  //157 / 155 = 1
    16'b10011101_10011100 : OUT <= 1;  //157 / 156 = 1
    16'b10011101_10011101 : OUT <= 1;  //157 / 157 = 1
    16'b10011101_10011110 : OUT <= 0;  //157 / 158 = 0
    16'b10011101_10011111 : OUT <= 0;  //157 / 159 = 0
    16'b10011101_10100000 : OUT <= 0;  //157 / 160 = 0
    16'b10011101_10100001 : OUT <= 0;  //157 / 161 = 0
    16'b10011101_10100010 : OUT <= 0;  //157 / 162 = 0
    16'b10011101_10100011 : OUT <= 0;  //157 / 163 = 0
    16'b10011101_10100100 : OUT <= 0;  //157 / 164 = 0
    16'b10011101_10100101 : OUT <= 0;  //157 / 165 = 0
    16'b10011101_10100110 : OUT <= 0;  //157 / 166 = 0
    16'b10011101_10100111 : OUT <= 0;  //157 / 167 = 0
    16'b10011101_10101000 : OUT <= 0;  //157 / 168 = 0
    16'b10011101_10101001 : OUT <= 0;  //157 / 169 = 0
    16'b10011101_10101010 : OUT <= 0;  //157 / 170 = 0
    16'b10011101_10101011 : OUT <= 0;  //157 / 171 = 0
    16'b10011101_10101100 : OUT <= 0;  //157 / 172 = 0
    16'b10011101_10101101 : OUT <= 0;  //157 / 173 = 0
    16'b10011101_10101110 : OUT <= 0;  //157 / 174 = 0
    16'b10011101_10101111 : OUT <= 0;  //157 / 175 = 0
    16'b10011101_10110000 : OUT <= 0;  //157 / 176 = 0
    16'b10011101_10110001 : OUT <= 0;  //157 / 177 = 0
    16'b10011101_10110010 : OUT <= 0;  //157 / 178 = 0
    16'b10011101_10110011 : OUT <= 0;  //157 / 179 = 0
    16'b10011101_10110100 : OUT <= 0;  //157 / 180 = 0
    16'b10011101_10110101 : OUT <= 0;  //157 / 181 = 0
    16'b10011101_10110110 : OUT <= 0;  //157 / 182 = 0
    16'b10011101_10110111 : OUT <= 0;  //157 / 183 = 0
    16'b10011101_10111000 : OUT <= 0;  //157 / 184 = 0
    16'b10011101_10111001 : OUT <= 0;  //157 / 185 = 0
    16'b10011101_10111010 : OUT <= 0;  //157 / 186 = 0
    16'b10011101_10111011 : OUT <= 0;  //157 / 187 = 0
    16'b10011101_10111100 : OUT <= 0;  //157 / 188 = 0
    16'b10011101_10111101 : OUT <= 0;  //157 / 189 = 0
    16'b10011101_10111110 : OUT <= 0;  //157 / 190 = 0
    16'b10011101_10111111 : OUT <= 0;  //157 / 191 = 0
    16'b10011101_11000000 : OUT <= 0;  //157 / 192 = 0
    16'b10011101_11000001 : OUT <= 0;  //157 / 193 = 0
    16'b10011101_11000010 : OUT <= 0;  //157 / 194 = 0
    16'b10011101_11000011 : OUT <= 0;  //157 / 195 = 0
    16'b10011101_11000100 : OUT <= 0;  //157 / 196 = 0
    16'b10011101_11000101 : OUT <= 0;  //157 / 197 = 0
    16'b10011101_11000110 : OUT <= 0;  //157 / 198 = 0
    16'b10011101_11000111 : OUT <= 0;  //157 / 199 = 0
    16'b10011101_11001000 : OUT <= 0;  //157 / 200 = 0
    16'b10011101_11001001 : OUT <= 0;  //157 / 201 = 0
    16'b10011101_11001010 : OUT <= 0;  //157 / 202 = 0
    16'b10011101_11001011 : OUT <= 0;  //157 / 203 = 0
    16'b10011101_11001100 : OUT <= 0;  //157 / 204 = 0
    16'b10011101_11001101 : OUT <= 0;  //157 / 205 = 0
    16'b10011101_11001110 : OUT <= 0;  //157 / 206 = 0
    16'b10011101_11001111 : OUT <= 0;  //157 / 207 = 0
    16'b10011101_11010000 : OUT <= 0;  //157 / 208 = 0
    16'b10011101_11010001 : OUT <= 0;  //157 / 209 = 0
    16'b10011101_11010010 : OUT <= 0;  //157 / 210 = 0
    16'b10011101_11010011 : OUT <= 0;  //157 / 211 = 0
    16'b10011101_11010100 : OUT <= 0;  //157 / 212 = 0
    16'b10011101_11010101 : OUT <= 0;  //157 / 213 = 0
    16'b10011101_11010110 : OUT <= 0;  //157 / 214 = 0
    16'b10011101_11010111 : OUT <= 0;  //157 / 215 = 0
    16'b10011101_11011000 : OUT <= 0;  //157 / 216 = 0
    16'b10011101_11011001 : OUT <= 0;  //157 / 217 = 0
    16'b10011101_11011010 : OUT <= 0;  //157 / 218 = 0
    16'b10011101_11011011 : OUT <= 0;  //157 / 219 = 0
    16'b10011101_11011100 : OUT <= 0;  //157 / 220 = 0
    16'b10011101_11011101 : OUT <= 0;  //157 / 221 = 0
    16'b10011101_11011110 : OUT <= 0;  //157 / 222 = 0
    16'b10011101_11011111 : OUT <= 0;  //157 / 223 = 0
    16'b10011101_11100000 : OUT <= 0;  //157 / 224 = 0
    16'b10011101_11100001 : OUT <= 0;  //157 / 225 = 0
    16'b10011101_11100010 : OUT <= 0;  //157 / 226 = 0
    16'b10011101_11100011 : OUT <= 0;  //157 / 227 = 0
    16'b10011101_11100100 : OUT <= 0;  //157 / 228 = 0
    16'b10011101_11100101 : OUT <= 0;  //157 / 229 = 0
    16'b10011101_11100110 : OUT <= 0;  //157 / 230 = 0
    16'b10011101_11100111 : OUT <= 0;  //157 / 231 = 0
    16'b10011101_11101000 : OUT <= 0;  //157 / 232 = 0
    16'b10011101_11101001 : OUT <= 0;  //157 / 233 = 0
    16'b10011101_11101010 : OUT <= 0;  //157 / 234 = 0
    16'b10011101_11101011 : OUT <= 0;  //157 / 235 = 0
    16'b10011101_11101100 : OUT <= 0;  //157 / 236 = 0
    16'b10011101_11101101 : OUT <= 0;  //157 / 237 = 0
    16'b10011101_11101110 : OUT <= 0;  //157 / 238 = 0
    16'b10011101_11101111 : OUT <= 0;  //157 / 239 = 0
    16'b10011101_11110000 : OUT <= 0;  //157 / 240 = 0
    16'b10011101_11110001 : OUT <= 0;  //157 / 241 = 0
    16'b10011101_11110010 : OUT <= 0;  //157 / 242 = 0
    16'b10011101_11110011 : OUT <= 0;  //157 / 243 = 0
    16'b10011101_11110100 : OUT <= 0;  //157 / 244 = 0
    16'b10011101_11110101 : OUT <= 0;  //157 / 245 = 0
    16'b10011101_11110110 : OUT <= 0;  //157 / 246 = 0
    16'b10011101_11110111 : OUT <= 0;  //157 / 247 = 0
    16'b10011101_11111000 : OUT <= 0;  //157 / 248 = 0
    16'b10011101_11111001 : OUT <= 0;  //157 / 249 = 0
    16'b10011101_11111010 : OUT <= 0;  //157 / 250 = 0
    16'b10011101_11111011 : OUT <= 0;  //157 / 251 = 0
    16'b10011101_11111100 : OUT <= 0;  //157 / 252 = 0
    16'b10011101_11111101 : OUT <= 0;  //157 / 253 = 0
    16'b10011101_11111110 : OUT <= 0;  //157 / 254 = 0
    16'b10011101_11111111 : OUT <= 0;  //157 / 255 = 0
    16'b10011110_00000000 : OUT <= 0;  //158 / 0 = 0
    16'b10011110_00000001 : OUT <= 158;  //158 / 1 = 158
    16'b10011110_00000010 : OUT <= 79;  //158 / 2 = 79
    16'b10011110_00000011 : OUT <= 52;  //158 / 3 = 52
    16'b10011110_00000100 : OUT <= 39;  //158 / 4 = 39
    16'b10011110_00000101 : OUT <= 31;  //158 / 5 = 31
    16'b10011110_00000110 : OUT <= 26;  //158 / 6 = 26
    16'b10011110_00000111 : OUT <= 22;  //158 / 7 = 22
    16'b10011110_00001000 : OUT <= 19;  //158 / 8 = 19
    16'b10011110_00001001 : OUT <= 17;  //158 / 9 = 17
    16'b10011110_00001010 : OUT <= 15;  //158 / 10 = 15
    16'b10011110_00001011 : OUT <= 14;  //158 / 11 = 14
    16'b10011110_00001100 : OUT <= 13;  //158 / 12 = 13
    16'b10011110_00001101 : OUT <= 12;  //158 / 13 = 12
    16'b10011110_00001110 : OUT <= 11;  //158 / 14 = 11
    16'b10011110_00001111 : OUT <= 10;  //158 / 15 = 10
    16'b10011110_00010000 : OUT <= 9;  //158 / 16 = 9
    16'b10011110_00010001 : OUT <= 9;  //158 / 17 = 9
    16'b10011110_00010010 : OUT <= 8;  //158 / 18 = 8
    16'b10011110_00010011 : OUT <= 8;  //158 / 19 = 8
    16'b10011110_00010100 : OUT <= 7;  //158 / 20 = 7
    16'b10011110_00010101 : OUT <= 7;  //158 / 21 = 7
    16'b10011110_00010110 : OUT <= 7;  //158 / 22 = 7
    16'b10011110_00010111 : OUT <= 6;  //158 / 23 = 6
    16'b10011110_00011000 : OUT <= 6;  //158 / 24 = 6
    16'b10011110_00011001 : OUT <= 6;  //158 / 25 = 6
    16'b10011110_00011010 : OUT <= 6;  //158 / 26 = 6
    16'b10011110_00011011 : OUT <= 5;  //158 / 27 = 5
    16'b10011110_00011100 : OUT <= 5;  //158 / 28 = 5
    16'b10011110_00011101 : OUT <= 5;  //158 / 29 = 5
    16'b10011110_00011110 : OUT <= 5;  //158 / 30 = 5
    16'b10011110_00011111 : OUT <= 5;  //158 / 31 = 5
    16'b10011110_00100000 : OUT <= 4;  //158 / 32 = 4
    16'b10011110_00100001 : OUT <= 4;  //158 / 33 = 4
    16'b10011110_00100010 : OUT <= 4;  //158 / 34 = 4
    16'b10011110_00100011 : OUT <= 4;  //158 / 35 = 4
    16'b10011110_00100100 : OUT <= 4;  //158 / 36 = 4
    16'b10011110_00100101 : OUT <= 4;  //158 / 37 = 4
    16'b10011110_00100110 : OUT <= 4;  //158 / 38 = 4
    16'b10011110_00100111 : OUT <= 4;  //158 / 39 = 4
    16'b10011110_00101000 : OUT <= 3;  //158 / 40 = 3
    16'b10011110_00101001 : OUT <= 3;  //158 / 41 = 3
    16'b10011110_00101010 : OUT <= 3;  //158 / 42 = 3
    16'b10011110_00101011 : OUT <= 3;  //158 / 43 = 3
    16'b10011110_00101100 : OUT <= 3;  //158 / 44 = 3
    16'b10011110_00101101 : OUT <= 3;  //158 / 45 = 3
    16'b10011110_00101110 : OUT <= 3;  //158 / 46 = 3
    16'b10011110_00101111 : OUT <= 3;  //158 / 47 = 3
    16'b10011110_00110000 : OUT <= 3;  //158 / 48 = 3
    16'b10011110_00110001 : OUT <= 3;  //158 / 49 = 3
    16'b10011110_00110010 : OUT <= 3;  //158 / 50 = 3
    16'b10011110_00110011 : OUT <= 3;  //158 / 51 = 3
    16'b10011110_00110100 : OUT <= 3;  //158 / 52 = 3
    16'b10011110_00110101 : OUT <= 2;  //158 / 53 = 2
    16'b10011110_00110110 : OUT <= 2;  //158 / 54 = 2
    16'b10011110_00110111 : OUT <= 2;  //158 / 55 = 2
    16'b10011110_00111000 : OUT <= 2;  //158 / 56 = 2
    16'b10011110_00111001 : OUT <= 2;  //158 / 57 = 2
    16'b10011110_00111010 : OUT <= 2;  //158 / 58 = 2
    16'b10011110_00111011 : OUT <= 2;  //158 / 59 = 2
    16'b10011110_00111100 : OUT <= 2;  //158 / 60 = 2
    16'b10011110_00111101 : OUT <= 2;  //158 / 61 = 2
    16'b10011110_00111110 : OUT <= 2;  //158 / 62 = 2
    16'b10011110_00111111 : OUT <= 2;  //158 / 63 = 2
    16'b10011110_01000000 : OUT <= 2;  //158 / 64 = 2
    16'b10011110_01000001 : OUT <= 2;  //158 / 65 = 2
    16'b10011110_01000010 : OUT <= 2;  //158 / 66 = 2
    16'b10011110_01000011 : OUT <= 2;  //158 / 67 = 2
    16'b10011110_01000100 : OUT <= 2;  //158 / 68 = 2
    16'b10011110_01000101 : OUT <= 2;  //158 / 69 = 2
    16'b10011110_01000110 : OUT <= 2;  //158 / 70 = 2
    16'b10011110_01000111 : OUT <= 2;  //158 / 71 = 2
    16'b10011110_01001000 : OUT <= 2;  //158 / 72 = 2
    16'b10011110_01001001 : OUT <= 2;  //158 / 73 = 2
    16'b10011110_01001010 : OUT <= 2;  //158 / 74 = 2
    16'b10011110_01001011 : OUT <= 2;  //158 / 75 = 2
    16'b10011110_01001100 : OUT <= 2;  //158 / 76 = 2
    16'b10011110_01001101 : OUT <= 2;  //158 / 77 = 2
    16'b10011110_01001110 : OUT <= 2;  //158 / 78 = 2
    16'b10011110_01001111 : OUT <= 2;  //158 / 79 = 2
    16'b10011110_01010000 : OUT <= 1;  //158 / 80 = 1
    16'b10011110_01010001 : OUT <= 1;  //158 / 81 = 1
    16'b10011110_01010010 : OUT <= 1;  //158 / 82 = 1
    16'b10011110_01010011 : OUT <= 1;  //158 / 83 = 1
    16'b10011110_01010100 : OUT <= 1;  //158 / 84 = 1
    16'b10011110_01010101 : OUT <= 1;  //158 / 85 = 1
    16'b10011110_01010110 : OUT <= 1;  //158 / 86 = 1
    16'b10011110_01010111 : OUT <= 1;  //158 / 87 = 1
    16'b10011110_01011000 : OUT <= 1;  //158 / 88 = 1
    16'b10011110_01011001 : OUT <= 1;  //158 / 89 = 1
    16'b10011110_01011010 : OUT <= 1;  //158 / 90 = 1
    16'b10011110_01011011 : OUT <= 1;  //158 / 91 = 1
    16'b10011110_01011100 : OUT <= 1;  //158 / 92 = 1
    16'b10011110_01011101 : OUT <= 1;  //158 / 93 = 1
    16'b10011110_01011110 : OUT <= 1;  //158 / 94 = 1
    16'b10011110_01011111 : OUT <= 1;  //158 / 95 = 1
    16'b10011110_01100000 : OUT <= 1;  //158 / 96 = 1
    16'b10011110_01100001 : OUT <= 1;  //158 / 97 = 1
    16'b10011110_01100010 : OUT <= 1;  //158 / 98 = 1
    16'b10011110_01100011 : OUT <= 1;  //158 / 99 = 1
    16'b10011110_01100100 : OUT <= 1;  //158 / 100 = 1
    16'b10011110_01100101 : OUT <= 1;  //158 / 101 = 1
    16'b10011110_01100110 : OUT <= 1;  //158 / 102 = 1
    16'b10011110_01100111 : OUT <= 1;  //158 / 103 = 1
    16'b10011110_01101000 : OUT <= 1;  //158 / 104 = 1
    16'b10011110_01101001 : OUT <= 1;  //158 / 105 = 1
    16'b10011110_01101010 : OUT <= 1;  //158 / 106 = 1
    16'b10011110_01101011 : OUT <= 1;  //158 / 107 = 1
    16'b10011110_01101100 : OUT <= 1;  //158 / 108 = 1
    16'b10011110_01101101 : OUT <= 1;  //158 / 109 = 1
    16'b10011110_01101110 : OUT <= 1;  //158 / 110 = 1
    16'b10011110_01101111 : OUT <= 1;  //158 / 111 = 1
    16'b10011110_01110000 : OUT <= 1;  //158 / 112 = 1
    16'b10011110_01110001 : OUT <= 1;  //158 / 113 = 1
    16'b10011110_01110010 : OUT <= 1;  //158 / 114 = 1
    16'b10011110_01110011 : OUT <= 1;  //158 / 115 = 1
    16'b10011110_01110100 : OUT <= 1;  //158 / 116 = 1
    16'b10011110_01110101 : OUT <= 1;  //158 / 117 = 1
    16'b10011110_01110110 : OUT <= 1;  //158 / 118 = 1
    16'b10011110_01110111 : OUT <= 1;  //158 / 119 = 1
    16'b10011110_01111000 : OUT <= 1;  //158 / 120 = 1
    16'b10011110_01111001 : OUT <= 1;  //158 / 121 = 1
    16'b10011110_01111010 : OUT <= 1;  //158 / 122 = 1
    16'b10011110_01111011 : OUT <= 1;  //158 / 123 = 1
    16'b10011110_01111100 : OUT <= 1;  //158 / 124 = 1
    16'b10011110_01111101 : OUT <= 1;  //158 / 125 = 1
    16'b10011110_01111110 : OUT <= 1;  //158 / 126 = 1
    16'b10011110_01111111 : OUT <= 1;  //158 / 127 = 1
    16'b10011110_10000000 : OUT <= 1;  //158 / 128 = 1
    16'b10011110_10000001 : OUT <= 1;  //158 / 129 = 1
    16'b10011110_10000010 : OUT <= 1;  //158 / 130 = 1
    16'b10011110_10000011 : OUT <= 1;  //158 / 131 = 1
    16'b10011110_10000100 : OUT <= 1;  //158 / 132 = 1
    16'b10011110_10000101 : OUT <= 1;  //158 / 133 = 1
    16'b10011110_10000110 : OUT <= 1;  //158 / 134 = 1
    16'b10011110_10000111 : OUT <= 1;  //158 / 135 = 1
    16'b10011110_10001000 : OUT <= 1;  //158 / 136 = 1
    16'b10011110_10001001 : OUT <= 1;  //158 / 137 = 1
    16'b10011110_10001010 : OUT <= 1;  //158 / 138 = 1
    16'b10011110_10001011 : OUT <= 1;  //158 / 139 = 1
    16'b10011110_10001100 : OUT <= 1;  //158 / 140 = 1
    16'b10011110_10001101 : OUT <= 1;  //158 / 141 = 1
    16'b10011110_10001110 : OUT <= 1;  //158 / 142 = 1
    16'b10011110_10001111 : OUT <= 1;  //158 / 143 = 1
    16'b10011110_10010000 : OUT <= 1;  //158 / 144 = 1
    16'b10011110_10010001 : OUT <= 1;  //158 / 145 = 1
    16'b10011110_10010010 : OUT <= 1;  //158 / 146 = 1
    16'b10011110_10010011 : OUT <= 1;  //158 / 147 = 1
    16'b10011110_10010100 : OUT <= 1;  //158 / 148 = 1
    16'b10011110_10010101 : OUT <= 1;  //158 / 149 = 1
    16'b10011110_10010110 : OUT <= 1;  //158 / 150 = 1
    16'b10011110_10010111 : OUT <= 1;  //158 / 151 = 1
    16'b10011110_10011000 : OUT <= 1;  //158 / 152 = 1
    16'b10011110_10011001 : OUT <= 1;  //158 / 153 = 1
    16'b10011110_10011010 : OUT <= 1;  //158 / 154 = 1
    16'b10011110_10011011 : OUT <= 1;  //158 / 155 = 1
    16'b10011110_10011100 : OUT <= 1;  //158 / 156 = 1
    16'b10011110_10011101 : OUT <= 1;  //158 / 157 = 1
    16'b10011110_10011110 : OUT <= 1;  //158 / 158 = 1
    16'b10011110_10011111 : OUT <= 0;  //158 / 159 = 0
    16'b10011110_10100000 : OUT <= 0;  //158 / 160 = 0
    16'b10011110_10100001 : OUT <= 0;  //158 / 161 = 0
    16'b10011110_10100010 : OUT <= 0;  //158 / 162 = 0
    16'b10011110_10100011 : OUT <= 0;  //158 / 163 = 0
    16'b10011110_10100100 : OUT <= 0;  //158 / 164 = 0
    16'b10011110_10100101 : OUT <= 0;  //158 / 165 = 0
    16'b10011110_10100110 : OUT <= 0;  //158 / 166 = 0
    16'b10011110_10100111 : OUT <= 0;  //158 / 167 = 0
    16'b10011110_10101000 : OUT <= 0;  //158 / 168 = 0
    16'b10011110_10101001 : OUT <= 0;  //158 / 169 = 0
    16'b10011110_10101010 : OUT <= 0;  //158 / 170 = 0
    16'b10011110_10101011 : OUT <= 0;  //158 / 171 = 0
    16'b10011110_10101100 : OUT <= 0;  //158 / 172 = 0
    16'b10011110_10101101 : OUT <= 0;  //158 / 173 = 0
    16'b10011110_10101110 : OUT <= 0;  //158 / 174 = 0
    16'b10011110_10101111 : OUT <= 0;  //158 / 175 = 0
    16'b10011110_10110000 : OUT <= 0;  //158 / 176 = 0
    16'b10011110_10110001 : OUT <= 0;  //158 / 177 = 0
    16'b10011110_10110010 : OUT <= 0;  //158 / 178 = 0
    16'b10011110_10110011 : OUT <= 0;  //158 / 179 = 0
    16'b10011110_10110100 : OUT <= 0;  //158 / 180 = 0
    16'b10011110_10110101 : OUT <= 0;  //158 / 181 = 0
    16'b10011110_10110110 : OUT <= 0;  //158 / 182 = 0
    16'b10011110_10110111 : OUT <= 0;  //158 / 183 = 0
    16'b10011110_10111000 : OUT <= 0;  //158 / 184 = 0
    16'b10011110_10111001 : OUT <= 0;  //158 / 185 = 0
    16'b10011110_10111010 : OUT <= 0;  //158 / 186 = 0
    16'b10011110_10111011 : OUT <= 0;  //158 / 187 = 0
    16'b10011110_10111100 : OUT <= 0;  //158 / 188 = 0
    16'b10011110_10111101 : OUT <= 0;  //158 / 189 = 0
    16'b10011110_10111110 : OUT <= 0;  //158 / 190 = 0
    16'b10011110_10111111 : OUT <= 0;  //158 / 191 = 0
    16'b10011110_11000000 : OUT <= 0;  //158 / 192 = 0
    16'b10011110_11000001 : OUT <= 0;  //158 / 193 = 0
    16'b10011110_11000010 : OUT <= 0;  //158 / 194 = 0
    16'b10011110_11000011 : OUT <= 0;  //158 / 195 = 0
    16'b10011110_11000100 : OUT <= 0;  //158 / 196 = 0
    16'b10011110_11000101 : OUT <= 0;  //158 / 197 = 0
    16'b10011110_11000110 : OUT <= 0;  //158 / 198 = 0
    16'b10011110_11000111 : OUT <= 0;  //158 / 199 = 0
    16'b10011110_11001000 : OUT <= 0;  //158 / 200 = 0
    16'b10011110_11001001 : OUT <= 0;  //158 / 201 = 0
    16'b10011110_11001010 : OUT <= 0;  //158 / 202 = 0
    16'b10011110_11001011 : OUT <= 0;  //158 / 203 = 0
    16'b10011110_11001100 : OUT <= 0;  //158 / 204 = 0
    16'b10011110_11001101 : OUT <= 0;  //158 / 205 = 0
    16'b10011110_11001110 : OUT <= 0;  //158 / 206 = 0
    16'b10011110_11001111 : OUT <= 0;  //158 / 207 = 0
    16'b10011110_11010000 : OUT <= 0;  //158 / 208 = 0
    16'b10011110_11010001 : OUT <= 0;  //158 / 209 = 0
    16'b10011110_11010010 : OUT <= 0;  //158 / 210 = 0
    16'b10011110_11010011 : OUT <= 0;  //158 / 211 = 0
    16'b10011110_11010100 : OUT <= 0;  //158 / 212 = 0
    16'b10011110_11010101 : OUT <= 0;  //158 / 213 = 0
    16'b10011110_11010110 : OUT <= 0;  //158 / 214 = 0
    16'b10011110_11010111 : OUT <= 0;  //158 / 215 = 0
    16'b10011110_11011000 : OUT <= 0;  //158 / 216 = 0
    16'b10011110_11011001 : OUT <= 0;  //158 / 217 = 0
    16'b10011110_11011010 : OUT <= 0;  //158 / 218 = 0
    16'b10011110_11011011 : OUT <= 0;  //158 / 219 = 0
    16'b10011110_11011100 : OUT <= 0;  //158 / 220 = 0
    16'b10011110_11011101 : OUT <= 0;  //158 / 221 = 0
    16'b10011110_11011110 : OUT <= 0;  //158 / 222 = 0
    16'b10011110_11011111 : OUT <= 0;  //158 / 223 = 0
    16'b10011110_11100000 : OUT <= 0;  //158 / 224 = 0
    16'b10011110_11100001 : OUT <= 0;  //158 / 225 = 0
    16'b10011110_11100010 : OUT <= 0;  //158 / 226 = 0
    16'b10011110_11100011 : OUT <= 0;  //158 / 227 = 0
    16'b10011110_11100100 : OUT <= 0;  //158 / 228 = 0
    16'b10011110_11100101 : OUT <= 0;  //158 / 229 = 0
    16'b10011110_11100110 : OUT <= 0;  //158 / 230 = 0
    16'b10011110_11100111 : OUT <= 0;  //158 / 231 = 0
    16'b10011110_11101000 : OUT <= 0;  //158 / 232 = 0
    16'b10011110_11101001 : OUT <= 0;  //158 / 233 = 0
    16'b10011110_11101010 : OUT <= 0;  //158 / 234 = 0
    16'b10011110_11101011 : OUT <= 0;  //158 / 235 = 0
    16'b10011110_11101100 : OUT <= 0;  //158 / 236 = 0
    16'b10011110_11101101 : OUT <= 0;  //158 / 237 = 0
    16'b10011110_11101110 : OUT <= 0;  //158 / 238 = 0
    16'b10011110_11101111 : OUT <= 0;  //158 / 239 = 0
    16'b10011110_11110000 : OUT <= 0;  //158 / 240 = 0
    16'b10011110_11110001 : OUT <= 0;  //158 / 241 = 0
    16'b10011110_11110010 : OUT <= 0;  //158 / 242 = 0
    16'b10011110_11110011 : OUT <= 0;  //158 / 243 = 0
    16'b10011110_11110100 : OUT <= 0;  //158 / 244 = 0
    16'b10011110_11110101 : OUT <= 0;  //158 / 245 = 0
    16'b10011110_11110110 : OUT <= 0;  //158 / 246 = 0
    16'b10011110_11110111 : OUT <= 0;  //158 / 247 = 0
    16'b10011110_11111000 : OUT <= 0;  //158 / 248 = 0
    16'b10011110_11111001 : OUT <= 0;  //158 / 249 = 0
    16'b10011110_11111010 : OUT <= 0;  //158 / 250 = 0
    16'b10011110_11111011 : OUT <= 0;  //158 / 251 = 0
    16'b10011110_11111100 : OUT <= 0;  //158 / 252 = 0
    16'b10011110_11111101 : OUT <= 0;  //158 / 253 = 0
    16'b10011110_11111110 : OUT <= 0;  //158 / 254 = 0
    16'b10011110_11111111 : OUT <= 0;  //158 / 255 = 0
    16'b10011111_00000000 : OUT <= 0;  //159 / 0 = 0
    16'b10011111_00000001 : OUT <= 159;  //159 / 1 = 159
    16'b10011111_00000010 : OUT <= 79;  //159 / 2 = 79
    16'b10011111_00000011 : OUT <= 53;  //159 / 3 = 53
    16'b10011111_00000100 : OUT <= 39;  //159 / 4 = 39
    16'b10011111_00000101 : OUT <= 31;  //159 / 5 = 31
    16'b10011111_00000110 : OUT <= 26;  //159 / 6 = 26
    16'b10011111_00000111 : OUT <= 22;  //159 / 7 = 22
    16'b10011111_00001000 : OUT <= 19;  //159 / 8 = 19
    16'b10011111_00001001 : OUT <= 17;  //159 / 9 = 17
    16'b10011111_00001010 : OUT <= 15;  //159 / 10 = 15
    16'b10011111_00001011 : OUT <= 14;  //159 / 11 = 14
    16'b10011111_00001100 : OUT <= 13;  //159 / 12 = 13
    16'b10011111_00001101 : OUT <= 12;  //159 / 13 = 12
    16'b10011111_00001110 : OUT <= 11;  //159 / 14 = 11
    16'b10011111_00001111 : OUT <= 10;  //159 / 15 = 10
    16'b10011111_00010000 : OUT <= 9;  //159 / 16 = 9
    16'b10011111_00010001 : OUT <= 9;  //159 / 17 = 9
    16'b10011111_00010010 : OUT <= 8;  //159 / 18 = 8
    16'b10011111_00010011 : OUT <= 8;  //159 / 19 = 8
    16'b10011111_00010100 : OUT <= 7;  //159 / 20 = 7
    16'b10011111_00010101 : OUT <= 7;  //159 / 21 = 7
    16'b10011111_00010110 : OUT <= 7;  //159 / 22 = 7
    16'b10011111_00010111 : OUT <= 6;  //159 / 23 = 6
    16'b10011111_00011000 : OUT <= 6;  //159 / 24 = 6
    16'b10011111_00011001 : OUT <= 6;  //159 / 25 = 6
    16'b10011111_00011010 : OUT <= 6;  //159 / 26 = 6
    16'b10011111_00011011 : OUT <= 5;  //159 / 27 = 5
    16'b10011111_00011100 : OUT <= 5;  //159 / 28 = 5
    16'b10011111_00011101 : OUT <= 5;  //159 / 29 = 5
    16'b10011111_00011110 : OUT <= 5;  //159 / 30 = 5
    16'b10011111_00011111 : OUT <= 5;  //159 / 31 = 5
    16'b10011111_00100000 : OUT <= 4;  //159 / 32 = 4
    16'b10011111_00100001 : OUT <= 4;  //159 / 33 = 4
    16'b10011111_00100010 : OUT <= 4;  //159 / 34 = 4
    16'b10011111_00100011 : OUT <= 4;  //159 / 35 = 4
    16'b10011111_00100100 : OUT <= 4;  //159 / 36 = 4
    16'b10011111_00100101 : OUT <= 4;  //159 / 37 = 4
    16'b10011111_00100110 : OUT <= 4;  //159 / 38 = 4
    16'b10011111_00100111 : OUT <= 4;  //159 / 39 = 4
    16'b10011111_00101000 : OUT <= 3;  //159 / 40 = 3
    16'b10011111_00101001 : OUT <= 3;  //159 / 41 = 3
    16'b10011111_00101010 : OUT <= 3;  //159 / 42 = 3
    16'b10011111_00101011 : OUT <= 3;  //159 / 43 = 3
    16'b10011111_00101100 : OUT <= 3;  //159 / 44 = 3
    16'b10011111_00101101 : OUT <= 3;  //159 / 45 = 3
    16'b10011111_00101110 : OUT <= 3;  //159 / 46 = 3
    16'b10011111_00101111 : OUT <= 3;  //159 / 47 = 3
    16'b10011111_00110000 : OUT <= 3;  //159 / 48 = 3
    16'b10011111_00110001 : OUT <= 3;  //159 / 49 = 3
    16'b10011111_00110010 : OUT <= 3;  //159 / 50 = 3
    16'b10011111_00110011 : OUT <= 3;  //159 / 51 = 3
    16'b10011111_00110100 : OUT <= 3;  //159 / 52 = 3
    16'b10011111_00110101 : OUT <= 3;  //159 / 53 = 3
    16'b10011111_00110110 : OUT <= 2;  //159 / 54 = 2
    16'b10011111_00110111 : OUT <= 2;  //159 / 55 = 2
    16'b10011111_00111000 : OUT <= 2;  //159 / 56 = 2
    16'b10011111_00111001 : OUT <= 2;  //159 / 57 = 2
    16'b10011111_00111010 : OUT <= 2;  //159 / 58 = 2
    16'b10011111_00111011 : OUT <= 2;  //159 / 59 = 2
    16'b10011111_00111100 : OUT <= 2;  //159 / 60 = 2
    16'b10011111_00111101 : OUT <= 2;  //159 / 61 = 2
    16'b10011111_00111110 : OUT <= 2;  //159 / 62 = 2
    16'b10011111_00111111 : OUT <= 2;  //159 / 63 = 2
    16'b10011111_01000000 : OUT <= 2;  //159 / 64 = 2
    16'b10011111_01000001 : OUT <= 2;  //159 / 65 = 2
    16'b10011111_01000010 : OUT <= 2;  //159 / 66 = 2
    16'b10011111_01000011 : OUT <= 2;  //159 / 67 = 2
    16'b10011111_01000100 : OUT <= 2;  //159 / 68 = 2
    16'b10011111_01000101 : OUT <= 2;  //159 / 69 = 2
    16'b10011111_01000110 : OUT <= 2;  //159 / 70 = 2
    16'b10011111_01000111 : OUT <= 2;  //159 / 71 = 2
    16'b10011111_01001000 : OUT <= 2;  //159 / 72 = 2
    16'b10011111_01001001 : OUT <= 2;  //159 / 73 = 2
    16'b10011111_01001010 : OUT <= 2;  //159 / 74 = 2
    16'b10011111_01001011 : OUT <= 2;  //159 / 75 = 2
    16'b10011111_01001100 : OUT <= 2;  //159 / 76 = 2
    16'b10011111_01001101 : OUT <= 2;  //159 / 77 = 2
    16'b10011111_01001110 : OUT <= 2;  //159 / 78 = 2
    16'b10011111_01001111 : OUT <= 2;  //159 / 79 = 2
    16'b10011111_01010000 : OUT <= 1;  //159 / 80 = 1
    16'b10011111_01010001 : OUT <= 1;  //159 / 81 = 1
    16'b10011111_01010010 : OUT <= 1;  //159 / 82 = 1
    16'b10011111_01010011 : OUT <= 1;  //159 / 83 = 1
    16'b10011111_01010100 : OUT <= 1;  //159 / 84 = 1
    16'b10011111_01010101 : OUT <= 1;  //159 / 85 = 1
    16'b10011111_01010110 : OUT <= 1;  //159 / 86 = 1
    16'b10011111_01010111 : OUT <= 1;  //159 / 87 = 1
    16'b10011111_01011000 : OUT <= 1;  //159 / 88 = 1
    16'b10011111_01011001 : OUT <= 1;  //159 / 89 = 1
    16'b10011111_01011010 : OUT <= 1;  //159 / 90 = 1
    16'b10011111_01011011 : OUT <= 1;  //159 / 91 = 1
    16'b10011111_01011100 : OUT <= 1;  //159 / 92 = 1
    16'b10011111_01011101 : OUT <= 1;  //159 / 93 = 1
    16'b10011111_01011110 : OUT <= 1;  //159 / 94 = 1
    16'b10011111_01011111 : OUT <= 1;  //159 / 95 = 1
    16'b10011111_01100000 : OUT <= 1;  //159 / 96 = 1
    16'b10011111_01100001 : OUT <= 1;  //159 / 97 = 1
    16'b10011111_01100010 : OUT <= 1;  //159 / 98 = 1
    16'b10011111_01100011 : OUT <= 1;  //159 / 99 = 1
    16'b10011111_01100100 : OUT <= 1;  //159 / 100 = 1
    16'b10011111_01100101 : OUT <= 1;  //159 / 101 = 1
    16'b10011111_01100110 : OUT <= 1;  //159 / 102 = 1
    16'b10011111_01100111 : OUT <= 1;  //159 / 103 = 1
    16'b10011111_01101000 : OUT <= 1;  //159 / 104 = 1
    16'b10011111_01101001 : OUT <= 1;  //159 / 105 = 1
    16'b10011111_01101010 : OUT <= 1;  //159 / 106 = 1
    16'b10011111_01101011 : OUT <= 1;  //159 / 107 = 1
    16'b10011111_01101100 : OUT <= 1;  //159 / 108 = 1
    16'b10011111_01101101 : OUT <= 1;  //159 / 109 = 1
    16'b10011111_01101110 : OUT <= 1;  //159 / 110 = 1
    16'b10011111_01101111 : OUT <= 1;  //159 / 111 = 1
    16'b10011111_01110000 : OUT <= 1;  //159 / 112 = 1
    16'b10011111_01110001 : OUT <= 1;  //159 / 113 = 1
    16'b10011111_01110010 : OUT <= 1;  //159 / 114 = 1
    16'b10011111_01110011 : OUT <= 1;  //159 / 115 = 1
    16'b10011111_01110100 : OUT <= 1;  //159 / 116 = 1
    16'b10011111_01110101 : OUT <= 1;  //159 / 117 = 1
    16'b10011111_01110110 : OUT <= 1;  //159 / 118 = 1
    16'b10011111_01110111 : OUT <= 1;  //159 / 119 = 1
    16'b10011111_01111000 : OUT <= 1;  //159 / 120 = 1
    16'b10011111_01111001 : OUT <= 1;  //159 / 121 = 1
    16'b10011111_01111010 : OUT <= 1;  //159 / 122 = 1
    16'b10011111_01111011 : OUT <= 1;  //159 / 123 = 1
    16'b10011111_01111100 : OUT <= 1;  //159 / 124 = 1
    16'b10011111_01111101 : OUT <= 1;  //159 / 125 = 1
    16'b10011111_01111110 : OUT <= 1;  //159 / 126 = 1
    16'b10011111_01111111 : OUT <= 1;  //159 / 127 = 1
    16'b10011111_10000000 : OUT <= 1;  //159 / 128 = 1
    16'b10011111_10000001 : OUT <= 1;  //159 / 129 = 1
    16'b10011111_10000010 : OUT <= 1;  //159 / 130 = 1
    16'b10011111_10000011 : OUT <= 1;  //159 / 131 = 1
    16'b10011111_10000100 : OUT <= 1;  //159 / 132 = 1
    16'b10011111_10000101 : OUT <= 1;  //159 / 133 = 1
    16'b10011111_10000110 : OUT <= 1;  //159 / 134 = 1
    16'b10011111_10000111 : OUT <= 1;  //159 / 135 = 1
    16'b10011111_10001000 : OUT <= 1;  //159 / 136 = 1
    16'b10011111_10001001 : OUT <= 1;  //159 / 137 = 1
    16'b10011111_10001010 : OUT <= 1;  //159 / 138 = 1
    16'b10011111_10001011 : OUT <= 1;  //159 / 139 = 1
    16'b10011111_10001100 : OUT <= 1;  //159 / 140 = 1
    16'b10011111_10001101 : OUT <= 1;  //159 / 141 = 1
    16'b10011111_10001110 : OUT <= 1;  //159 / 142 = 1
    16'b10011111_10001111 : OUT <= 1;  //159 / 143 = 1
    16'b10011111_10010000 : OUT <= 1;  //159 / 144 = 1
    16'b10011111_10010001 : OUT <= 1;  //159 / 145 = 1
    16'b10011111_10010010 : OUT <= 1;  //159 / 146 = 1
    16'b10011111_10010011 : OUT <= 1;  //159 / 147 = 1
    16'b10011111_10010100 : OUT <= 1;  //159 / 148 = 1
    16'b10011111_10010101 : OUT <= 1;  //159 / 149 = 1
    16'b10011111_10010110 : OUT <= 1;  //159 / 150 = 1
    16'b10011111_10010111 : OUT <= 1;  //159 / 151 = 1
    16'b10011111_10011000 : OUT <= 1;  //159 / 152 = 1
    16'b10011111_10011001 : OUT <= 1;  //159 / 153 = 1
    16'b10011111_10011010 : OUT <= 1;  //159 / 154 = 1
    16'b10011111_10011011 : OUT <= 1;  //159 / 155 = 1
    16'b10011111_10011100 : OUT <= 1;  //159 / 156 = 1
    16'b10011111_10011101 : OUT <= 1;  //159 / 157 = 1
    16'b10011111_10011110 : OUT <= 1;  //159 / 158 = 1
    16'b10011111_10011111 : OUT <= 1;  //159 / 159 = 1
    16'b10011111_10100000 : OUT <= 0;  //159 / 160 = 0
    16'b10011111_10100001 : OUT <= 0;  //159 / 161 = 0
    16'b10011111_10100010 : OUT <= 0;  //159 / 162 = 0
    16'b10011111_10100011 : OUT <= 0;  //159 / 163 = 0
    16'b10011111_10100100 : OUT <= 0;  //159 / 164 = 0
    16'b10011111_10100101 : OUT <= 0;  //159 / 165 = 0
    16'b10011111_10100110 : OUT <= 0;  //159 / 166 = 0
    16'b10011111_10100111 : OUT <= 0;  //159 / 167 = 0
    16'b10011111_10101000 : OUT <= 0;  //159 / 168 = 0
    16'b10011111_10101001 : OUT <= 0;  //159 / 169 = 0
    16'b10011111_10101010 : OUT <= 0;  //159 / 170 = 0
    16'b10011111_10101011 : OUT <= 0;  //159 / 171 = 0
    16'b10011111_10101100 : OUT <= 0;  //159 / 172 = 0
    16'b10011111_10101101 : OUT <= 0;  //159 / 173 = 0
    16'b10011111_10101110 : OUT <= 0;  //159 / 174 = 0
    16'b10011111_10101111 : OUT <= 0;  //159 / 175 = 0
    16'b10011111_10110000 : OUT <= 0;  //159 / 176 = 0
    16'b10011111_10110001 : OUT <= 0;  //159 / 177 = 0
    16'b10011111_10110010 : OUT <= 0;  //159 / 178 = 0
    16'b10011111_10110011 : OUT <= 0;  //159 / 179 = 0
    16'b10011111_10110100 : OUT <= 0;  //159 / 180 = 0
    16'b10011111_10110101 : OUT <= 0;  //159 / 181 = 0
    16'b10011111_10110110 : OUT <= 0;  //159 / 182 = 0
    16'b10011111_10110111 : OUT <= 0;  //159 / 183 = 0
    16'b10011111_10111000 : OUT <= 0;  //159 / 184 = 0
    16'b10011111_10111001 : OUT <= 0;  //159 / 185 = 0
    16'b10011111_10111010 : OUT <= 0;  //159 / 186 = 0
    16'b10011111_10111011 : OUT <= 0;  //159 / 187 = 0
    16'b10011111_10111100 : OUT <= 0;  //159 / 188 = 0
    16'b10011111_10111101 : OUT <= 0;  //159 / 189 = 0
    16'b10011111_10111110 : OUT <= 0;  //159 / 190 = 0
    16'b10011111_10111111 : OUT <= 0;  //159 / 191 = 0
    16'b10011111_11000000 : OUT <= 0;  //159 / 192 = 0
    16'b10011111_11000001 : OUT <= 0;  //159 / 193 = 0
    16'b10011111_11000010 : OUT <= 0;  //159 / 194 = 0
    16'b10011111_11000011 : OUT <= 0;  //159 / 195 = 0
    16'b10011111_11000100 : OUT <= 0;  //159 / 196 = 0
    16'b10011111_11000101 : OUT <= 0;  //159 / 197 = 0
    16'b10011111_11000110 : OUT <= 0;  //159 / 198 = 0
    16'b10011111_11000111 : OUT <= 0;  //159 / 199 = 0
    16'b10011111_11001000 : OUT <= 0;  //159 / 200 = 0
    16'b10011111_11001001 : OUT <= 0;  //159 / 201 = 0
    16'b10011111_11001010 : OUT <= 0;  //159 / 202 = 0
    16'b10011111_11001011 : OUT <= 0;  //159 / 203 = 0
    16'b10011111_11001100 : OUT <= 0;  //159 / 204 = 0
    16'b10011111_11001101 : OUT <= 0;  //159 / 205 = 0
    16'b10011111_11001110 : OUT <= 0;  //159 / 206 = 0
    16'b10011111_11001111 : OUT <= 0;  //159 / 207 = 0
    16'b10011111_11010000 : OUT <= 0;  //159 / 208 = 0
    16'b10011111_11010001 : OUT <= 0;  //159 / 209 = 0
    16'b10011111_11010010 : OUT <= 0;  //159 / 210 = 0
    16'b10011111_11010011 : OUT <= 0;  //159 / 211 = 0
    16'b10011111_11010100 : OUT <= 0;  //159 / 212 = 0
    16'b10011111_11010101 : OUT <= 0;  //159 / 213 = 0
    16'b10011111_11010110 : OUT <= 0;  //159 / 214 = 0
    16'b10011111_11010111 : OUT <= 0;  //159 / 215 = 0
    16'b10011111_11011000 : OUT <= 0;  //159 / 216 = 0
    16'b10011111_11011001 : OUT <= 0;  //159 / 217 = 0
    16'b10011111_11011010 : OUT <= 0;  //159 / 218 = 0
    16'b10011111_11011011 : OUT <= 0;  //159 / 219 = 0
    16'b10011111_11011100 : OUT <= 0;  //159 / 220 = 0
    16'b10011111_11011101 : OUT <= 0;  //159 / 221 = 0
    16'b10011111_11011110 : OUT <= 0;  //159 / 222 = 0
    16'b10011111_11011111 : OUT <= 0;  //159 / 223 = 0
    16'b10011111_11100000 : OUT <= 0;  //159 / 224 = 0
    16'b10011111_11100001 : OUT <= 0;  //159 / 225 = 0
    16'b10011111_11100010 : OUT <= 0;  //159 / 226 = 0
    16'b10011111_11100011 : OUT <= 0;  //159 / 227 = 0
    16'b10011111_11100100 : OUT <= 0;  //159 / 228 = 0
    16'b10011111_11100101 : OUT <= 0;  //159 / 229 = 0
    16'b10011111_11100110 : OUT <= 0;  //159 / 230 = 0
    16'b10011111_11100111 : OUT <= 0;  //159 / 231 = 0
    16'b10011111_11101000 : OUT <= 0;  //159 / 232 = 0
    16'b10011111_11101001 : OUT <= 0;  //159 / 233 = 0
    16'b10011111_11101010 : OUT <= 0;  //159 / 234 = 0
    16'b10011111_11101011 : OUT <= 0;  //159 / 235 = 0
    16'b10011111_11101100 : OUT <= 0;  //159 / 236 = 0
    16'b10011111_11101101 : OUT <= 0;  //159 / 237 = 0
    16'b10011111_11101110 : OUT <= 0;  //159 / 238 = 0
    16'b10011111_11101111 : OUT <= 0;  //159 / 239 = 0
    16'b10011111_11110000 : OUT <= 0;  //159 / 240 = 0
    16'b10011111_11110001 : OUT <= 0;  //159 / 241 = 0
    16'b10011111_11110010 : OUT <= 0;  //159 / 242 = 0
    16'b10011111_11110011 : OUT <= 0;  //159 / 243 = 0
    16'b10011111_11110100 : OUT <= 0;  //159 / 244 = 0
    16'b10011111_11110101 : OUT <= 0;  //159 / 245 = 0
    16'b10011111_11110110 : OUT <= 0;  //159 / 246 = 0
    16'b10011111_11110111 : OUT <= 0;  //159 / 247 = 0
    16'b10011111_11111000 : OUT <= 0;  //159 / 248 = 0
    16'b10011111_11111001 : OUT <= 0;  //159 / 249 = 0
    16'b10011111_11111010 : OUT <= 0;  //159 / 250 = 0
    16'b10011111_11111011 : OUT <= 0;  //159 / 251 = 0
    16'b10011111_11111100 : OUT <= 0;  //159 / 252 = 0
    16'b10011111_11111101 : OUT <= 0;  //159 / 253 = 0
    16'b10011111_11111110 : OUT <= 0;  //159 / 254 = 0
    16'b10011111_11111111 : OUT <= 0;  //159 / 255 = 0
    16'b10100000_00000000 : OUT <= 0;  //160 / 0 = 0
    16'b10100000_00000001 : OUT <= 160;  //160 / 1 = 160
    16'b10100000_00000010 : OUT <= 80;  //160 / 2 = 80
    16'b10100000_00000011 : OUT <= 53;  //160 / 3 = 53
    16'b10100000_00000100 : OUT <= 40;  //160 / 4 = 40
    16'b10100000_00000101 : OUT <= 32;  //160 / 5 = 32
    16'b10100000_00000110 : OUT <= 26;  //160 / 6 = 26
    16'b10100000_00000111 : OUT <= 22;  //160 / 7 = 22
    16'b10100000_00001000 : OUT <= 20;  //160 / 8 = 20
    16'b10100000_00001001 : OUT <= 17;  //160 / 9 = 17
    16'b10100000_00001010 : OUT <= 16;  //160 / 10 = 16
    16'b10100000_00001011 : OUT <= 14;  //160 / 11 = 14
    16'b10100000_00001100 : OUT <= 13;  //160 / 12 = 13
    16'b10100000_00001101 : OUT <= 12;  //160 / 13 = 12
    16'b10100000_00001110 : OUT <= 11;  //160 / 14 = 11
    16'b10100000_00001111 : OUT <= 10;  //160 / 15 = 10
    16'b10100000_00010000 : OUT <= 10;  //160 / 16 = 10
    16'b10100000_00010001 : OUT <= 9;  //160 / 17 = 9
    16'b10100000_00010010 : OUT <= 8;  //160 / 18 = 8
    16'b10100000_00010011 : OUT <= 8;  //160 / 19 = 8
    16'b10100000_00010100 : OUT <= 8;  //160 / 20 = 8
    16'b10100000_00010101 : OUT <= 7;  //160 / 21 = 7
    16'b10100000_00010110 : OUT <= 7;  //160 / 22 = 7
    16'b10100000_00010111 : OUT <= 6;  //160 / 23 = 6
    16'b10100000_00011000 : OUT <= 6;  //160 / 24 = 6
    16'b10100000_00011001 : OUT <= 6;  //160 / 25 = 6
    16'b10100000_00011010 : OUT <= 6;  //160 / 26 = 6
    16'b10100000_00011011 : OUT <= 5;  //160 / 27 = 5
    16'b10100000_00011100 : OUT <= 5;  //160 / 28 = 5
    16'b10100000_00011101 : OUT <= 5;  //160 / 29 = 5
    16'b10100000_00011110 : OUT <= 5;  //160 / 30 = 5
    16'b10100000_00011111 : OUT <= 5;  //160 / 31 = 5
    16'b10100000_00100000 : OUT <= 5;  //160 / 32 = 5
    16'b10100000_00100001 : OUT <= 4;  //160 / 33 = 4
    16'b10100000_00100010 : OUT <= 4;  //160 / 34 = 4
    16'b10100000_00100011 : OUT <= 4;  //160 / 35 = 4
    16'b10100000_00100100 : OUT <= 4;  //160 / 36 = 4
    16'b10100000_00100101 : OUT <= 4;  //160 / 37 = 4
    16'b10100000_00100110 : OUT <= 4;  //160 / 38 = 4
    16'b10100000_00100111 : OUT <= 4;  //160 / 39 = 4
    16'b10100000_00101000 : OUT <= 4;  //160 / 40 = 4
    16'b10100000_00101001 : OUT <= 3;  //160 / 41 = 3
    16'b10100000_00101010 : OUT <= 3;  //160 / 42 = 3
    16'b10100000_00101011 : OUT <= 3;  //160 / 43 = 3
    16'b10100000_00101100 : OUT <= 3;  //160 / 44 = 3
    16'b10100000_00101101 : OUT <= 3;  //160 / 45 = 3
    16'b10100000_00101110 : OUT <= 3;  //160 / 46 = 3
    16'b10100000_00101111 : OUT <= 3;  //160 / 47 = 3
    16'b10100000_00110000 : OUT <= 3;  //160 / 48 = 3
    16'b10100000_00110001 : OUT <= 3;  //160 / 49 = 3
    16'b10100000_00110010 : OUT <= 3;  //160 / 50 = 3
    16'b10100000_00110011 : OUT <= 3;  //160 / 51 = 3
    16'b10100000_00110100 : OUT <= 3;  //160 / 52 = 3
    16'b10100000_00110101 : OUT <= 3;  //160 / 53 = 3
    16'b10100000_00110110 : OUT <= 2;  //160 / 54 = 2
    16'b10100000_00110111 : OUT <= 2;  //160 / 55 = 2
    16'b10100000_00111000 : OUT <= 2;  //160 / 56 = 2
    16'b10100000_00111001 : OUT <= 2;  //160 / 57 = 2
    16'b10100000_00111010 : OUT <= 2;  //160 / 58 = 2
    16'b10100000_00111011 : OUT <= 2;  //160 / 59 = 2
    16'b10100000_00111100 : OUT <= 2;  //160 / 60 = 2
    16'b10100000_00111101 : OUT <= 2;  //160 / 61 = 2
    16'b10100000_00111110 : OUT <= 2;  //160 / 62 = 2
    16'b10100000_00111111 : OUT <= 2;  //160 / 63 = 2
    16'b10100000_01000000 : OUT <= 2;  //160 / 64 = 2
    16'b10100000_01000001 : OUT <= 2;  //160 / 65 = 2
    16'b10100000_01000010 : OUT <= 2;  //160 / 66 = 2
    16'b10100000_01000011 : OUT <= 2;  //160 / 67 = 2
    16'b10100000_01000100 : OUT <= 2;  //160 / 68 = 2
    16'b10100000_01000101 : OUT <= 2;  //160 / 69 = 2
    16'b10100000_01000110 : OUT <= 2;  //160 / 70 = 2
    16'b10100000_01000111 : OUT <= 2;  //160 / 71 = 2
    16'b10100000_01001000 : OUT <= 2;  //160 / 72 = 2
    16'b10100000_01001001 : OUT <= 2;  //160 / 73 = 2
    16'b10100000_01001010 : OUT <= 2;  //160 / 74 = 2
    16'b10100000_01001011 : OUT <= 2;  //160 / 75 = 2
    16'b10100000_01001100 : OUT <= 2;  //160 / 76 = 2
    16'b10100000_01001101 : OUT <= 2;  //160 / 77 = 2
    16'b10100000_01001110 : OUT <= 2;  //160 / 78 = 2
    16'b10100000_01001111 : OUT <= 2;  //160 / 79 = 2
    16'b10100000_01010000 : OUT <= 2;  //160 / 80 = 2
    16'b10100000_01010001 : OUT <= 1;  //160 / 81 = 1
    16'b10100000_01010010 : OUT <= 1;  //160 / 82 = 1
    16'b10100000_01010011 : OUT <= 1;  //160 / 83 = 1
    16'b10100000_01010100 : OUT <= 1;  //160 / 84 = 1
    16'b10100000_01010101 : OUT <= 1;  //160 / 85 = 1
    16'b10100000_01010110 : OUT <= 1;  //160 / 86 = 1
    16'b10100000_01010111 : OUT <= 1;  //160 / 87 = 1
    16'b10100000_01011000 : OUT <= 1;  //160 / 88 = 1
    16'b10100000_01011001 : OUT <= 1;  //160 / 89 = 1
    16'b10100000_01011010 : OUT <= 1;  //160 / 90 = 1
    16'b10100000_01011011 : OUT <= 1;  //160 / 91 = 1
    16'b10100000_01011100 : OUT <= 1;  //160 / 92 = 1
    16'b10100000_01011101 : OUT <= 1;  //160 / 93 = 1
    16'b10100000_01011110 : OUT <= 1;  //160 / 94 = 1
    16'b10100000_01011111 : OUT <= 1;  //160 / 95 = 1
    16'b10100000_01100000 : OUT <= 1;  //160 / 96 = 1
    16'b10100000_01100001 : OUT <= 1;  //160 / 97 = 1
    16'b10100000_01100010 : OUT <= 1;  //160 / 98 = 1
    16'b10100000_01100011 : OUT <= 1;  //160 / 99 = 1
    16'b10100000_01100100 : OUT <= 1;  //160 / 100 = 1
    16'b10100000_01100101 : OUT <= 1;  //160 / 101 = 1
    16'b10100000_01100110 : OUT <= 1;  //160 / 102 = 1
    16'b10100000_01100111 : OUT <= 1;  //160 / 103 = 1
    16'b10100000_01101000 : OUT <= 1;  //160 / 104 = 1
    16'b10100000_01101001 : OUT <= 1;  //160 / 105 = 1
    16'b10100000_01101010 : OUT <= 1;  //160 / 106 = 1
    16'b10100000_01101011 : OUT <= 1;  //160 / 107 = 1
    16'b10100000_01101100 : OUT <= 1;  //160 / 108 = 1
    16'b10100000_01101101 : OUT <= 1;  //160 / 109 = 1
    16'b10100000_01101110 : OUT <= 1;  //160 / 110 = 1
    16'b10100000_01101111 : OUT <= 1;  //160 / 111 = 1
    16'b10100000_01110000 : OUT <= 1;  //160 / 112 = 1
    16'b10100000_01110001 : OUT <= 1;  //160 / 113 = 1
    16'b10100000_01110010 : OUT <= 1;  //160 / 114 = 1
    16'b10100000_01110011 : OUT <= 1;  //160 / 115 = 1
    16'b10100000_01110100 : OUT <= 1;  //160 / 116 = 1
    16'b10100000_01110101 : OUT <= 1;  //160 / 117 = 1
    16'b10100000_01110110 : OUT <= 1;  //160 / 118 = 1
    16'b10100000_01110111 : OUT <= 1;  //160 / 119 = 1
    16'b10100000_01111000 : OUT <= 1;  //160 / 120 = 1
    16'b10100000_01111001 : OUT <= 1;  //160 / 121 = 1
    16'b10100000_01111010 : OUT <= 1;  //160 / 122 = 1
    16'b10100000_01111011 : OUT <= 1;  //160 / 123 = 1
    16'b10100000_01111100 : OUT <= 1;  //160 / 124 = 1
    16'b10100000_01111101 : OUT <= 1;  //160 / 125 = 1
    16'b10100000_01111110 : OUT <= 1;  //160 / 126 = 1
    16'b10100000_01111111 : OUT <= 1;  //160 / 127 = 1
    16'b10100000_10000000 : OUT <= 1;  //160 / 128 = 1
    16'b10100000_10000001 : OUT <= 1;  //160 / 129 = 1
    16'b10100000_10000010 : OUT <= 1;  //160 / 130 = 1
    16'b10100000_10000011 : OUT <= 1;  //160 / 131 = 1
    16'b10100000_10000100 : OUT <= 1;  //160 / 132 = 1
    16'b10100000_10000101 : OUT <= 1;  //160 / 133 = 1
    16'b10100000_10000110 : OUT <= 1;  //160 / 134 = 1
    16'b10100000_10000111 : OUT <= 1;  //160 / 135 = 1
    16'b10100000_10001000 : OUT <= 1;  //160 / 136 = 1
    16'b10100000_10001001 : OUT <= 1;  //160 / 137 = 1
    16'b10100000_10001010 : OUT <= 1;  //160 / 138 = 1
    16'b10100000_10001011 : OUT <= 1;  //160 / 139 = 1
    16'b10100000_10001100 : OUT <= 1;  //160 / 140 = 1
    16'b10100000_10001101 : OUT <= 1;  //160 / 141 = 1
    16'b10100000_10001110 : OUT <= 1;  //160 / 142 = 1
    16'b10100000_10001111 : OUT <= 1;  //160 / 143 = 1
    16'b10100000_10010000 : OUT <= 1;  //160 / 144 = 1
    16'b10100000_10010001 : OUT <= 1;  //160 / 145 = 1
    16'b10100000_10010010 : OUT <= 1;  //160 / 146 = 1
    16'b10100000_10010011 : OUT <= 1;  //160 / 147 = 1
    16'b10100000_10010100 : OUT <= 1;  //160 / 148 = 1
    16'b10100000_10010101 : OUT <= 1;  //160 / 149 = 1
    16'b10100000_10010110 : OUT <= 1;  //160 / 150 = 1
    16'b10100000_10010111 : OUT <= 1;  //160 / 151 = 1
    16'b10100000_10011000 : OUT <= 1;  //160 / 152 = 1
    16'b10100000_10011001 : OUT <= 1;  //160 / 153 = 1
    16'b10100000_10011010 : OUT <= 1;  //160 / 154 = 1
    16'b10100000_10011011 : OUT <= 1;  //160 / 155 = 1
    16'b10100000_10011100 : OUT <= 1;  //160 / 156 = 1
    16'b10100000_10011101 : OUT <= 1;  //160 / 157 = 1
    16'b10100000_10011110 : OUT <= 1;  //160 / 158 = 1
    16'b10100000_10011111 : OUT <= 1;  //160 / 159 = 1
    16'b10100000_10100000 : OUT <= 1;  //160 / 160 = 1
    16'b10100000_10100001 : OUT <= 0;  //160 / 161 = 0
    16'b10100000_10100010 : OUT <= 0;  //160 / 162 = 0
    16'b10100000_10100011 : OUT <= 0;  //160 / 163 = 0
    16'b10100000_10100100 : OUT <= 0;  //160 / 164 = 0
    16'b10100000_10100101 : OUT <= 0;  //160 / 165 = 0
    16'b10100000_10100110 : OUT <= 0;  //160 / 166 = 0
    16'b10100000_10100111 : OUT <= 0;  //160 / 167 = 0
    16'b10100000_10101000 : OUT <= 0;  //160 / 168 = 0
    16'b10100000_10101001 : OUT <= 0;  //160 / 169 = 0
    16'b10100000_10101010 : OUT <= 0;  //160 / 170 = 0
    16'b10100000_10101011 : OUT <= 0;  //160 / 171 = 0
    16'b10100000_10101100 : OUT <= 0;  //160 / 172 = 0
    16'b10100000_10101101 : OUT <= 0;  //160 / 173 = 0
    16'b10100000_10101110 : OUT <= 0;  //160 / 174 = 0
    16'b10100000_10101111 : OUT <= 0;  //160 / 175 = 0
    16'b10100000_10110000 : OUT <= 0;  //160 / 176 = 0
    16'b10100000_10110001 : OUT <= 0;  //160 / 177 = 0
    16'b10100000_10110010 : OUT <= 0;  //160 / 178 = 0
    16'b10100000_10110011 : OUT <= 0;  //160 / 179 = 0
    16'b10100000_10110100 : OUT <= 0;  //160 / 180 = 0
    16'b10100000_10110101 : OUT <= 0;  //160 / 181 = 0
    16'b10100000_10110110 : OUT <= 0;  //160 / 182 = 0
    16'b10100000_10110111 : OUT <= 0;  //160 / 183 = 0
    16'b10100000_10111000 : OUT <= 0;  //160 / 184 = 0
    16'b10100000_10111001 : OUT <= 0;  //160 / 185 = 0
    16'b10100000_10111010 : OUT <= 0;  //160 / 186 = 0
    16'b10100000_10111011 : OUT <= 0;  //160 / 187 = 0
    16'b10100000_10111100 : OUT <= 0;  //160 / 188 = 0
    16'b10100000_10111101 : OUT <= 0;  //160 / 189 = 0
    16'b10100000_10111110 : OUT <= 0;  //160 / 190 = 0
    16'b10100000_10111111 : OUT <= 0;  //160 / 191 = 0
    16'b10100000_11000000 : OUT <= 0;  //160 / 192 = 0
    16'b10100000_11000001 : OUT <= 0;  //160 / 193 = 0
    16'b10100000_11000010 : OUT <= 0;  //160 / 194 = 0
    16'b10100000_11000011 : OUT <= 0;  //160 / 195 = 0
    16'b10100000_11000100 : OUT <= 0;  //160 / 196 = 0
    16'b10100000_11000101 : OUT <= 0;  //160 / 197 = 0
    16'b10100000_11000110 : OUT <= 0;  //160 / 198 = 0
    16'b10100000_11000111 : OUT <= 0;  //160 / 199 = 0
    16'b10100000_11001000 : OUT <= 0;  //160 / 200 = 0
    16'b10100000_11001001 : OUT <= 0;  //160 / 201 = 0
    16'b10100000_11001010 : OUT <= 0;  //160 / 202 = 0
    16'b10100000_11001011 : OUT <= 0;  //160 / 203 = 0
    16'b10100000_11001100 : OUT <= 0;  //160 / 204 = 0
    16'b10100000_11001101 : OUT <= 0;  //160 / 205 = 0
    16'b10100000_11001110 : OUT <= 0;  //160 / 206 = 0
    16'b10100000_11001111 : OUT <= 0;  //160 / 207 = 0
    16'b10100000_11010000 : OUT <= 0;  //160 / 208 = 0
    16'b10100000_11010001 : OUT <= 0;  //160 / 209 = 0
    16'b10100000_11010010 : OUT <= 0;  //160 / 210 = 0
    16'b10100000_11010011 : OUT <= 0;  //160 / 211 = 0
    16'b10100000_11010100 : OUT <= 0;  //160 / 212 = 0
    16'b10100000_11010101 : OUT <= 0;  //160 / 213 = 0
    16'b10100000_11010110 : OUT <= 0;  //160 / 214 = 0
    16'b10100000_11010111 : OUT <= 0;  //160 / 215 = 0
    16'b10100000_11011000 : OUT <= 0;  //160 / 216 = 0
    16'b10100000_11011001 : OUT <= 0;  //160 / 217 = 0
    16'b10100000_11011010 : OUT <= 0;  //160 / 218 = 0
    16'b10100000_11011011 : OUT <= 0;  //160 / 219 = 0
    16'b10100000_11011100 : OUT <= 0;  //160 / 220 = 0
    16'b10100000_11011101 : OUT <= 0;  //160 / 221 = 0
    16'b10100000_11011110 : OUT <= 0;  //160 / 222 = 0
    16'b10100000_11011111 : OUT <= 0;  //160 / 223 = 0
    16'b10100000_11100000 : OUT <= 0;  //160 / 224 = 0
    16'b10100000_11100001 : OUT <= 0;  //160 / 225 = 0
    16'b10100000_11100010 : OUT <= 0;  //160 / 226 = 0
    16'b10100000_11100011 : OUT <= 0;  //160 / 227 = 0
    16'b10100000_11100100 : OUT <= 0;  //160 / 228 = 0
    16'b10100000_11100101 : OUT <= 0;  //160 / 229 = 0
    16'b10100000_11100110 : OUT <= 0;  //160 / 230 = 0
    16'b10100000_11100111 : OUT <= 0;  //160 / 231 = 0
    16'b10100000_11101000 : OUT <= 0;  //160 / 232 = 0
    16'b10100000_11101001 : OUT <= 0;  //160 / 233 = 0
    16'b10100000_11101010 : OUT <= 0;  //160 / 234 = 0
    16'b10100000_11101011 : OUT <= 0;  //160 / 235 = 0
    16'b10100000_11101100 : OUT <= 0;  //160 / 236 = 0
    16'b10100000_11101101 : OUT <= 0;  //160 / 237 = 0
    16'b10100000_11101110 : OUT <= 0;  //160 / 238 = 0
    16'b10100000_11101111 : OUT <= 0;  //160 / 239 = 0
    16'b10100000_11110000 : OUT <= 0;  //160 / 240 = 0
    16'b10100000_11110001 : OUT <= 0;  //160 / 241 = 0
    16'b10100000_11110010 : OUT <= 0;  //160 / 242 = 0
    16'b10100000_11110011 : OUT <= 0;  //160 / 243 = 0
    16'b10100000_11110100 : OUT <= 0;  //160 / 244 = 0
    16'b10100000_11110101 : OUT <= 0;  //160 / 245 = 0
    16'b10100000_11110110 : OUT <= 0;  //160 / 246 = 0
    16'b10100000_11110111 : OUT <= 0;  //160 / 247 = 0
    16'b10100000_11111000 : OUT <= 0;  //160 / 248 = 0
    16'b10100000_11111001 : OUT <= 0;  //160 / 249 = 0
    16'b10100000_11111010 : OUT <= 0;  //160 / 250 = 0
    16'b10100000_11111011 : OUT <= 0;  //160 / 251 = 0
    16'b10100000_11111100 : OUT <= 0;  //160 / 252 = 0
    16'b10100000_11111101 : OUT <= 0;  //160 / 253 = 0
    16'b10100000_11111110 : OUT <= 0;  //160 / 254 = 0
    16'b10100000_11111111 : OUT <= 0;  //160 / 255 = 0
    16'b10100001_00000000 : OUT <= 0;  //161 / 0 = 0
    16'b10100001_00000001 : OUT <= 161;  //161 / 1 = 161
    16'b10100001_00000010 : OUT <= 80;  //161 / 2 = 80
    16'b10100001_00000011 : OUT <= 53;  //161 / 3 = 53
    16'b10100001_00000100 : OUT <= 40;  //161 / 4 = 40
    16'b10100001_00000101 : OUT <= 32;  //161 / 5 = 32
    16'b10100001_00000110 : OUT <= 26;  //161 / 6 = 26
    16'b10100001_00000111 : OUT <= 23;  //161 / 7 = 23
    16'b10100001_00001000 : OUT <= 20;  //161 / 8 = 20
    16'b10100001_00001001 : OUT <= 17;  //161 / 9 = 17
    16'b10100001_00001010 : OUT <= 16;  //161 / 10 = 16
    16'b10100001_00001011 : OUT <= 14;  //161 / 11 = 14
    16'b10100001_00001100 : OUT <= 13;  //161 / 12 = 13
    16'b10100001_00001101 : OUT <= 12;  //161 / 13 = 12
    16'b10100001_00001110 : OUT <= 11;  //161 / 14 = 11
    16'b10100001_00001111 : OUT <= 10;  //161 / 15 = 10
    16'b10100001_00010000 : OUT <= 10;  //161 / 16 = 10
    16'b10100001_00010001 : OUT <= 9;  //161 / 17 = 9
    16'b10100001_00010010 : OUT <= 8;  //161 / 18 = 8
    16'b10100001_00010011 : OUT <= 8;  //161 / 19 = 8
    16'b10100001_00010100 : OUT <= 8;  //161 / 20 = 8
    16'b10100001_00010101 : OUT <= 7;  //161 / 21 = 7
    16'b10100001_00010110 : OUT <= 7;  //161 / 22 = 7
    16'b10100001_00010111 : OUT <= 7;  //161 / 23 = 7
    16'b10100001_00011000 : OUT <= 6;  //161 / 24 = 6
    16'b10100001_00011001 : OUT <= 6;  //161 / 25 = 6
    16'b10100001_00011010 : OUT <= 6;  //161 / 26 = 6
    16'b10100001_00011011 : OUT <= 5;  //161 / 27 = 5
    16'b10100001_00011100 : OUT <= 5;  //161 / 28 = 5
    16'b10100001_00011101 : OUT <= 5;  //161 / 29 = 5
    16'b10100001_00011110 : OUT <= 5;  //161 / 30 = 5
    16'b10100001_00011111 : OUT <= 5;  //161 / 31 = 5
    16'b10100001_00100000 : OUT <= 5;  //161 / 32 = 5
    16'b10100001_00100001 : OUT <= 4;  //161 / 33 = 4
    16'b10100001_00100010 : OUT <= 4;  //161 / 34 = 4
    16'b10100001_00100011 : OUT <= 4;  //161 / 35 = 4
    16'b10100001_00100100 : OUT <= 4;  //161 / 36 = 4
    16'b10100001_00100101 : OUT <= 4;  //161 / 37 = 4
    16'b10100001_00100110 : OUT <= 4;  //161 / 38 = 4
    16'b10100001_00100111 : OUT <= 4;  //161 / 39 = 4
    16'b10100001_00101000 : OUT <= 4;  //161 / 40 = 4
    16'b10100001_00101001 : OUT <= 3;  //161 / 41 = 3
    16'b10100001_00101010 : OUT <= 3;  //161 / 42 = 3
    16'b10100001_00101011 : OUT <= 3;  //161 / 43 = 3
    16'b10100001_00101100 : OUT <= 3;  //161 / 44 = 3
    16'b10100001_00101101 : OUT <= 3;  //161 / 45 = 3
    16'b10100001_00101110 : OUT <= 3;  //161 / 46 = 3
    16'b10100001_00101111 : OUT <= 3;  //161 / 47 = 3
    16'b10100001_00110000 : OUT <= 3;  //161 / 48 = 3
    16'b10100001_00110001 : OUT <= 3;  //161 / 49 = 3
    16'b10100001_00110010 : OUT <= 3;  //161 / 50 = 3
    16'b10100001_00110011 : OUT <= 3;  //161 / 51 = 3
    16'b10100001_00110100 : OUT <= 3;  //161 / 52 = 3
    16'b10100001_00110101 : OUT <= 3;  //161 / 53 = 3
    16'b10100001_00110110 : OUT <= 2;  //161 / 54 = 2
    16'b10100001_00110111 : OUT <= 2;  //161 / 55 = 2
    16'b10100001_00111000 : OUT <= 2;  //161 / 56 = 2
    16'b10100001_00111001 : OUT <= 2;  //161 / 57 = 2
    16'b10100001_00111010 : OUT <= 2;  //161 / 58 = 2
    16'b10100001_00111011 : OUT <= 2;  //161 / 59 = 2
    16'b10100001_00111100 : OUT <= 2;  //161 / 60 = 2
    16'b10100001_00111101 : OUT <= 2;  //161 / 61 = 2
    16'b10100001_00111110 : OUT <= 2;  //161 / 62 = 2
    16'b10100001_00111111 : OUT <= 2;  //161 / 63 = 2
    16'b10100001_01000000 : OUT <= 2;  //161 / 64 = 2
    16'b10100001_01000001 : OUT <= 2;  //161 / 65 = 2
    16'b10100001_01000010 : OUT <= 2;  //161 / 66 = 2
    16'b10100001_01000011 : OUT <= 2;  //161 / 67 = 2
    16'b10100001_01000100 : OUT <= 2;  //161 / 68 = 2
    16'b10100001_01000101 : OUT <= 2;  //161 / 69 = 2
    16'b10100001_01000110 : OUT <= 2;  //161 / 70 = 2
    16'b10100001_01000111 : OUT <= 2;  //161 / 71 = 2
    16'b10100001_01001000 : OUT <= 2;  //161 / 72 = 2
    16'b10100001_01001001 : OUT <= 2;  //161 / 73 = 2
    16'b10100001_01001010 : OUT <= 2;  //161 / 74 = 2
    16'b10100001_01001011 : OUT <= 2;  //161 / 75 = 2
    16'b10100001_01001100 : OUT <= 2;  //161 / 76 = 2
    16'b10100001_01001101 : OUT <= 2;  //161 / 77 = 2
    16'b10100001_01001110 : OUT <= 2;  //161 / 78 = 2
    16'b10100001_01001111 : OUT <= 2;  //161 / 79 = 2
    16'b10100001_01010000 : OUT <= 2;  //161 / 80 = 2
    16'b10100001_01010001 : OUT <= 1;  //161 / 81 = 1
    16'b10100001_01010010 : OUT <= 1;  //161 / 82 = 1
    16'b10100001_01010011 : OUT <= 1;  //161 / 83 = 1
    16'b10100001_01010100 : OUT <= 1;  //161 / 84 = 1
    16'b10100001_01010101 : OUT <= 1;  //161 / 85 = 1
    16'b10100001_01010110 : OUT <= 1;  //161 / 86 = 1
    16'b10100001_01010111 : OUT <= 1;  //161 / 87 = 1
    16'b10100001_01011000 : OUT <= 1;  //161 / 88 = 1
    16'b10100001_01011001 : OUT <= 1;  //161 / 89 = 1
    16'b10100001_01011010 : OUT <= 1;  //161 / 90 = 1
    16'b10100001_01011011 : OUT <= 1;  //161 / 91 = 1
    16'b10100001_01011100 : OUT <= 1;  //161 / 92 = 1
    16'b10100001_01011101 : OUT <= 1;  //161 / 93 = 1
    16'b10100001_01011110 : OUT <= 1;  //161 / 94 = 1
    16'b10100001_01011111 : OUT <= 1;  //161 / 95 = 1
    16'b10100001_01100000 : OUT <= 1;  //161 / 96 = 1
    16'b10100001_01100001 : OUT <= 1;  //161 / 97 = 1
    16'b10100001_01100010 : OUT <= 1;  //161 / 98 = 1
    16'b10100001_01100011 : OUT <= 1;  //161 / 99 = 1
    16'b10100001_01100100 : OUT <= 1;  //161 / 100 = 1
    16'b10100001_01100101 : OUT <= 1;  //161 / 101 = 1
    16'b10100001_01100110 : OUT <= 1;  //161 / 102 = 1
    16'b10100001_01100111 : OUT <= 1;  //161 / 103 = 1
    16'b10100001_01101000 : OUT <= 1;  //161 / 104 = 1
    16'b10100001_01101001 : OUT <= 1;  //161 / 105 = 1
    16'b10100001_01101010 : OUT <= 1;  //161 / 106 = 1
    16'b10100001_01101011 : OUT <= 1;  //161 / 107 = 1
    16'b10100001_01101100 : OUT <= 1;  //161 / 108 = 1
    16'b10100001_01101101 : OUT <= 1;  //161 / 109 = 1
    16'b10100001_01101110 : OUT <= 1;  //161 / 110 = 1
    16'b10100001_01101111 : OUT <= 1;  //161 / 111 = 1
    16'b10100001_01110000 : OUT <= 1;  //161 / 112 = 1
    16'b10100001_01110001 : OUT <= 1;  //161 / 113 = 1
    16'b10100001_01110010 : OUT <= 1;  //161 / 114 = 1
    16'b10100001_01110011 : OUT <= 1;  //161 / 115 = 1
    16'b10100001_01110100 : OUT <= 1;  //161 / 116 = 1
    16'b10100001_01110101 : OUT <= 1;  //161 / 117 = 1
    16'b10100001_01110110 : OUT <= 1;  //161 / 118 = 1
    16'b10100001_01110111 : OUT <= 1;  //161 / 119 = 1
    16'b10100001_01111000 : OUT <= 1;  //161 / 120 = 1
    16'b10100001_01111001 : OUT <= 1;  //161 / 121 = 1
    16'b10100001_01111010 : OUT <= 1;  //161 / 122 = 1
    16'b10100001_01111011 : OUT <= 1;  //161 / 123 = 1
    16'b10100001_01111100 : OUT <= 1;  //161 / 124 = 1
    16'b10100001_01111101 : OUT <= 1;  //161 / 125 = 1
    16'b10100001_01111110 : OUT <= 1;  //161 / 126 = 1
    16'b10100001_01111111 : OUT <= 1;  //161 / 127 = 1
    16'b10100001_10000000 : OUT <= 1;  //161 / 128 = 1
    16'b10100001_10000001 : OUT <= 1;  //161 / 129 = 1
    16'b10100001_10000010 : OUT <= 1;  //161 / 130 = 1
    16'b10100001_10000011 : OUT <= 1;  //161 / 131 = 1
    16'b10100001_10000100 : OUT <= 1;  //161 / 132 = 1
    16'b10100001_10000101 : OUT <= 1;  //161 / 133 = 1
    16'b10100001_10000110 : OUT <= 1;  //161 / 134 = 1
    16'b10100001_10000111 : OUT <= 1;  //161 / 135 = 1
    16'b10100001_10001000 : OUT <= 1;  //161 / 136 = 1
    16'b10100001_10001001 : OUT <= 1;  //161 / 137 = 1
    16'b10100001_10001010 : OUT <= 1;  //161 / 138 = 1
    16'b10100001_10001011 : OUT <= 1;  //161 / 139 = 1
    16'b10100001_10001100 : OUT <= 1;  //161 / 140 = 1
    16'b10100001_10001101 : OUT <= 1;  //161 / 141 = 1
    16'b10100001_10001110 : OUT <= 1;  //161 / 142 = 1
    16'b10100001_10001111 : OUT <= 1;  //161 / 143 = 1
    16'b10100001_10010000 : OUT <= 1;  //161 / 144 = 1
    16'b10100001_10010001 : OUT <= 1;  //161 / 145 = 1
    16'b10100001_10010010 : OUT <= 1;  //161 / 146 = 1
    16'b10100001_10010011 : OUT <= 1;  //161 / 147 = 1
    16'b10100001_10010100 : OUT <= 1;  //161 / 148 = 1
    16'b10100001_10010101 : OUT <= 1;  //161 / 149 = 1
    16'b10100001_10010110 : OUT <= 1;  //161 / 150 = 1
    16'b10100001_10010111 : OUT <= 1;  //161 / 151 = 1
    16'b10100001_10011000 : OUT <= 1;  //161 / 152 = 1
    16'b10100001_10011001 : OUT <= 1;  //161 / 153 = 1
    16'b10100001_10011010 : OUT <= 1;  //161 / 154 = 1
    16'b10100001_10011011 : OUT <= 1;  //161 / 155 = 1
    16'b10100001_10011100 : OUT <= 1;  //161 / 156 = 1
    16'b10100001_10011101 : OUT <= 1;  //161 / 157 = 1
    16'b10100001_10011110 : OUT <= 1;  //161 / 158 = 1
    16'b10100001_10011111 : OUT <= 1;  //161 / 159 = 1
    16'b10100001_10100000 : OUT <= 1;  //161 / 160 = 1
    16'b10100001_10100001 : OUT <= 1;  //161 / 161 = 1
    16'b10100001_10100010 : OUT <= 0;  //161 / 162 = 0
    16'b10100001_10100011 : OUT <= 0;  //161 / 163 = 0
    16'b10100001_10100100 : OUT <= 0;  //161 / 164 = 0
    16'b10100001_10100101 : OUT <= 0;  //161 / 165 = 0
    16'b10100001_10100110 : OUT <= 0;  //161 / 166 = 0
    16'b10100001_10100111 : OUT <= 0;  //161 / 167 = 0
    16'b10100001_10101000 : OUT <= 0;  //161 / 168 = 0
    16'b10100001_10101001 : OUT <= 0;  //161 / 169 = 0
    16'b10100001_10101010 : OUT <= 0;  //161 / 170 = 0
    16'b10100001_10101011 : OUT <= 0;  //161 / 171 = 0
    16'b10100001_10101100 : OUT <= 0;  //161 / 172 = 0
    16'b10100001_10101101 : OUT <= 0;  //161 / 173 = 0
    16'b10100001_10101110 : OUT <= 0;  //161 / 174 = 0
    16'b10100001_10101111 : OUT <= 0;  //161 / 175 = 0
    16'b10100001_10110000 : OUT <= 0;  //161 / 176 = 0
    16'b10100001_10110001 : OUT <= 0;  //161 / 177 = 0
    16'b10100001_10110010 : OUT <= 0;  //161 / 178 = 0
    16'b10100001_10110011 : OUT <= 0;  //161 / 179 = 0
    16'b10100001_10110100 : OUT <= 0;  //161 / 180 = 0
    16'b10100001_10110101 : OUT <= 0;  //161 / 181 = 0
    16'b10100001_10110110 : OUT <= 0;  //161 / 182 = 0
    16'b10100001_10110111 : OUT <= 0;  //161 / 183 = 0
    16'b10100001_10111000 : OUT <= 0;  //161 / 184 = 0
    16'b10100001_10111001 : OUT <= 0;  //161 / 185 = 0
    16'b10100001_10111010 : OUT <= 0;  //161 / 186 = 0
    16'b10100001_10111011 : OUT <= 0;  //161 / 187 = 0
    16'b10100001_10111100 : OUT <= 0;  //161 / 188 = 0
    16'b10100001_10111101 : OUT <= 0;  //161 / 189 = 0
    16'b10100001_10111110 : OUT <= 0;  //161 / 190 = 0
    16'b10100001_10111111 : OUT <= 0;  //161 / 191 = 0
    16'b10100001_11000000 : OUT <= 0;  //161 / 192 = 0
    16'b10100001_11000001 : OUT <= 0;  //161 / 193 = 0
    16'b10100001_11000010 : OUT <= 0;  //161 / 194 = 0
    16'b10100001_11000011 : OUT <= 0;  //161 / 195 = 0
    16'b10100001_11000100 : OUT <= 0;  //161 / 196 = 0
    16'b10100001_11000101 : OUT <= 0;  //161 / 197 = 0
    16'b10100001_11000110 : OUT <= 0;  //161 / 198 = 0
    16'b10100001_11000111 : OUT <= 0;  //161 / 199 = 0
    16'b10100001_11001000 : OUT <= 0;  //161 / 200 = 0
    16'b10100001_11001001 : OUT <= 0;  //161 / 201 = 0
    16'b10100001_11001010 : OUT <= 0;  //161 / 202 = 0
    16'b10100001_11001011 : OUT <= 0;  //161 / 203 = 0
    16'b10100001_11001100 : OUT <= 0;  //161 / 204 = 0
    16'b10100001_11001101 : OUT <= 0;  //161 / 205 = 0
    16'b10100001_11001110 : OUT <= 0;  //161 / 206 = 0
    16'b10100001_11001111 : OUT <= 0;  //161 / 207 = 0
    16'b10100001_11010000 : OUT <= 0;  //161 / 208 = 0
    16'b10100001_11010001 : OUT <= 0;  //161 / 209 = 0
    16'b10100001_11010010 : OUT <= 0;  //161 / 210 = 0
    16'b10100001_11010011 : OUT <= 0;  //161 / 211 = 0
    16'b10100001_11010100 : OUT <= 0;  //161 / 212 = 0
    16'b10100001_11010101 : OUT <= 0;  //161 / 213 = 0
    16'b10100001_11010110 : OUT <= 0;  //161 / 214 = 0
    16'b10100001_11010111 : OUT <= 0;  //161 / 215 = 0
    16'b10100001_11011000 : OUT <= 0;  //161 / 216 = 0
    16'b10100001_11011001 : OUT <= 0;  //161 / 217 = 0
    16'b10100001_11011010 : OUT <= 0;  //161 / 218 = 0
    16'b10100001_11011011 : OUT <= 0;  //161 / 219 = 0
    16'b10100001_11011100 : OUT <= 0;  //161 / 220 = 0
    16'b10100001_11011101 : OUT <= 0;  //161 / 221 = 0
    16'b10100001_11011110 : OUT <= 0;  //161 / 222 = 0
    16'b10100001_11011111 : OUT <= 0;  //161 / 223 = 0
    16'b10100001_11100000 : OUT <= 0;  //161 / 224 = 0
    16'b10100001_11100001 : OUT <= 0;  //161 / 225 = 0
    16'b10100001_11100010 : OUT <= 0;  //161 / 226 = 0
    16'b10100001_11100011 : OUT <= 0;  //161 / 227 = 0
    16'b10100001_11100100 : OUT <= 0;  //161 / 228 = 0
    16'b10100001_11100101 : OUT <= 0;  //161 / 229 = 0
    16'b10100001_11100110 : OUT <= 0;  //161 / 230 = 0
    16'b10100001_11100111 : OUT <= 0;  //161 / 231 = 0
    16'b10100001_11101000 : OUT <= 0;  //161 / 232 = 0
    16'b10100001_11101001 : OUT <= 0;  //161 / 233 = 0
    16'b10100001_11101010 : OUT <= 0;  //161 / 234 = 0
    16'b10100001_11101011 : OUT <= 0;  //161 / 235 = 0
    16'b10100001_11101100 : OUT <= 0;  //161 / 236 = 0
    16'b10100001_11101101 : OUT <= 0;  //161 / 237 = 0
    16'b10100001_11101110 : OUT <= 0;  //161 / 238 = 0
    16'b10100001_11101111 : OUT <= 0;  //161 / 239 = 0
    16'b10100001_11110000 : OUT <= 0;  //161 / 240 = 0
    16'b10100001_11110001 : OUT <= 0;  //161 / 241 = 0
    16'b10100001_11110010 : OUT <= 0;  //161 / 242 = 0
    16'b10100001_11110011 : OUT <= 0;  //161 / 243 = 0
    16'b10100001_11110100 : OUT <= 0;  //161 / 244 = 0
    16'b10100001_11110101 : OUT <= 0;  //161 / 245 = 0
    16'b10100001_11110110 : OUT <= 0;  //161 / 246 = 0
    16'b10100001_11110111 : OUT <= 0;  //161 / 247 = 0
    16'b10100001_11111000 : OUT <= 0;  //161 / 248 = 0
    16'b10100001_11111001 : OUT <= 0;  //161 / 249 = 0
    16'b10100001_11111010 : OUT <= 0;  //161 / 250 = 0
    16'b10100001_11111011 : OUT <= 0;  //161 / 251 = 0
    16'b10100001_11111100 : OUT <= 0;  //161 / 252 = 0
    16'b10100001_11111101 : OUT <= 0;  //161 / 253 = 0
    16'b10100001_11111110 : OUT <= 0;  //161 / 254 = 0
    16'b10100001_11111111 : OUT <= 0;  //161 / 255 = 0
    16'b10100010_00000000 : OUT <= 0;  //162 / 0 = 0
    16'b10100010_00000001 : OUT <= 162;  //162 / 1 = 162
    16'b10100010_00000010 : OUT <= 81;  //162 / 2 = 81
    16'b10100010_00000011 : OUT <= 54;  //162 / 3 = 54
    16'b10100010_00000100 : OUT <= 40;  //162 / 4 = 40
    16'b10100010_00000101 : OUT <= 32;  //162 / 5 = 32
    16'b10100010_00000110 : OUT <= 27;  //162 / 6 = 27
    16'b10100010_00000111 : OUT <= 23;  //162 / 7 = 23
    16'b10100010_00001000 : OUT <= 20;  //162 / 8 = 20
    16'b10100010_00001001 : OUT <= 18;  //162 / 9 = 18
    16'b10100010_00001010 : OUT <= 16;  //162 / 10 = 16
    16'b10100010_00001011 : OUT <= 14;  //162 / 11 = 14
    16'b10100010_00001100 : OUT <= 13;  //162 / 12 = 13
    16'b10100010_00001101 : OUT <= 12;  //162 / 13 = 12
    16'b10100010_00001110 : OUT <= 11;  //162 / 14 = 11
    16'b10100010_00001111 : OUT <= 10;  //162 / 15 = 10
    16'b10100010_00010000 : OUT <= 10;  //162 / 16 = 10
    16'b10100010_00010001 : OUT <= 9;  //162 / 17 = 9
    16'b10100010_00010010 : OUT <= 9;  //162 / 18 = 9
    16'b10100010_00010011 : OUT <= 8;  //162 / 19 = 8
    16'b10100010_00010100 : OUT <= 8;  //162 / 20 = 8
    16'b10100010_00010101 : OUT <= 7;  //162 / 21 = 7
    16'b10100010_00010110 : OUT <= 7;  //162 / 22 = 7
    16'b10100010_00010111 : OUT <= 7;  //162 / 23 = 7
    16'b10100010_00011000 : OUT <= 6;  //162 / 24 = 6
    16'b10100010_00011001 : OUT <= 6;  //162 / 25 = 6
    16'b10100010_00011010 : OUT <= 6;  //162 / 26 = 6
    16'b10100010_00011011 : OUT <= 6;  //162 / 27 = 6
    16'b10100010_00011100 : OUT <= 5;  //162 / 28 = 5
    16'b10100010_00011101 : OUT <= 5;  //162 / 29 = 5
    16'b10100010_00011110 : OUT <= 5;  //162 / 30 = 5
    16'b10100010_00011111 : OUT <= 5;  //162 / 31 = 5
    16'b10100010_00100000 : OUT <= 5;  //162 / 32 = 5
    16'b10100010_00100001 : OUT <= 4;  //162 / 33 = 4
    16'b10100010_00100010 : OUT <= 4;  //162 / 34 = 4
    16'b10100010_00100011 : OUT <= 4;  //162 / 35 = 4
    16'b10100010_00100100 : OUT <= 4;  //162 / 36 = 4
    16'b10100010_00100101 : OUT <= 4;  //162 / 37 = 4
    16'b10100010_00100110 : OUT <= 4;  //162 / 38 = 4
    16'b10100010_00100111 : OUT <= 4;  //162 / 39 = 4
    16'b10100010_00101000 : OUT <= 4;  //162 / 40 = 4
    16'b10100010_00101001 : OUT <= 3;  //162 / 41 = 3
    16'b10100010_00101010 : OUT <= 3;  //162 / 42 = 3
    16'b10100010_00101011 : OUT <= 3;  //162 / 43 = 3
    16'b10100010_00101100 : OUT <= 3;  //162 / 44 = 3
    16'b10100010_00101101 : OUT <= 3;  //162 / 45 = 3
    16'b10100010_00101110 : OUT <= 3;  //162 / 46 = 3
    16'b10100010_00101111 : OUT <= 3;  //162 / 47 = 3
    16'b10100010_00110000 : OUT <= 3;  //162 / 48 = 3
    16'b10100010_00110001 : OUT <= 3;  //162 / 49 = 3
    16'b10100010_00110010 : OUT <= 3;  //162 / 50 = 3
    16'b10100010_00110011 : OUT <= 3;  //162 / 51 = 3
    16'b10100010_00110100 : OUT <= 3;  //162 / 52 = 3
    16'b10100010_00110101 : OUT <= 3;  //162 / 53 = 3
    16'b10100010_00110110 : OUT <= 3;  //162 / 54 = 3
    16'b10100010_00110111 : OUT <= 2;  //162 / 55 = 2
    16'b10100010_00111000 : OUT <= 2;  //162 / 56 = 2
    16'b10100010_00111001 : OUT <= 2;  //162 / 57 = 2
    16'b10100010_00111010 : OUT <= 2;  //162 / 58 = 2
    16'b10100010_00111011 : OUT <= 2;  //162 / 59 = 2
    16'b10100010_00111100 : OUT <= 2;  //162 / 60 = 2
    16'b10100010_00111101 : OUT <= 2;  //162 / 61 = 2
    16'b10100010_00111110 : OUT <= 2;  //162 / 62 = 2
    16'b10100010_00111111 : OUT <= 2;  //162 / 63 = 2
    16'b10100010_01000000 : OUT <= 2;  //162 / 64 = 2
    16'b10100010_01000001 : OUT <= 2;  //162 / 65 = 2
    16'b10100010_01000010 : OUT <= 2;  //162 / 66 = 2
    16'b10100010_01000011 : OUT <= 2;  //162 / 67 = 2
    16'b10100010_01000100 : OUT <= 2;  //162 / 68 = 2
    16'b10100010_01000101 : OUT <= 2;  //162 / 69 = 2
    16'b10100010_01000110 : OUT <= 2;  //162 / 70 = 2
    16'b10100010_01000111 : OUT <= 2;  //162 / 71 = 2
    16'b10100010_01001000 : OUT <= 2;  //162 / 72 = 2
    16'b10100010_01001001 : OUT <= 2;  //162 / 73 = 2
    16'b10100010_01001010 : OUT <= 2;  //162 / 74 = 2
    16'b10100010_01001011 : OUT <= 2;  //162 / 75 = 2
    16'b10100010_01001100 : OUT <= 2;  //162 / 76 = 2
    16'b10100010_01001101 : OUT <= 2;  //162 / 77 = 2
    16'b10100010_01001110 : OUT <= 2;  //162 / 78 = 2
    16'b10100010_01001111 : OUT <= 2;  //162 / 79 = 2
    16'b10100010_01010000 : OUT <= 2;  //162 / 80 = 2
    16'b10100010_01010001 : OUT <= 2;  //162 / 81 = 2
    16'b10100010_01010010 : OUT <= 1;  //162 / 82 = 1
    16'b10100010_01010011 : OUT <= 1;  //162 / 83 = 1
    16'b10100010_01010100 : OUT <= 1;  //162 / 84 = 1
    16'b10100010_01010101 : OUT <= 1;  //162 / 85 = 1
    16'b10100010_01010110 : OUT <= 1;  //162 / 86 = 1
    16'b10100010_01010111 : OUT <= 1;  //162 / 87 = 1
    16'b10100010_01011000 : OUT <= 1;  //162 / 88 = 1
    16'b10100010_01011001 : OUT <= 1;  //162 / 89 = 1
    16'b10100010_01011010 : OUT <= 1;  //162 / 90 = 1
    16'b10100010_01011011 : OUT <= 1;  //162 / 91 = 1
    16'b10100010_01011100 : OUT <= 1;  //162 / 92 = 1
    16'b10100010_01011101 : OUT <= 1;  //162 / 93 = 1
    16'b10100010_01011110 : OUT <= 1;  //162 / 94 = 1
    16'b10100010_01011111 : OUT <= 1;  //162 / 95 = 1
    16'b10100010_01100000 : OUT <= 1;  //162 / 96 = 1
    16'b10100010_01100001 : OUT <= 1;  //162 / 97 = 1
    16'b10100010_01100010 : OUT <= 1;  //162 / 98 = 1
    16'b10100010_01100011 : OUT <= 1;  //162 / 99 = 1
    16'b10100010_01100100 : OUT <= 1;  //162 / 100 = 1
    16'b10100010_01100101 : OUT <= 1;  //162 / 101 = 1
    16'b10100010_01100110 : OUT <= 1;  //162 / 102 = 1
    16'b10100010_01100111 : OUT <= 1;  //162 / 103 = 1
    16'b10100010_01101000 : OUT <= 1;  //162 / 104 = 1
    16'b10100010_01101001 : OUT <= 1;  //162 / 105 = 1
    16'b10100010_01101010 : OUT <= 1;  //162 / 106 = 1
    16'b10100010_01101011 : OUT <= 1;  //162 / 107 = 1
    16'b10100010_01101100 : OUT <= 1;  //162 / 108 = 1
    16'b10100010_01101101 : OUT <= 1;  //162 / 109 = 1
    16'b10100010_01101110 : OUT <= 1;  //162 / 110 = 1
    16'b10100010_01101111 : OUT <= 1;  //162 / 111 = 1
    16'b10100010_01110000 : OUT <= 1;  //162 / 112 = 1
    16'b10100010_01110001 : OUT <= 1;  //162 / 113 = 1
    16'b10100010_01110010 : OUT <= 1;  //162 / 114 = 1
    16'b10100010_01110011 : OUT <= 1;  //162 / 115 = 1
    16'b10100010_01110100 : OUT <= 1;  //162 / 116 = 1
    16'b10100010_01110101 : OUT <= 1;  //162 / 117 = 1
    16'b10100010_01110110 : OUT <= 1;  //162 / 118 = 1
    16'b10100010_01110111 : OUT <= 1;  //162 / 119 = 1
    16'b10100010_01111000 : OUT <= 1;  //162 / 120 = 1
    16'b10100010_01111001 : OUT <= 1;  //162 / 121 = 1
    16'b10100010_01111010 : OUT <= 1;  //162 / 122 = 1
    16'b10100010_01111011 : OUT <= 1;  //162 / 123 = 1
    16'b10100010_01111100 : OUT <= 1;  //162 / 124 = 1
    16'b10100010_01111101 : OUT <= 1;  //162 / 125 = 1
    16'b10100010_01111110 : OUT <= 1;  //162 / 126 = 1
    16'b10100010_01111111 : OUT <= 1;  //162 / 127 = 1
    16'b10100010_10000000 : OUT <= 1;  //162 / 128 = 1
    16'b10100010_10000001 : OUT <= 1;  //162 / 129 = 1
    16'b10100010_10000010 : OUT <= 1;  //162 / 130 = 1
    16'b10100010_10000011 : OUT <= 1;  //162 / 131 = 1
    16'b10100010_10000100 : OUT <= 1;  //162 / 132 = 1
    16'b10100010_10000101 : OUT <= 1;  //162 / 133 = 1
    16'b10100010_10000110 : OUT <= 1;  //162 / 134 = 1
    16'b10100010_10000111 : OUT <= 1;  //162 / 135 = 1
    16'b10100010_10001000 : OUT <= 1;  //162 / 136 = 1
    16'b10100010_10001001 : OUT <= 1;  //162 / 137 = 1
    16'b10100010_10001010 : OUT <= 1;  //162 / 138 = 1
    16'b10100010_10001011 : OUT <= 1;  //162 / 139 = 1
    16'b10100010_10001100 : OUT <= 1;  //162 / 140 = 1
    16'b10100010_10001101 : OUT <= 1;  //162 / 141 = 1
    16'b10100010_10001110 : OUT <= 1;  //162 / 142 = 1
    16'b10100010_10001111 : OUT <= 1;  //162 / 143 = 1
    16'b10100010_10010000 : OUT <= 1;  //162 / 144 = 1
    16'b10100010_10010001 : OUT <= 1;  //162 / 145 = 1
    16'b10100010_10010010 : OUT <= 1;  //162 / 146 = 1
    16'b10100010_10010011 : OUT <= 1;  //162 / 147 = 1
    16'b10100010_10010100 : OUT <= 1;  //162 / 148 = 1
    16'b10100010_10010101 : OUT <= 1;  //162 / 149 = 1
    16'b10100010_10010110 : OUT <= 1;  //162 / 150 = 1
    16'b10100010_10010111 : OUT <= 1;  //162 / 151 = 1
    16'b10100010_10011000 : OUT <= 1;  //162 / 152 = 1
    16'b10100010_10011001 : OUT <= 1;  //162 / 153 = 1
    16'b10100010_10011010 : OUT <= 1;  //162 / 154 = 1
    16'b10100010_10011011 : OUT <= 1;  //162 / 155 = 1
    16'b10100010_10011100 : OUT <= 1;  //162 / 156 = 1
    16'b10100010_10011101 : OUT <= 1;  //162 / 157 = 1
    16'b10100010_10011110 : OUT <= 1;  //162 / 158 = 1
    16'b10100010_10011111 : OUT <= 1;  //162 / 159 = 1
    16'b10100010_10100000 : OUT <= 1;  //162 / 160 = 1
    16'b10100010_10100001 : OUT <= 1;  //162 / 161 = 1
    16'b10100010_10100010 : OUT <= 1;  //162 / 162 = 1
    16'b10100010_10100011 : OUT <= 0;  //162 / 163 = 0
    16'b10100010_10100100 : OUT <= 0;  //162 / 164 = 0
    16'b10100010_10100101 : OUT <= 0;  //162 / 165 = 0
    16'b10100010_10100110 : OUT <= 0;  //162 / 166 = 0
    16'b10100010_10100111 : OUT <= 0;  //162 / 167 = 0
    16'b10100010_10101000 : OUT <= 0;  //162 / 168 = 0
    16'b10100010_10101001 : OUT <= 0;  //162 / 169 = 0
    16'b10100010_10101010 : OUT <= 0;  //162 / 170 = 0
    16'b10100010_10101011 : OUT <= 0;  //162 / 171 = 0
    16'b10100010_10101100 : OUT <= 0;  //162 / 172 = 0
    16'b10100010_10101101 : OUT <= 0;  //162 / 173 = 0
    16'b10100010_10101110 : OUT <= 0;  //162 / 174 = 0
    16'b10100010_10101111 : OUT <= 0;  //162 / 175 = 0
    16'b10100010_10110000 : OUT <= 0;  //162 / 176 = 0
    16'b10100010_10110001 : OUT <= 0;  //162 / 177 = 0
    16'b10100010_10110010 : OUT <= 0;  //162 / 178 = 0
    16'b10100010_10110011 : OUT <= 0;  //162 / 179 = 0
    16'b10100010_10110100 : OUT <= 0;  //162 / 180 = 0
    16'b10100010_10110101 : OUT <= 0;  //162 / 181 = 0
    16'b10100010_10110110 : OUT <= 0;  //162 / 182 = 0
    16'b10100010_10110111 : OUT <= 0;  //162 / 183 = 0
    16'b10100010_10111000 : OUT <= 0;  //162 / 184 = 0
    16'b10100010_10111001 : OUT <= 0;  //162 / 185 = 0
    16'b10100010_10111010 : OUT <= 0;  //162 / 186 = 0
    16'b10100010_10111011 : OUT <= 0;  //162 / 187 = 0
    16'b10100010_10111100 : OUT <= 0;  //162 / 188 = 0
    16'b10100010_10111101 : OUT <= 0;  //162 / 189 = 0
    16'b10100010_10111110 : OUT <= 0;  //162 / 190 = 0
    16'b10100010_10111111 : OUT <= 0;  //162 / 191 = 0
    16'b10100010_11000000 : OUT <= 0;  //162 / 192 = 0
    16'b10100010_11000001 : OUT <= 0;  //162 / 193 = 0
    16'b10100010_11000010 : OUT <= 0;  //162 / 194 = 0
    16'b10100010_11000011 : OUT <= 0;  //162 / 195 = 0
    16'b10100010_11000100 : OUT <= 0;  //162 / 196 = 0
    16'b10100010_11000101 : OUT <= 0;  //162 / 197 = 0
    16'b10100010_11000110 : OUT <= 0;  //162 / 198 = 0
    16'b10100010_11000111 : OUT <= 0;  //162 / 199 = 0
    16'b10100010_11001000 : OUT <= 0;  //162 / 200 = 0
    16'b10100010_11001001 : OUT <= 0;  //162 / 201 = 0
    16'b10100010_11001010 : OUT <= 0;  //162 / 202 = 0
    16'b10100010_11001011 : OUT <= 0;  //162 / 203 = 0
    16'b10100010_11001100 : OUT <= 0;  //162 / 204 = 0
    16'b10100010_11001101 : OUT <= 0;  //162 / 205 = 0
    16'b10100010_11001110 : OUT <= 0;  //162 / 206 = 0
    16'b10100010_11001111 : OUT <= 0;  //162 / 207 = 0
    16'b10100010_11010000 : OUT <= 0;  //162 / 208 = 0
    16'b10100010_11010001 : OUT <= 0;  //162 / 209 = 0
    16'b10100010_11010010 : OUT <= 0;  //162 / 210 = 0
    16'b10100010_11010011 : OUT <= 0;  //162 / 211 = 0
    16'b10100010_11010100 : OUT <= 0;  //162 / 212 = 0
    16'b10100010_11010101 : OUT <= 0;  //162 / 213 = 0
    16'b10100010_11010110 : OUT <= 0;  //162 / 214 = 0
    16'b10100010_11010111 : OUT <= 0;  //162 / 215 = 0
    16'b10100010_11011000 : OUT <= 0;  //162 / 216 = 0
    16'b10100010_11011001 : OUT <= 0;  //162 / 217 = 0
    16'b10100010_11011010 : OUT <= 0;  //162 / 218 = 0
    16'b10100010_11011011 : OUT <= 0;  //162 / 219 = 0
    16'b10100010_11011100 : OUT <= 0;  //162 / 220 = 0
    16'b10100010_11011101 : OUT <= 0;  //162 / 221 = 0
    16'b10100010_11011110 : OUT <= 0;  //162 / 222 = 0
    16'b10100010_11011111 : OUT <= 0;  //162 / 223 = 0
    16'b10100010_11100000 : OUT <= 0;  //162 / 224 = 0
    16'b10100010_11100001 : OUT <= 0;  //162 / 225 = 0
    16'b10100010_11100010 : OUT <= 0;  //162 / 226 = 0
    16'b10100010_11100011 : OUT <= 0;  //162 / 227 = 0
    16'b10100010_11100100 : OUT <= 0;  //162 / 228 = 0
    16'b10100010_11100101 : OUT <= 0;  //162 / 229 = 0
    16'b10100010_11100110 : OUT <= 0;  //162 / 230 = 0
    16'b10100010_11100111 : OUT <= 0;  //162 / 231 = 0
    16'b10100010_11101000 : OUT <= 0;  //162 / 232 = 0
    16'b10100010_11101001 : OUT <= 0;  //162 / 233 = 0
    16'b10100010_11101010 : OUT <= 0;  //162 / 234 = 0
    16'b10100010_11101011 : OUT <= 0;  //162 / 235 = 0
    16'b10100010_11101100 : OUT <= 0;  //162 / 236 = 0
    16'b10100010_11101101 : OUT <= 0;  //162 / 237 = 0
    16'b10100010_11101110 : OUT <= 0;  //162 / 238 = 0
    16'b10100010_11101111 : OUT <= 0;  //162 / 239 = 0
    16'b10100010_11110000 : OUT <= 0;  //162 / 240 = 0
    16'b10100010_11110001 : OUT <= 0;  //162 / 241 = 0
    16'b10100010_11110010 : OUT <= 0;  //162 / 242 = 0
    16'b10100010_11110011 : OUT <= 0;  //162 / 243 = 0
    16'b10100010_11110100 : OUT <= 0;  //162 / 244 = 0
    16'b10100010_11110101 : OUT <= 0;  //162 / 245 = 0
    16'b10100010_11110110 : OUT <= 0;  //162 / 246 = 0
    16'b10100010_11110111 : OUT <= 0;  //162 / 247 = 0
    16'b10100010_11111000 : OUT <= 0;  //162 / 248 = 0
    16'b10100010_11111001 : OUT <= 0;  //162 / 249 = 0
    16'b10100010_11111010 : OUT <= 0;  //162 / 250 = 0
    16'b10100010_11111011 : OUT <= 0;  //162 / 251 = 0
    16'b10100010_11111100 : OUT <= 0;  //162 / 252 = 0
    16'b10100010_11111101 : OUT <= 0;  //162 / 253 = 0
    16'b10100010_11111110 : OUT <= 0;  //162 / 254 = 0
    16'b10100010_11111111 : OUT <= 0;  //162 / 255 = 0
    16'b10100011_00000000 : OUT <= 0;  //163 / 0 = 0
    16'b10100011_00000001 : OUT <= 163;  //163 / 1 = 163
    16'b10100011_00000010 : OUT <= 81;  //163 / 2 = 81
    16'b10100011_00000011 : OUT <= 54;  //163 / 3 = 54
    16'b10100011_00000100 : OUT <= 40;  //163 / 4 = 40
    16'b10100011_00000101 : OUT <= 32;  //163 / 5 = 32
    16'b10100011_00000110 : OUT <= 27;  //163 / 6 = 27
    16'b10100011_00000111 : OUT <= 23;  //163 / 7 = 23
    16'b10100011_00001000 : OUT <= 20;  //163 / 8 = 20
    16'b10100011_00001001 : OUT <= 18;  //163 / 9 = 18
    16'b10100011_00001010 : OUT <= 16;  //163 / 10 = 16
    16'b10100011_00001011 : OUT <= 14;  //163 / 11 = 14
    16'b10100011_00001100 : OUT <= 13;  //163 / 12 = 13
    16'b10100011_00001101 : OUT <= 12;  //163 / 13 = 12
    16'b10100011_00001110 : OUT <= 11;  //163 / 14 = 11
    16'b10100011_00001111 : OUT <= 10;  //163 / 15 = 10
    16'b10100011_00010000 : OUT <= 10;  //163 / 16 = 10
    16'b10100011_00010001 : OUT <= 9;  //163 / 17 = 9
    16'b10100011_00010010 : OUT <= 9;  //163 / 18 = 9
    16'b10100011_00010011 : OUT <= 8;  //163 / 19 = 8
    16'b10100011_00010100 : OUT <= 8;  //163 / 20 = 8
    16'b10100011_00010101 : OUT <= 7;  //163 / 21 = 7
    16'b10100011_00010110 : OUT <= 7;  //163 / 22 = 7
    16'b10100011_00010111 : OUT <= 7;  //163 / 23 = 7
    16'b10100011_00011000 : OUT <= 6;  //163 / 24 = 6
    16'b10100011_00011001 : OUT <= 6;  //163 / 25 = 6
    16'b10100011_00011010 : OUT <= 6;  //163 / 26 = 6
    16'b10100011_00011011 : OUT <= 6;  //163 / 27 = 6
    16'b10100011_00011100 : OUT <= 5;  //163 / 28 = 5
    16'b10100011_00011101 : OUT <= 5;  //163 / 29 = 5
    16'b10100011_00011110 : OUT <= 5;  //163 / 30 = 5
    16'b10100011_00011111 : OUT <= 5;  //163 / 31 = 5
    16'b10100011_00100000 : OUT <= 5;  //163 / 32 = 5
    16'b10100011_00100001 : OUT <= 4;  //163 / 33 = 4
    16'b10100011_00100010 : OUT <= 4;  //163 / 34 = 4
    16'b10100011_00100011 : OUT <= 4;  //163 / 35 = 4
    16'b10100011_00100100 : OUT <= 4;  //163 / 36 = 4
    16'b10100011_00100101 : OUT <= 4;  //163 / 37 = 4
    16'b10100011_00100110 : OUT <= 4;  //163 / 38 = 4
    16'b10100011_00100111 : OUT <= 4;  //163 / 39 = 4
    16'b10100011_00101000 : OUT <= 4;  //163 / 40 = 4
    16'b10100011_00101001 : OUT <= 3;  //163 / 41 = 3
    16'b10100011_00101010 : OUT <= 3;  //163 / 42 = 3
    16'b10100011_00101011 : OUT <= 3;  //163 / 43 = 3
    16'b10100011_00101100 : OUT <= 3;  //163 / 44 = 3
    16'b10100011_00101101 : OUT <= 3;  //163 / 45 = 3
    16'b10100011_00101110 : OUT <= 3;  //163 / 46 = 3
    16'b10100011_00101111 : OUT <= 3;  //163 / 47 = 3
    16'b10100011_00110000 : OUT <= 3;  //163 / 48 = 3
    16'b10100011_00110001 : OUT <= 3;  //163 / 49 = 3
    16'b10100011_00110010 : OUT <= 3;  //163 / 50 = 3
    16'b10100011_00110011 : OUT <= 3;  //163 / 51 = 3
    16'b10100011_00110100 : OUT <= 3;  //163 / 52 = 3
    16'b10100011_00110101 : OUT <= 3;  //163 / 53 = 3
    16'b10100011_00110110 : OUT <= 3;  //163 / 54 = 3
    16'b10100011_00110111 : OUT <= 2;  //163 / 55 = 2
    16'b10100011_00111000 : OUT <= 2;  //163 / 56 = 2
    16'b10100011_00111001 : OUT <= 2;  //163 / 57 = 2
    16'b10100011_00111010 : OUT <= 2;  //163 / 58 = 2
    16'b10100011_00111011 : OUT <= 2;  //163 / 59 = 2
    16'b10100011_00111100 : OUT <= 2;  //163 / 60 = 2
    16'b10100011_00111101 : OUT <= 2;  //163 / 61 = 2
    16'b10100011_00111110 : OUT <= 2;  //163 / 62 = 2
    16'b10100011_00111111 : OUT <= 2;  //163 / 63 = 2
    16'b10100011_01000000 : OUT <= 2;  //163 / 64 = 2
    16'b10100011_01000001 : OUT <= 2;  //163 / 65 = 2
    16'b10100011_01000010 : OUT <= 2;  //163 / 66 = 2
    16'b10100011_01000011 : OUT <= 2;  //163 / 67 = 2
    16'b10100011_01000100 : OUT <= 2;  //163 / 68 = 2
    16'b10100011_01000101 : OUT <= 2;  //163 / 69 = 2
    16'b10100011_01000110 : OUT <= 2;  //163 / 70 = 2
    16'b10100011_01000111 : OUT <= 2;  //163 / 71 = 2
    16'b10100011_01001000 : OUT <= 2;  //163 / 72 = 2
    16'b10100011_01001001 : OUT <= 2;  //163 / 73 = 2
    16'b10100011_01001010 : OUT <= 2;  //163 / 74 = 2
    16'b10100011_01001011 : OUT <= 2;  //163 / 75 = 2
    16'b10100011_01001100 : OUT <= 2;  //163 / 76 = 2
    16'b10100011_01001101 : OUT <= 2;  //163 / 77 = 2
    16'b10100011_01001110 : OUT <= 2;  //163 / 78 = 2
    16'b10100011_01001111 : OUT <= 2;  //163 / 79 = 2
    16'b10100011_01010000 : OUT <= 2;  //163 / 80 = 2
    16'b10100011_01010001 : OUT <= 2;  //163 / 81 = 2
    16'b10100011_01010010 : OUT <= 1;  //163 / 82 = 1
    16'b10100011_01010011 : OUT <= 1;  //163 / 83 = 1
    16'b10100011_01010100 : OUT <= 1;  //163 / 84 = 1
    16'b10100011_01010101 : OUT <= 1;  //163 / 85 = 1
    16'b10100011_01010110 : OUT <= 1;  //163 / 86 = 1
    16'b10100011_01010111 : OUT <= 1;  //163 / 87 = 1
    16'b10100011_01011000 : OUT <= 1;  //163 / 88 = 1
    16'b10100011_01011001 : OUT <= 1;  //163 / 89 = 1
    16'b10100011_01011010 : OUT <= 1;  //163 / 90 = 1
    16'b10100011_01011011 : OUT <= 1;  //163 / 91 = 1
    16'b10100011_01011100 : OUT <= 1;  //163 / 92 = 1
    16'b10100011_01011101 : OUT <= 1;  //163 / 93 = 1
    16'b10100011_01011110 : OUT <= 1;  //163 / 94 = 1
    16'b10100011_01011111 : OUT <= 1;  //163 / 95 = 1
    16'b10100011_01100000 : OUT <= 1;  //163 / 96 = 1
    16'b10100011_01100001 : OUT <= 1;  //163 / 97 = 1
    16'b10100011_01100010 : OUT <= 1;  //163 / 98 = 1
    16'b10100011_01100011 : OUT <= 1;  //163 / 99 = 1
    16'b10100011_01100100 : OUT <= 1;  //163 / 100 = 1
    16'b10100011_01100101 : OUT <= 1;  //163 / 101 = 1
    16'b10100011_01100110 : OUT <= 1;  //163 / 102 = 1
    16'b10100011_01100111 : OUT <= 1;  //163 / 103 = 1
    16'b10100011_01101000 : OUT <= 1;  //163 / 104 = 1
    16'b10100011_01101001 : OUT <= 1;  //163 / 105 = 1
    16'b10100011_01101010 : OUT <= 1;  //163 / 106 = 1
    16'b10100011_01101011 : OUT <= 1;  //163 / 107 = 1
    16'b10100011_01101100 : OUT <= 1;  //163 / 108 = 1
    16'b10100011_01101101 : OUT <= 1;  //163 / 109 = 1
    16'b10100011_01101110 : OUT <= 1;  //163 / 110 = 1
    16'b10100011_01101111 : OUT <= 1;  //163 / 111 = 1
    16'b10100011_01110000 : OUT <= 1;  //163 / 112 = 1
    16'b10100011_01110001 : OUT <= 1;  //163 / 113 = 1
    16'b10100011_01110010 : OUT <= 1;  //163 / 114 = 1
    16'b10100011_01110011 : OUT <= 1;  //163 / 115 = 1
    16'b10100011_01110100 : OUT <= 1;  //163 / 116 = 1
    16'b10100011_01110101 : OUT <= 1;  //163 / 117 = 1
    16'b10100011_01110110 : OUT <= 1;  //163 / 118 = 1
    16'b10100011_01110111 : OUT <= 1;  //163 / 119 = 1
    16'b10100011_01111000 : OUT <= 1;  //163 / 120 = 1
    16'b10100011_01111001 : OUT <= 1;  //163 / 121 = 1
    16'b10100011_01111010 : OUT <= 1;  //163 / 122 = 1
    16'b10100011_01111011 : OUT <= 1;  //163 / 123 = 1
    16'b10100011_01111100 : OUT <= 1;  //163 / 124 = 1
    16'b10100011_01111101 : OUT <= 1;  //163 / 125 = 1
    16'b10100011_01111110 : OUT <= 1;  //163 / 126 = 1
    16'b10100011_01111111 : OUT <= 1;  //163 / 127 = 1
    16'b10100011_10000000 : OUT <= 1;  //163 / 128 = 1
    16'b10100011_10000001 : OUT <= 1;  //163 / 129 = 1
    16'b10100011_10000010 : OUT <= 1;  //163 / 130 = 1
    16'b10100011_10000011 : OUT <= 1;  //163 / 131 = 1
    16'b10100011_10000100 : OUT <= 1;  //163 / 132 = 1
    16'b10100011_10000101 : OUT <= 1;  //163 / 133 = 1
    16'b10100011_10000110 : OUT <= 1;  //163 / 134 = 1
    16'b10100011_10000111 : OUT <= 1;  //163 / 135 = 1
    16'b10100011_10001000 : OUT <= 1;  //163 / 136 = 1
    16'b10100011_10001001 : OUT <= 1;  //163 / 137 = 1
    16'b10100011_10001010 : OUT <= 1;  //163 / 138 = 1
    16'b10100011_10001011 : OUT <= 1;  //163 / 139 = 1
    16'b10100011_10001100 : OUT <= 1;  //163 / 140 = 1
    16'b10100011_10001101 : OUT <= 1;  //163 / 141 = 1
    16'b10100011_10001110 : OUT <= 1;  //163 / 142 = 1
    16'b10100011_10001111 : OUT <= 1;  //163 / 143 = 1
    16'b10100011_10010000 : OUT <= 1;  //163 / 144 = 1
    16'b10100011_10010001 : OUT <= 1;  //163 / 145 = 1
    16'b10100011_10010010 : OUT <= 1;  //163 / 146 = 1
    16'b10100011_10010011 : OUT <= 1;  //163 / 147 = 1
    16'b10100011_10010100 : OUT <= 1;  //163 / 148 = 1
    16'b10100011_10010101 : OUT <= 1;  //163 / 149 = 1
    16'b10100011_10010110 : OUT <= 1;  //163 / 150 = 1
    16'b10100011_10010111 : OUT <= 1;  //163 / 151 = 1
    16'b10100011_10011000 : OUT <= 1;  //163 / 152 = 1
    16'b10100011_10011001 : OUT <= 1;  //163 / 153 = 1
    16'b10100011_10011010 : OUT <= 1;  //163 / 154 = 1
    16'b10100011_10011011 : OUT <= 1;  //163 / 155 = 1
    16'b10100011_10011100 : OUT <= 1;  //163 / 156 = 1
    16'b10100011_10011101 : OUT <= 1;  //163 / 157 = 1
    16'b10100011_10011110 : OUT <= 1;  //163 / 158 = 1
    16'b10100011_10011111 : OUT <= 1;  //163 / 159 = 1
    16'b10100011_10100000 : OUT <= 1;  //163 / 160 = 1
    16'b10100011_10100001 : OUT <= 1;  //163 / 161 = 1
    16'b10100011_10100010 : OUT <= 1;  //163 / 162 = 1
    16'b10100011_10100011 : OUT <= 1;  //163 / 163 = 1
    16'b10100011_10100100 : OUT <= 0;  //163 / 164 = 0
    16'b10100011_10100101 : OUT <= 0;  //163 / 165 = 0
    16'b10100011_10100110 : OUT <= 0;  //163 / 166 = 0
    16'b10100011_10100111 : OUT <= 0;  //163 / 167 = 0
    16'b10100011_10101000 : OUT <= 0;  //163 / 168 = 0
    16'b10100011_10101001 : OUT <= 0;  //163 / 169 = 0
    16'b10100011_10101010 : OUT <= 0;  //163 / 170 = 0
    16'b10100011_10101011 : OUT <= 0;  //163 / 171 = 0
    16'b10100011_10101100 : OUT <= 0;  //163 / 172 = 0
    16'b10100011_10101101 : OUT <= 0;  //163 / 173 = 0
    16'b10100011_10101110 : OUT <= 0;  //163 / 174 = 0
    16'b10100011_10101111 : OUT <= 0;  //163 / 175 = 0
    16'b10100011_10110000 : OUT <= 0;  //163 / 176 = 0
    16'b10100011_10110001 : OUT <= 0;  //163 / 177 = 0
    16'b10100011_10110010 : OUT <= 0;  //163 / 178 = 0
    16'b10100011_10110011 : OUT <= 0;  //163 / 179 = 0
    16'b10100011_10110100 : OUT <= 0;  //163 / 180 = 0
    16'b10100011_10110101 : OUT <= 0;  //163 / 181 = 0
    16'b10100011_10110110 : OUT <= 0;  //163 / 182 = 0
    16'b10100011_10110111 : OUT <= 0;  //163 / 183 = 0
    16'b10100011_10111000 : OUT <= 0;  //163 / 184 = 0
    16'b10100011_10111001 : OUT <= 0;  //163 / 185 = 0
    16'b10100011_10111010 : OUT <= 0;  //163 / 186 = 0
    16'b10100011_10111011 : OUT <= 0;  //163 / 187 = 0
    16'b10100011_10111100 : OUT <= 0;  //163 / 188 = 0
    16'b10100011_10111101 : OUT <= 0;  //163 / 189 = 0
    16'b10100011_10111110 : OUT <= 0;  //163 / 190 = 0
    16'b10100011_10111111 : OUT <= 0;  //163 / 191 = 0
    16'b10100011_11000000 : OUT <= 0;  //163 / 192 = 0
    16'b10100011_11000001 : OUT <= 0;  //163 / 193 = 0
    16'b10100011_11000010 : OUT <= 0;  //163 / 194 = 0
    16'b10100011_11000011 : OUT <= 0;  //163 / 195 = 0
    16'b10100011_11000100 : OUT <= 0;  //163 / 196 = 0
    16'b10100011_11000101 : OUT <= 0;  //163 / 197 = 0
    16'b10100011_11000110 : OUT <= 0;  //163 / 198 = 0
    16'b10100011_11000111 : OUT <= 0;  //163 / 199 = 0
    16'b10100011_11001000 : OUT <= 0;  //163 / 200 = 0
    16'b10100011_11001001 : OUT <= 0;  //163 / 201 = 0
    16'b10100011_11001010 : OUT <= 0;  //163 / 202 = 0
    16'b10100011_11001011 : OUT <= 0;  //163 / 203 = 0
    16'b10100011_11001100 : OUT <= 0;  //163 / 204 = 0
    16'b10100011_11001101 : OUT <= 0;  //163 / 205 = 0
    16'b10100011_11001110 : OUT <= 0;  //163 / 206 = 0
    16'b10100011_11001111 : OUT <= 0;  //163 / 207 = 0
    16'b10100011_11010000 : OUT <= 0;  //163 / 208 = 0
    16'b10100011_11010001 : OUT <= 0;  //163 / 209 = 0
    16'b10100011_11010010 : OUT <= 0;  //163 / 210 = 0
    16'b10100011_11010011 : OUT <= 0;  //163 / 211 = 0
    16'b10100011_11010100 : OUT <= 0;  //163 / 212 = 0
    16'b10100011_11010101 : OUT <= 0;  //163 / 213 = 0
    16'b10100011_11010110 : OUT <= 0;  //163 / 214 = 0
    16'b10100011_11010111 : OUT <= 0;  //163 / 215 = 0
    16'b10100011_11011000 : OUT <= 0;  //163 / 216 = 0
    16'b10100011_11011001 : OUT <= 0;  //163 / 217 = 0
    16'b10100011_11011010 : OUT <= 0;  //163 / 218 = 0
    16'b10100011_11011011 : OUT <= 0;  //163 / 219 = 0
    16'b10100011_11011100 : OUT <= 0;  //163 / 220 = 0
    16'b10100011_11011101 : OUT <= 0;  //163 / 221 = 0
    16'b10100011_11011110 : OUT <= 0;  //163 / 222 = 0
    16'b10100011_11011111 : OUT <= 0;  //163 / 223 = 0
    16'b10100011_11100000 : OUT <= 0;  //163 / 224 = 0
    16'b10100011_11100001 : OUT <= 0;  //163 / 225 = 0
    16'b10100011_11100010 : OUT <= 0;  //163 / 226 = 0
    16'b10100011_11100011 : OUT <= 0;  //163 / 227 = 0
    16'b10100011_11100100 : OUT <= 0;  //163 / 228 = 0
    16'b10100011_11100101 : OUT <= 0;  //163 / 229 = 0
    16'b10100011_11100110 : OUT <= 0;  //163 / 230 = 0
    16'b10100011_11100111 : OUT <= 0;  //163 / 231 = 0
    16'b10100011_11101000 : OUT <= 0;  //163 / 232 = 0
    16'b10100011_11101001 : OUT <= 0;  //163 / 233 = 0
    16'b10100011_11101010 : OUT <= 0;  //163 / 234 = 0
    16'b10100011_11101011 : OUT <= 0;  //163 / 235 = 0
    16'b10100011_11101100 : OUT <= 0;  //163 / 236 = 0
    16'b10100011_11101101 : OUT <= 0;  //163 / 237 = 0
    16'b10100011_11101110 : OUT <= 0;  //163 / 238 = 0
    16'b10100011_11101111 : OUT <= 0;  //163 / 239 = 0
    16'b10100011_11110000 : OUT <= 0;  //163 / 240 = 0
    16'b10100011_11110001 : OUT <= 0;  //163 / 241 = 0
    16'b10100011_11110010 : OUT <= 0;  //163 / 242 = 0
    16'b10100011_11110011 : OUT <= 0;  //163 / 243 = 0
    16'b10100011_11110100 : OUT <= 0;  //163 / 244 = 0
    16'b10100011_11110101 : OUT <= 0;  //163 / 245 = 0
    16'b10100011_11110110 : OUT <= 0;  //163 / 246 = 0
    16'b10100011_11110111 : OUT <= 0;  //163 / 247 = 0
    16'b10100011_11111000 : OUT <= 0;  //163 / 248 = 0
    16'b10100011_11111001 : OUT <= 0;  //163 / 249 = 0
    16'b10100011_11111010 : OUT <= 0;  //163 / 250 = 0
    16'b10100011_11111011 : OUT <= 0;  //163 / 251 = 0
    16'b10100011_11111100 : OUT <= 0;  //163 / 252 = 0
    16'b10100011_11111101 : OUT <= 0;  //163 / 253 = 0
    16'b10100011_11111110 : OUT <= 0;  //163 / 254 = 0
    16'b10100011_11111111 : OUT <= 0;  //163 / 255 = 0
    16'b10100100_00000000 : OUT <= 0;  //164 / 0 = 0
    16'b10100100_00000001 : OUT <= 164;  //164 / 1 = 164
    16'b10100100_00000010 : OUT <= 82;  //164 / 2 = 82
    16'b10100100_00000011 : OUT <= 54;  //164 / 3 = 54
    16'b10100100_00000100 : OUT <= 41;  //164 / 4 = 41
    16'b10100100_00000101 : OUT <= 32;  //164 / 5 = 32
    16'b10100100_00000110 : OUT <= 27;  //164 / 6 = 27
    16'b10100100_00000111 : OUT <= 23;  //164 / 7 = 23
    16'b10100100_00001000 : OUT <= 20;  //164 / 8 = 20
    16'b10100100_00001001 : OUT <= 18;  //164 / 9 = 18
    16'b10100100_00001010 : OUT <= 16;  //164 / 10 = 16
    16'b10100100_00001011 : OUT <= 14;  //164 / 11 = 14
    16'b10100100_00001100 : OUT <= 13;  //164 / 12 = 13
    16'b10100100_00001101 : OUT <= 12;  //164 / 13 = 12
    16'b10100100_00001110 : OUT <= 11;  //164 / 14 = 11
    16'b10100100_00001111 : OUT <= 10;  //164 / 15 = 10
    16'b10100100_00010000 : OUT <= 10;  //164 / 16 = 10
    16'b10100100_00010001 : OUT <= 9;  //164 / 17 = 9
    16'b10100100_00010010 : OUT <= 9;  //164 / 18 = 9
    16'b10100100_00010011 : OUT <= 8;  //164 / 19 = 8
    16'b10100100_00010100 : OUT <= 8;  //164 / 20 = 8
    16'b10100100_00010101 : OUT <= 7;  //164 / 21 = 7
    16'b10100100_00010110 : OUT <= 7;  //164 / 22 = 7
    16'b10100100_00010111 : OUT <= 7;  //164 / 23 = 7
    16'b10100100_00011000 : OUT <= 6;  //164 / 24 = 6
    16'b10100100_00011001 : OUT <= 6;  //164 / 25 = 6
    16'b10100100_00011010 : OUT <= 6;  //164 / 26 = 6
    16'b10100100_00011011 : OUT <= 6;  //164 / 27 = 6
    16'b10100100_00011100 : OUT <= 5;  //164 / 28 = 5
    16'b10100100_00011101 : OUT <= 5;  //164 / 29 = 5
    16'b10100100_00011110 : OUT <= 5;  //164 / 30 = 5
    16'b10100100_00011111 : OUT <= 5;  //164 / 31 = 5
    16'b10100100_00100000 : OUT <= 5;  //164 / 32 = 5
    16'b10100100_00100001 : OUT <= 4;  //164 / 33 = 4
    16'b10100100_00100010 : OUT <= 4;  //164 / 34 = 4
    16'b10100100_00100011 : OUT <= 4;  //164 / 35 = 4
    16'b10100100_00100100 : OUT <= 4;  //164 / 36 = 4
    16'b10100100_00100101 : OUT <= 4;  //164 / 37 = 4
    16'b10100100_00100110 : OUT <= 4;  //164 / 38 = 4
    16'b10100100_00100111 : OUT <= 4;  //164 / 39 = 4
    16'b10100100_00101000 : OUT <= 4;  //164 / 40 = 4
    16'b10100100_00101001 : OUT <= 4;  //164 / 41 = 4
    16'b10100100_00101010 : OUT <= 3;  //164 / 42 = 3
    16'b10100100_00101011 : OUT <= 3;  //164 / 43 = 3
    16'b10100100_00101100 : OUT <= 3;  //164 / 44 = 3
    16'b10100100_00101101 : OUT <= 3;  //164 / 45 = 3
    16'b10100100_00101110 : OUT <= 3;  //164 / 46 = 3
    16'b10100100_00101111 : OUT <= 3;  //164 / 47 = 3
    16'b10100100_00110000 : OUT <= 3;  //164 / 48 = 3
    16'b10100100_00110001 : OUT <= 3;  //164 / 49 = 3
    16'b10100100_00110010 : OUT <= 3;  //164 / 50 = 3
    16'b10100100_00110011 : OUT <= 3;  //164 / 51 = 3
    16'b10100100_00110100 : OUT <= 3;  //164 / 52 = 3
    16'b10100100_00110101 : OUT <= 3;  //164 / 53 = 3
    16'b10100100_00110110 : OUT <= 3;  //164 / 54 = 3
    16'b10100100_00110111 : OUT <= 2;  //164 / 55 = 2
    16'b10100100_00111000 : OUT <= 2;  //164 / 56 = 2
    16'b10100100_00111001 : OUT <= 2;  //164 / 57 = 2
    16'b10100100_00111010 : OUT <= 2;  //164 / 58 = 2
    16'b10100100_00111011 : OUT <= 2;  //164 / 59 = 2
    16'b10100100_00111100 : OUT <= 2;  //164 / 60 = 2
    16'b10100100_00111101 : OUT <= 2;  //164 / 61 = 2
    16'b10100100_00111110 : OUT <= 2;  //164 / 62 = 2
    16'b10100100_00111111 : OUT <= 2;  //164 / 63 = 2
    16'b10100100_01000000 : OUT <= 2;  //164 / 64 = 2
    16'b10100100_01000001 : OUT <= 2;  //164 / 65 = 2
    16'b10100100_01000010 : OUT <= 2;  //164 / 66 = 2
    16'b10100100_01000011 : OUT <= 2;  //164 / 67 = 2
    16'b10100100_01000100 : OUT <= 2;  //164 / 68 = 2
    16'b10100100_01000101 : OUT <= 2;  //164 / 69 = 2
    16'b10100100_01000110 : OUT <= 2;  //164 / 70 = 2
    16'b10100100_01000111 : OUT <= 2;  //164 / 71 = 2
    16'b10100100_01001000 : OUT <= 2;  //164 / 72 = 2
    16'b10100100_01001001 : OUT <= 2;  //164 / 73 = 2
    16'b10100100_01001010 : OUT <= 2;  //164 / 74 = 2
    16'b10100100_01001011 : OUT <= 2;  //164 / 75 = 2
    16'b10100100_01001100 : OUT <= 2;  //164 / 76 = 2
    16'b10100100_01001101 : OUT <= 2;  //164 / 77 = 2
    16'b10100100_01001110 : OUT <= 2;  //164 / 78 = 2
    16'b10100100_01001111 : OUT <= 2;  //164 / 79 = 2
    16'b10100100_01010000 : OUT <= 2;  //164 / 80 = 2
    16'b10100100_01010001 : OUT <= 2;  //164 / 81 = 2
    16'b10100100_01010010 : OUT <= 2;  //164 / 82 = 2
    16'b10100100_01010011 : OUT <= 1;  //164 / 83 = 1
    16'b10100100_01010100 : OUT <= 1;  //164 / 84 = 1
    16'b10100100_01010101 : OUT <= 1;  //164 / 85 = 1
    16'b10100100_01010110 : OUT <= 1;  //164 / 86 = 1
    16'b10100100_01010111 : OUT <= 1;  //164 / 87 = 1
    16'b10100100_01011000 : OUT <= 1;  //164 / 88 = 1
    16'b10100100_01011001 : OUT <= 1;  //164 / 89 = 1
    16'b10100100_01011010 : OUT <= 1;  //164 / 90 = 1
    16'b10100100_01011011 : OUT <= 1;  //164 / 91 = 1
    16'b10100100_01011100 : OUT <= 1;  //164 / 92 = 1
    16'b10100100_01011101 : OUT <= 1;  //164 / 93 = 1
    16'b10100100_01011110 : OUT <= 1;  //164 / 94 = 1
    16'b10100100_01011111 : OUT <= 1;  //164 / 95 = 1
    16'b10100100_01100000 : OUT <= 1;  //164 / 96 = 1
    16'b10100100_01100001 : OUT <= 1;  //164 / 97 = 1
    16'b10100100_01100010 : OUT <= 1;  //164 / 98 = 1
    16'b10100100_01100011 : OUT <= 1;  //164 / 99 = 1
    16'b10100100_01100100 : OUT <= 1;  //164 / 100 = 1
    16'b10100100_01100101 : OUT <= 1;  //164 / 101 = 1
    16'b10100100_01100110 : OUT <= 1;  //164 / 102 = 1
    16'b10100100_01100111 : OUT <= 1;  //164 / 103 = 1
    16'b10100100_01101000 : OUT <= 1;  //164 / 104 = 1
    16'b10100100_01101001 : OUT <= 1;  //164 / 105 = 1
    16'b10100100_01101010 : OUT <= 1;  //164 / 106 = 1
    16'b10100100_01101011 : OUT <= 1;  //164 / 107 = 1
    16'b10100100_01101100 : OUT <= 1;  //164 / 108 = 1
    16'b10100100_01101101 : OUT <= 1;  //164 / 109 = 1
    16'b10100100_01101110 : OUT <= 1;  //164 / 110 = 1
    16'b10100100_01101111 : OUT <= 1;  //164 / 111 = 1
    16'b10100100_01110000 : OUT <= 1;  //164 / 112 = 1
    16'b10100100_01110001 : OUT <= 1;  //164 / 113 = 1
    16'b10100100_01110010 : OUT <= 1;  //164 / 114 = 1
    16'b10100100_01110011 : OUT <= 1;  //164 / 115 = 1
    16'b10100100_01110100 : OUT <= 1;  //164 / 116 = 1
    16'b10100100_01110101 : OUT <= 1;  //164 / 117 = 1
    16'b10100100_01110110 : OUT <= 1;  //164 / 118 = 1
    16'b10100100_01110111 : OUT <= 1;  //164 / 119 = 1
    16'b10100100_01111000 : OUT <= 1;  //164 / 120 = 1
    16'b10100100_01111001 : OUT <= 1;  //164 / 121 = 1
    16'b10100100_01111010 : OUT <= 1;  //164 / 122 = 1
    16'b10100100_01111011 : OUT <= 1;  //164 / 123 = 1
    16'b10100100_01111100 : OUT <= 1;  //164 / 124 = 1
    16'b10100100_01111101 : OUT <= 1;  //164 / 125 = 1
    16'b10100100_01111110 : OUT <= 1;  //164 / 126 = 1
    16'b10100100_01111111 : OUT <= 1;  //164 / 127 = 1
    16'b10100100_10000000 : OUT <= 1;  //164 / 128 = 1
    16'b10100100_10000001 : OUT <= 1;  //164 / 129 = 1
    16'b10100100_10000010 : OUT <= 1;  //164 / 130 = 1
    16'b10100100_10000011 : OUT <= 1;  //164 / 131 = 1
    16'b10100100_10000100 : OUT <= 1;  //164 / 132 = 1
    16'b10100100_10000101 : OUT <= 1;  //164 / 133 = 1
    16'b10100100_10000110 : OUT <= 1;  //164 / 134 = 1
    16'b10100100_10000111 : OUT <= 1;  //164 / 135 = 1
    16'b10100100_10001000 : OUT <= 1;  //164 / 136 = 1
    16'b10100100_10001001 : OUT <= 1;  //164 / 137 = 1
    16'b10100100_10001010 : OUT <= 1;  //164 / 138 = 1
    16'b10100100_10001011 : OUT <= 1;  //164 / 139 = 1
    16'b10100100_10001100 : OUT <= 1;  //164 / 140 = 1
    16'b10100100_10001101 : OUT <= 1;  //164 / 141 = 1
    16'b10100100_10001110 : OUT <= 1;  //164 / 142 = 1
    16'b10100100_10001111 : OUT <= 1;  //164 / 143 = 1
    16'b10100100_10010000 : OUT <= 1;  //164 / 144 = 1
    16'b10100100_10010001 : OUT <= 1;  //164 / 145 = 1
    16'b10100100_10010010 : OUT <= 1;  //164 / 146 = 1
    16'b10100100_10010011 : OUT <= 1;  //164 / 147 = 1
    16'b10100100_10010100 : OUT <= 1;  //164 / 148 = 1
    16'b10100100_10010101 : OUT <= 1;  //164 / 149 = 1
    16'b10100100_10010110 : OUT <= 1;  //164 / 150 = 1
    16'b10100100_10010111 : OUT <= 1;  //164 / 151 = 1
    16'b10100100_10011000 : OUT <= 1;  //164 / 152 = 1
    16'b10100100_10011001 : OUT <= 1;  //164 / 153 = 1
    16'b10100100_10011010 : OUT <= 1;  //164 / 154 = 1
    16'b10100100_10011011 : OUT <= 1;  //164 / 155 = 1
    16'b10100100_10011100 : OUT <= 1;  //164 / 156 = 1
    16'b10100100_10011101 : OUT <= 1;  //164 / 157 = 1
    16'b10100100_10011110 : OUT <= 1;  //164 / 158 = 1
    16'b10100100_10011111 : OUT <= 1;  //164 / 159 = 1
    16'b10100100_10100000 : OUT <= 1;  //164 / 160 = 1
    16'b10100100_10100001 : OUT <= 1;  //164 / 161 = 1
    16'b10100100_10100010 : OUT <= 1;  //164 / 162 = 1
    16'b10100100_10100011 : OUT <= 1;  //164 / 163 = 1
    16'b10100100_10100100 : OUT <= 1;  //164 / 164 = 1
    16'b10100100_10100101 : OUT <= 0;  //164 / 165 = 0
    16'b10100100_10100110 : OUT <= 0;  //164 / 166 = 0
    16'b10100100_10100111 : OUT <= 0;  //164 / 167 = 0
    16'b10100100_10101000 : OUT <= 0;  //164 / 168 = 0
    16'b10100100_10101001 : OUT <= 0;  //164 / 169 = 0
    16'b10100100_10101010 : OUT <= 0;  //164 / 170 = 0
    16'b10100100_10101011 : OUT <= 0;  //164 / 171 = 0
    16'b10100100_10101100 : OUT <= 0;  //164 / 172 = 0
    16'b10100100_10101101 : OUT <= 0;  //164 / 173 = 0
    16'b10100100_10101110 : OUT <= 0;  //164 / 174 = 0
    16'b10100100_10101111 : OUT <= 0;  //164 / 175 = 0
    16'b10100100_10110000 : OUT <= 0;  //164 / 176 = 0
    16'b10100100_10110001 : OUT <= 0;  //164 / 177 = 0
    16'b10100100_10110010 : OUT <= 0;  //164 / 178 = 0
    16'b10100100_10110011 : OUT <= 0;  //164 / 179 = 0
    16'b10100100_10110100 : OUT <= 0;  //164 / 180 = 0
    16'b10100100_10110101 : OUT <= 0;  //164 / 181 = 0
    16'b10100100_10110110 : OUT <= 0;  //164 / 182 = 0
    16'b10100100_10110111 : OUT <= 0;  //164 / 183 = 0
    16'b10100100_10111000 : OUT <= 0;  //164 / 184 = 0
    16'b10100100_10111001 : OUT <= 0;  //164 / 185 = 0
    16'b10100100_10111010 : OUT <= 0;  //164 / 186 = 0
    16'b10100100_10111011 : OUT <= 0;  //164 / 187 = 0
    16'b10100100_10111100 : OUT <= 0;  //164 / 188 = 0
    16'b10100100_10111101 : OUT <= 0;  //164 / 189 = 0
    16'b10100100_10111110 : OUT <= 0;  //164 / 190 = 0
    16'b10100100_10111111 : OUT <= 0;  //164 / 191 = 0
    16'b10100100_11000000 : OUT <= 0;  //164 / 192 = 0
    16'b10100100_11000001 : OUT <= 0;  //164 / 193 = 0
    16'b10100100_11000010 : OUT <= 0;  //164 / 194 = 0
    16'b10100100_11000011 : OUT <= 0;  //164 / 195 = 0
    16'b10100100_11000100 : OUT <= 0;  //164 / 196 = 0
    16'b10100100_11000101 : OUT <= 0;  //164 / 197 = 0
    16'b10100100_11000110 : OUT <= 0;  //164 / 198 = 0
    16'b10100100_11000111 : OUT <= 0;  //164 / 199 = 0
    16'b10100100_11001000 : OUT <= 0;  //164 / 200 = 0
    16'b10100100_11001001 : OUT <= 0;  //164 / 201 = 0
    16'b10100100_11001010 : OUT <= 0;  //164 / 202 = 0
    16'b10100100_11001011 : OUT <= 0;  //164 / 203 = 0
    16'b10100100_11001100 : OUT <= 0;  //164 / 204 = 0
    16'b10100100_11001101 : OUT <= 0;  //164 / 205 = 0
    16'b10100100_11001110 : OUT <= 0;  //164 / 206 = 0
    16'b10100100_11001111 : OUT <= 0;  //164 / 207 = 0
    16'b10100100_11010000 : OUT <= 0;  //164 / 208 = 0
    16'b10100100_11010001 : OUT <= 0;  //164 / 209 = 0
    16'b10100100_11010010 : OUT <= 0;  //164 / 210 = 0
    16'b10100100_11010011 : OUT <= 0;  //164 / 211 = 0
    16'b10100100_11010100 : OUT <= 0;  //164 / 212 = 0
    16'b10100100_11010101 : OUT <= 0;  //164 / 213 = 0
    16'b10100100_11010110 : OUT <= 0;  //164 / 214 = 0
    16'b10100100_11010111 : OUT <= 0;  //164 / 215 = 0
    16'b10100100_11011000 : OUT <= 0;  //164 / 216 = 0
    16'b10100100_11011001 : OUT <= 0;  //164 / 217 = 0
    16'b10100100_11011010 : OUT <= 0;  //164 / 218 = 0
    16'b10100100_11011011 : OUT <= 0;  //164 / 219 = 0
    16'b10100100_11011100 : OUT <= 0;  //164 / 220 = 0
    16'b10100100_11011101 : OUT <= 0;  //164 / 221 = 0
    16'b10100100_11011110 : OUT <= 0;  //164 / 222 = 0
    16'b10100100_11011111 : OUT <= 0;  //164 / 223 = 0
    16'b10100100_11100000 : OUT <= 0;  //164 / 224 = 0
    16'b10100100_11100001 : OUT <= 0;  //164 / 225 = 0
    16'b10100100_11100010 : OUT <= 0;  //164 / 226 = 0
    16'b10100100_11100011 : OUT <= 0;  //164 / 227 = 0
    16'b10100100_11100100 : OUT <= 0;  //164 / 228 = 0
    16'b10100100_11100101 : OUT <= 0;  //164 / 229 = 0
    16'b10100100_11100110 : OUT <= 0;  //164 / 230 = 0
    16'b10100100_11100111 : OUT <= 0;  //164 / 231 = 0
    16'b10100100_11101000 : OUT <= 0;  //164 / 232 = 0
    16'b10100100_11101001 : OUT <= 0;  //164 / 233 = 0
    16'b10100100_11101010 : OUT <= 0;  //164 / 234 = 0
    16'b10100100_11101011 : OUT <= 0;  //164 / 235 = 0
    16'b10100100_11101100 : OUT <= 0;  //164 / 236 = 0
    16'b10100100_11101101 : OUT <= 0;  //164 / 237 = 0
    16'b10100100_11101110 : OUT <= 0;  //164 / 238 = 0
    16'b10100100_11101111 : OUT <= 0;  //164 / 239 = 0
    16'b10100100_11110000 : OUT <= 0;  //164 / 240 = 0
    16'b10100100_11110001 : OUT <= 0;  //164 / 241 = 0
    16'b10100100_11110010 : OUT <= 0;  //164 / 242 = 0
    16'b10100100_11110011 : OUT <= 0;  //164 / 243 = 0
    16'b10100100_11110100 : OUT <= 0;  //164 / 244 = 0
    16'b10100100_11110101 : OUT <= 0;  //164 / 245 = 0
    16'b10100100_11110110 : OUT <= 0;  //164 / 246 = 0
    16'b10100100_11110111 : OUT <= 0;  //164 / 247 = 0
    16'b10100100_11111000 : OUT <= 0;  //164 / 248 = 0
    16'b10100100_11111001 : OUT <= 0;  //164 / 249 = 0
    16'b10100100_11111010 : OUT <= 0;  //164 / 250 = 0
    16'b10100100_11111011 : OUT <= 0;  //164 / 251 = 0
    16'b10100100_11111100 : OUT <= 0;  //164 / 252 = 0
    16'b10100100_11111101 : OUT <= 0;  //164 / 253 = 0
    16'b10100100_11111110 : OUT <= 0;  //164 / 254 = 0
    16'b10100100_11111111 : OUT <= 0;  //164 / 255 = 0
    16'b10100101_00000000 : OUT <= 0;  //165 / 0 = 0
    16'b10100101_00000001 : OUT <= 165;  //165 / 1 = 165
    16'b10100101_00000010 : OUT <= 82;  //165 / 2 = 82
    16'b10100101_00000011 : OUT <= 55;  //165 / 3 = 55
    16'b10100101_00000100 : OUT <= 41;  //165 / 4 = 41
    16'b10100101_00000101 : OUT <= 33;  //165 / 5 = 33
    16'b10100101_00000110 : OUT <= 27;  //165 / 6 = 27
    16'b10100101_00000111 : OUT <= 23;  //165 / 7 = 23
    16'b10100101_00001000 : OUT <= 20;  //165 / 8 = 20
    16'b10100101_00001001 : OUT <= 18;  //165 / 9 = 18
    16'b10100101_00001010 : OUT <= 16;  //165 / 10 = 16
    16'b10100101_00001011 : OUT <= 15;  //165 / 11 = 15
    16'b10100101_00001100 : OUT <= 13;  //165 / 12 = 13
    16'b10100101_00001101 : OUT <= 12;  //165 / 13 = 12
    16'b10100101_00001110 : OUT <= 11;  //165 / 14 = 11
    16'b10100101_00001111 : OUT <= 11;  //165 / 15 = 11
    16'b10100101_00010000 : OUT <= 10;  //165 / 16 = 10
    16'b10100101_00010001 : OUT <= 9;  //165 / 17 = 9
    16'b10100101_00010010 : OUT <= 9;  //165 / 18 = 9
    16'b10100101_00010011 : OUT <= 8;  //165 / 19 = 8
    16'b10100101_00010100 : OUT <= 8;  //165 / 20 = 8
    16'b10100101_00010101 : OUT <= 7;  //165 / 21 = 7
    16'b10100101_00010110 : OUT <= 7;  //165 / 22 = 7
    16'b10100101_00010111 : OUT <= 7;  //165 / 23 = 7
    16'b10100101_00011000 : OUT <= 6;  //165 / 24 = 6
    16'b10100101_00011001 : OUT <= 6;  //165 / 25 = 6
    16'b10100101_00011010 : OUT <= 6;  //165 / 26 = 6
    16'b10100101_00011011 : OUT <= 6;  //165 / 27 = 6
    16'b10100101_00011100 : OUT <= 5;  //165 / 28 = 5
    16'b10100101_00011101 : OUT <= 5;  //165 / 29 = 5
    16'b10100101_00011110 : OUT <= 5;  //165 / 30 = 5
    16'b10100101_00011111 : OUT <= 5;  //165 / 31 = 5
    16'b10100101_00100000 : OUT <= 5;  //165 / 32 = 5
    16'b10100101_00100001 : OUT <= 5;  //165 / 33 = 5
    16'b10100101_00100010 : OUT <= 4;  //165 / 34 = 4
    16'b10100101_00100011 : OUT <= 4;  //165 / 35 = 4
    16'b10100101_00100100 : OUT <= 4;  //165 / 36 = 4
    16'b10100101_00100101 : OUT <= 4;  //165 / 37 = 4
    16'b10100101_00100110 : OUT <= 4;  //165 / 38 = 4
    16'b10100101_00100111 : OUT <= 4;  //165 / 39 = 4
    16'b10100101_00101000 : OUT <= 4;  //165 / 40 = 4
    16'b10100101_00101001 : OUT <= 4;  //165 / 41 = 4
    16'b10100101_00101010 : OUT <= 3;  //165 / 42 = 3
    16'b10100101_00101011 : OUT <= 3;  //165 / 43 = 3
    16'b10100101_00101100 : OUT <= 3;  //165 / 44 = 3
    16'b10100101_00101101 : OUT <= 3;  //165 / 45 = 3
    16'b10100101_00101110 : OUT <= 3;  //165 / 46 = 3
    16'b10100101_00101111 : OUT <= 3;  //165 / 47 = 3
    16'b10100101_00110000 : OUT <= 3;  //165 / 48 = 3
    16'b10100101_00110001 : OUT <= 3;  //165 / 49 = 3
    16'b10100101_00110010 : OUT <= 3;  //165 / 50 = 3
    16'b10100101_00110011 : OUT <= 3;  //165 / 51 = 3
    16'b10100101_00110100 : OUT <= 3;  //165 / 52 = 3
    16'b10100101_00110101 : OUT <= 3;  //165 / 53 = 3
    16'b10100101_00110110 : OUT <= 3;  //165 / 54 = 3
    16'b10100101_00110111 : OUT <= 3;  //165 / 55 = 3
    16'b10100101_00111000 : OUT <= 2;  //165 / 56 = 2
    16'b10100101_00111001 : OUT <= 2;  //165 / 57 = 2
    16'b10100101_00111010 : OUT <= 2;  //165 / 58 = 2
    16'b10100101_00111011 : OUT <= 2;  //165 / 59 = 2
    16'b10100101_00111100 : OUT <= 2;  //165 / 60 = 2
    16'b10100101_00111101 : OUT <= 2;  //165 / 61 = 2
    16'b10100101_00111110 : OUT <= 2;  //165 / 62 = 2
    16'b10100101_00111111 : OUT <= 2;  //165 / 63 = 2
    16'b10100101_01000000 : OUT <= 2;  //165 / 64 = 2
    16'b10100101_01000001 : OUT <= 2;  //165 / 65 = 2
    16'b10100101_01000010 : OUT <= 2;  //165 / 66 = 2
    16'b10100101_01000011 : OUT <= 2;  //165 / 67 = 2
    16'b10100101_01000100 : OUT <= 2;  //165 / 68 = 2
    16'b10100101_01000101 : OUT <= 2;  //165 / 69 = 2
    16'b10100101_01000110 : OUT <= 2;  //165 / 70 = 2
    16'b10100101_01000111 : OUT <= 2;  //165 / 71 = 2
    16'b10100101_01001000 : OUT <= 2;  //165 / 72 = 2
    16'b10100101_01001001 : OUT <= 2;  //165 / 73 = 2
    16'b10100101_01001010 : OUT <= 2;  //165 / 74 = 2
    16'b10100101_01001011 : OUT <= 2;  //165 / 75 = 2
    16'b10100101_01001100 : OUT <= 2;  //165 / 76 = 2
    16'b10100101_01001101 : OUT <= 2;  //165 / 77 = 2
    16'b10100101_01001110 : OUT <= 2;  //165 / 78 = 2
    16'b10100101_01001111 : OUT <= 2;  //165 / 79 = 2
    16'b10100101_01010000 : OUT <= 2;  //165 / 80 = 2
    16'b10100101_01010001 : OUT <= 2;  //165 / 81 = 2
    16'b10100101_01010010 : OUT <= 2;  //165 / 82 = 2
    16'b10100101_01010011 : OUT <= 1;  //165 / 83 = 1
    16'b10100101_01010100 : OUT <= 1;  //165 / 84 = 1
    16'b10100101_01010101 : OUT <= 1;  //165 / 85 = 1
    16'b10100101_01010110 : OUT <= 1;  //165 / 86 = 1
    16'b10100101_01010111 : OUT <= 1;  //165 / 87 = 1
    16'b10100101_01011000 : OUT <= 1;  //165 / 88 = 1
    16'b10100101_01011001 : OUT <= 1;  //165 / 89 = 1
    16'b10100101_01011010 : OUT <= 1;  //165 / 90 = 1
    16'b10100101_01011011 : OUT <= 1;  //165 / 91 = 1
    16'b10100101_01011100 : OUT <= 1;  //165 / 92 = 1
    16'b10100101_01011101 : OUT <= 1;  //165 / 93 = 1
    16'b10100101_01011110 : OUT <= 1;  //165 / 94 = 1
    16'b10100101_01011111 : OUT <= 1;  //165 / 95 = 1
    16'b10100101_01100000 : OUT <= 1;  //165 / 96 = 1
    16'b10100101_01100001 : OUT <= 1;  //165 / 97 = 1
    16'b10100101_01100010 : OUT <= 1;  //165 / 98 = 1
    16'b10100101_01100011 : OUT <= 1;  //165 / 99 = 1
    16'b10100101_01100100 : OUT <= 1;  //165 / 100 = 1
    16'b10100101_01100101 : OUT <= 1;  //165 / 101 = 1
    16'b10100101_01100110 : OUT <= 1;  //165 / 102 = 1
    16'b10100101_01100111 : OUT <= 1;  //165 / 103 = 1
    16'b10100101_01101000 : OUT <= 1;  //165 / 104 = 1
    16'b10100101_01101001 : OUT <= 1;  //165 / 105 = 1
    16'b10100101_01101010 : OUT <= 1;  //165 / 106 = 1
    16'b10100101_01101011 : OUT <= 1;  //165 / 107 = 1
    16'b10100101_01101100 : OUT <= 1;  //165 / 108 = 1
    16'b10100101_01101101 : OUT <= 1;  //165 / 109 = 1
    16'b10100101_01101110 : OUT <= 1;  //165 / 110 = 1
    16'b10100101_01101111 : OUT <= 1;  //165 / 111 = 1
    16'b10100101_01110000 : OUT <= 1;  //165 / 112 = 1
    16'b10100101_01110001 : OUT <= 1;  //165 / 113 = 1
    16'b10100101_01110010 : OUT <= 1;  //165 / 114 = 1
    16'b10100101_01110011 : OUT <= 1;  //165 / 115 = 1
    16'b10100101_01110100 : OUT <= 1;  //165 / 116 = 1
    16'b10100101_01110101 : OUT <= 1;  //165 / 117 = 1
    16'b10100101_01110110 : OUT <= 1;  //165 / 118 = 1
    16'b10100101_01110111 : OUT <= 1;  //165 / 119 = 1
    16'b10100101_01111000 : OUT <= 1;  //165 / 120 = 1
    16'b10100101_01111001 : OUT <= 1;  //165 / 121 = 1
    16'b10100101_01111010 : OUT <= 1;  //165 / 122 = 1
    16'b10100101_01111011 : OUT <= 1;  //165 / 123 = 1
    16'b10100101_01111100 : OUT <= 1;  //165 / 124 = 1
    16'b10100101_01111101 : OUT <= 1;  //165 / 125 = 1
    16'b10100101_01111110 : OUT <= 1;  //165 / 126 = 1
    16'b10100101_01111111 : OUT <= 1;  //165 / 127 = 1
    16'b10100101_10000000 : OUT <= 1;  //165 / 128 = 1
    16'b10100101_10000001 : OUT <= 1;  //165 / 129 = 1
    16'b10100101_10000010 : OUT <= 1;  //165 / 130 = 1
    16'b10100101_10000011 : OUT <= 1;  //165 / 131 = 1
    16'b10100101_10000100 : OUT <= 1;  //165 / 132 = 1
    16'b10100101_10000101 : OUT <= 1;  //165 / 133 = 1
    16'b10100101_10000110 : OUT <= 1;  //165 / 134 = 1
    16'b10100101_10000111 : OUT <= 1;  //165 / 135 = 1
    16'b10100101_10001000 : OUT <= 1;  //165 / 136 = 1
    16'b10100101_10001001 : OUT <= 1;  //165 / 137 = 1
    16'b10100101_10001010 : OUT <= 1;  //165 / 138 = 1
    16'b10100101_10001011 : OUT <= 1;  //165 / 139 = 1
    16'b10100101_10001100 : OUT <= 1;  //165 / 140 = 1
    16'b10100101_10001101 : OUT <= 1;  //165 / 141 = 1
    16'b10100101_10001110 : OUT <= 1;  //165 / 142 = 1
    16'b10100101_10001111 : OUT <= 1;  //165 / 143 = 1
    16'b10100101_10010000 : OUT <= 1;  //165 / 144 = 1
    16'b10100101_10010001 : OUT <= 1;  //165 / 145 = 1
    16'b10100101_10010010 : OUT <= 1;  //165 / 146 = 1
    16'b10100101_10010011 : OUT <= 1;  //165 / 147 = 1
    16'b10100101_10010100 : OUT <= 1;  //165 / 148 = 1
    16'b10100101_10010101 : OUT <= 1;  //165 / 149 = 1
    16'b10100101_10010110 : OUT <= 1;  //165 / 150 = 1
    16'b10100101_10010111 : OUT <= 1;  //165 / 151 = 1
    16'b10100101_10011000 : OUT <= 1;  //165 / 152 = 1
    16'b10100101_10011001 : OUT <= 1;  //165 / 153 = 1
    16'b10100101_10011010 : OUT <= 1;  //165 / 154 = 1
    16'b10100101_10011011 : OUT <= 1;  //165 / 155 = 1
    16'b10100101_10011100 : OUT <= 1;  //165 / 156 = 1
    16'b10100101_10011101 : OUT <= 1;  //165 / 157 = 1
    16'b10100101_10011110 : OUT <= 1;  //165 / 158 = 1
    16'b10100101_10011111 : OUT <= 1;  //165 / 159 = 1
    16'b10100101_10100000 : OUT <= 1;  //165 / 160 = 1
    16'b10100101_10100001 : OUT <= 1;  //165 / 161 = 1
    16'b10100101_10100010 : OUT <= 1;  //165 / 162 = 1
    16'b10100101_10100011 : OUT <= 1;  //165 / 163 = 1
    16'b10100101_10100100 : OUT <= 1;  //165 / 164 = 1
    16'b10100101_10100101 : OUT <= 1;  //165 / 165 = 1
    16'b10100101_10100110 : OUT <= 0;  //165 / 166 = 0
    16'b10100101_10100111 : OUT <= 0;  //165 / 167 = 0
    16'b10100101_10101000 : OUT <= 0;  //165 / 168 = 0
    16'b10100101_10101001 : OUT <= 0;  //165 / 169 = 0
    16'b10100101_10101010 : OUT <= 0;  //165 / 170 = 0
    16'b10100101_10101011 : OUT <= 0;  //165 / 171 = 0
    16'b10100101_10101100 : OUT <= 0;  //165 / 172 = 0
    16'b10100101_10101101 : OUT <= 0;  //165 / 173 = 0
    16'b10100101_10101110 : OUT <= 0;  //165 / 174 = 0
    16'b10100101_10101111 : OUT <= 0;  //165 / 175 = 0
    16'b10100101_10110000 : OUT <= 0;  //165 / 176 = 0
    16'b10100101_10110001 : OUT <= 0;  //165 / 177 = 0
    16'b10100101_10110010 : OUT <= 0;  //165 / 178 = 0
    16'b10100101_10110011 : OUT <= 0;  //165 / 179 = 0
    16'b10100101_10110100 : OUT <= 0;  //165 / 180 = 0
    16'b10100101_10110101 : OUT <= 0;  //165 / 181 = 0
    16'b10100101_10110110 : OUT <= 0;  //165 / 182 = 0
    16'b10100101_10110111 : OUT <= 0;  //165 / 183 = 0
    16'b10100101_10111000 : OUT <= 0;  //165 / 184 = 0
    16'b10100101_10111001 : OUT <= 0;  //165 / 185 = 0
    16'b10100101_10111010 : OUT <= 0;  //165 / 186 = 0
    16'b10100101_10111011 : OUT <= 0;  //165 / 187 = 0
    16'b10100101_10111100 : OUT <= 0;  //165 / 188 = 0
    16'b10100101_10111101 : OUT <= 0;  //165 / 189 = 0
    16'b10100101_10111110 : OUT <= 0;  //165 / 190 = 0
    16'b10100101_10111111 : OUT <= 0;  //165 / 191 = 0
    16'b10100101_11000000 : OUT <= 0;  //165 / 192 = 0
    16'b10100101_11000001 : OUT <= 0;  //165 / 193 = 0
    16'b10100101_11000010 : OUT <= 0;  //165 / 194 = 0
    16'b10100101_11000011 : OUT <= 0;  //165 / 195 = 0
    16'b10100101_11000100 : OUT <= 0;  //165 / 196 = 0
    16'b10100101_11000101 : OUT <= 0;  //165 / 197 = 0
    16'b10100101_11000110 : OUT <= 0;  //165 / 198 = 0
    16'b10100101_11000111 : OUT <= 0;  //165 / 199 = 0
    16'b10100101_11001000 : OUT <= 0;  //165 / 200 = 0
    16'b10100101_11001001 : OUT <= 0;  //165 / 201 = 0
    16'b10100101_11001010 : OUT <= 0;  //165 / 202 = 0
    16'b10100101_11001011 : OUT <= 0;  //165 / 203 = 0
    16'b10100101_11001100 : OUT <= 0;  //165 / 204 = 0
    16'b10100101_11001101 : OUT <= 0;  //165 / 205 = 0
    16'b10100101_11001110 : OUT <= 0;  //165 / 206 = 0
    16'b10100101_11001111 : OUT <= 0;  //165 / 207 = 0
    16'b10100101_11010000 : OUT <= 0;  //165 / 208 = 0
    16'b10100101_11010001 : OUT <= 0;  //165 / 209 = 0
    16'b10100101_11010010 : OUT <= 0;  //165 / 210 = 0
    16'b10100101_11010011 : OUT <= 0;  //165 / 211 = 0
    16'b10100101_11010100 : OUT <= 0;  //165 / 212 = 0
    16'b10100101_11010101 : OUT <= 0;  //165 / 213 = 0
    16'b10100101_11010110 : OUT <= 0;  //165 / 214 = 0
    16'b10100101_11010111 : OUT <= 0;  //165 / 215 = 0
    16'b10100101_11011000 : OUT <= 0;  //165 / 216 = 0
    16'b10100101_11011001 : OUT <= 0;  //165 / 217 = 0
    16'b10100101_11011010 : OUT <= 0;  //165 / 218 = 0
    16'b10100101_11011011 : OUT <= 0;  //165 / 219 = 0
    16'b10100101_11011100 : OUT <= 0;  //165 / 220 = 0
    16'b10100101_11011101 : OUT <= 0;  //165 / 221 = 0
    16'b10100101_11011110 : OUT <= 0;  //165 / 222 = 0
    16'b10100101_11011111 : OUT <= 0;  //165 / 223 = 0
    16'b10100101_11100000 : OUT <= 0;  //165 / 224 = 0
    16'b10100101_11100001 : OUT <= 0;  //165 / 225 = 0
    16'b10100101_11100010 : OUT <= 0;  //165 / 226 = 0
    16'b10100101_11100011 : OUT <= 0;  //165 / 227 = 0
    16'b10100101_11100100 : OUT <= 0;  //165 / 228 = 0
    16'b10100101_11100101 : OUT <= 0;  //165 / 229 = 0
    16'b10100101_11100110 : OUT <= 0;  //165 / 230 = 0
    16'b10100101_11100111 : OUT <= 0;  //165 / 231 = 0
    16'b10100101_11101000 : OUT <= 0;  //165 / 232 = 0
    16'b10100101_11101001 : OUT <= 0;  //165 / 233 = 0
    16'b10100101_11101010 : OUT <= 0;  //165 / 234 = 0
    16'b10100101_11101011 : OUT <= 0;  //165 / 235 = 0
    16'b10100101_11101100 : OUT <= 0;  //165 / 236 = 0
    16'b10100101_11101101 : OUT <= 0;  //165 / 237 = 0
    16'b10100101_11101110 : OUT <= 0;  //165 / 238 = 0
    16'b10100101_11101111 : OUT <= 0;  //165 / 239 = 0
    16'b10100101_11110000 : OUT <= 0;  //165 / 240 = 0
    16'b10100101_11110001 : OUT <= 0;  //165 / 241 = 0
    16'b10100101_11110010 : OUT <= 0;  //165 / 242 = 0
    16'b10100101_11110011 : OUT <= 0;  //165 / 243 = 0
    16'b10100101_11110100 : OUT <= 0;  //165 / 244 = 0
    16'b10100101_11110101 : OUT <= 0;  //165 / 245 = 0
    16'b10100101_11110110 : OUT <= 0;  //165 / 246 = 0
    16'b10100101_11110111 : OUT <= 0;  //165 / 247 = 0
    16'b10100101_11111000 : OUT <= 0;  //165 / 248 = 0
    16'b10100101_11111001 : OUT <= 0;  //165 / 249 = 0
    16'b10100101_11111010 : OUT <= 0;  //165 / 250 = 0
    16'b10100101_11111011 : OUT <= 0;  //165 / 251 = 0
    16'b10100101_11111100 : OUT <= 0;  //165 / 252 = 0
    16'b10100101_11111101 : OUT <= 0;  //165 / 253 = 0
    16'b10100101_11111110 : OUT <= 0;  //165 / 254 = 0
    16'b10100101_11111111 : OUT <= 0;  //165 / 255 = 0
    16'b10100110_00000000 : OUT <= 0;  //166 / 0 = 0
    16'b10100110_00000001 : OUT <= 166;  //166 / 1 = 166
    16'b10100110_00000010 : OUT <= 83;  //166 / 2 = 83
    16'b10100110_00000011 : OUT <= 55;  //166 / 3 = 55
    16'b10100110_00000100 : OUT <= 41;  //166 / 4 = 41
    16'b10100110_00000101 : OUT <= 33;  //166 / 5 = 33
    16'b10100110_00000110 : OUT <= 27;  //166 / 6 = 27
    16'b10100110_00000111 : OUT <= 23;  //166 / 7 = 23
    16'b10100110_00001000 : OUT <= 20;  //166 / 8 = 20
    16'b10100110_00001001 : OUT <= 18;  //166 / 9 = 18
    16'b10100110_00001010 : OUT <= 16;  //166 / 10 = 16
    16'b10100110_00001011 : OUT <= 15;  //166 / 11 = 15
    16'b10100110_00001100 : OUT <= 13;  //166 / 12 = 13
    16'b10100110_00001101 : OUT <= 12;  //166 / 13 = 12
    16'b10100110_00001110 : OUT <= 11;  //166 / 14 = 11
    16'b10100110_00001111 : OUT <= 11;  //166 / 15 = 11
    16'b10100110_00010000 : OUT <= 10;  //166 / 16 = 10
    16'b10100110_00010001 : OUT <= 9;  //166 / 17 = 9
    16'b10100110_00010010 : OUT <= 9;  //166 / 18 = 9
    16'b10100110_00010011 : OUT <= 8;  //166 / 19 = 8
    16'b10100110_00010100 : OUT <= 8;  //166 / 20 = 8
    16'b10100110_00010101 : OUT <= 7;  //166 / 21 = 7
    16'b10100110_00010110 : OUT <= 7;  //166 / 22 = 7
    16'b10100110_00010111 : OUT <= 7;  //166 / 23 = 7
    16'b10100110_00011000 : OUT <= 6;  //166 / 24 = 6
    16'b10100110_00011001 : OUT <= 6;  //166 / 25 = 6
    16'b10100110_00011010 : OUT <= 6;  //166 / 26 = 6
    16'b10100110_00011011 : OUT <= 6;  //166 / 27 = 6
    16'b10100110_00011100 : OUT <= 5;  //166 / 28 = 5
    16'b10100110_00011101 : OUT <= 5;  //166 / 29 = 5
    16'b10100110_00011110 : OUT <= 5;  //166 / 30 = 5
    16'b10100110_00011111 : OUT <= 5;  //166 / 31 = 5
    16'b10100110_00100000 : OUT <= 5;  //166 / 32 = 5
    16'b10100110_00100001 : OUT <= 5;  //166 / 33 = 5
    16'b10100110_00100010 : OUT <= 4;  //166 / 34 = 4
    16'b10100110_00100011 : OUT <= 4;  //166 / 35 = 4
    16'b10100110_00100100 : OUT <= 4;  //166 / 36 = 4
    16'b10100110_00100101 : OUT <= 4;  //166 / 37 = 4
    16'b10100110_00100110 : OUT <= 4;  //166 / 38 = 4
    16'b10100110_00100111 : OUT <= 4;  //166 / 39 = 4
    16'b10100110_00101000 : OUT <= 4;  //166 / 40 = 4
    16'b10100110_00101001 : OUT <= 4;  //166 / 41 = 4
    16'b10100110_00101010 : OUT <= 3;  //166 / 42 = 3
    16'b10100110_00101011 : OUT <= 3;  //166 / 43 = 3
    16'b10100110_00101100 : OUT <= 3;  //166 / 44 = 3
    16'b10100110_00101101 : OUT <= 3;  //166 / 45 = 3
    16'b10100110_00101110 : OUT <= 3;  //166 / 46 = 3
    16'b10100110_00101111 : OUT <= 3;  //166 / 47 = 3
    16'b10100110_00110000 : OUT <= 3;  //166 / 48 = 3
    16'b10100110_00110001 : OUT <= 3;  //166 / 49 = 3
    16'b10100110_00110010 : OUT <= 3;  //166 / 50 = 3
    16'b10100110_00110011 : OUT <= 3;  //166 / 51 = 3
    16'b10100110_00110100 : OUT <= 3;  //166 / 52 = 3
    16'b10100110_00110101 : OUT <= 3;  //166 / 53 = 3
    16'b10100110_00110110 : OUT <= 3;  //166 / 54 = 3
    16'b10100110_00110111 : OUT <= 3;  //166 / 55 = 3
    16'b10100110_00111000 : OUT <= 2;  //166 / 56 = 2
    16'b10100110_00111001 : OUT <= 2;  //166 / 57 = 2
    16'b10100110_00111010 : OUT <= 2;  //166 / 58 = 2
    16'b10100110_00111011 : OUT <= 2;  //166 / 59 = 2
    16'b10100110_00111100 : OUT <= 2;  //166 / 60 = 2
    16'b10100110_00111101 : OUT <= 2;  //166 / 61 = 2
    16'b10100110_00111110 : OUT <= 2;  //166 / 62 = 2
    16'b10100110_00111111 : OUT <= 2;  //166 / 63 = 2
    16'b10100110_01000000 : OUT <= 2;  //166 / 64 = 2
    16'b10100110_01000001 : OUT <= 2;  //166 / 65 = 2
    16'b10100110_01000010 : OUT <= 2;  //166 / 66 = 2
    16'b10100110_01000011 : OUT <= 2;  //166 / 67 = 2
    16'b10100110_01000100 : OUT <= 2;  //166 / 68 = 2
    16'b10100110_01000101 : OUT <= 2;  //166 / 69 = 2
    16'b10100110_01000110 : OUT <= 2;  //166 / 70 = 2
    16'b10100110_01000111 : OUT <= 2;  //166 / 71 = 2
    16'b10100110_01001000 : OUT <= 2;  //166 / 72 = 2
    16'b10100110_01001001 : OUT <= 2;  //166 / 73 = 2
    16'b10100110_01001010 : OUT <= 2;  //166 / 74 = 2
    16'b10100110_01001011 : OUT <= 2;  //166 / 75 = 2
    16'b10100110_01001100 : OUT <= 2;  //166 / 76 = 2
    16'b10100110_01001101 : OUT <= 2;  //166 / 77 = 2
    16'b10100110_01001110 : OUT <= 2;  //166 / 78 = 2
    16'b10100110_01001111 : OUT <= 2;  //166 / 79 = 2
    16'b10100110_01010000 : OUT <= 2;  //166 / 80 = 2
    16'b10100110_01010001 : OUT <= 2;  //166 / 81 = 2
    16'b10100110_01010010 : OUT <= 2;  //166 / 82 = 2
    16'b10100110_01010011 : OUT <= 2;  //166 / 83 = 2
    16'b10100110_01010100 : OUT <= 1;  //166 / 84 = 1
    16'b10100110_01010101 : OUT <= 1;  //166 / 85 = 1
    16'b10100110_01010110 : OUT <= 1;  //166 / 86 = 1
    16'b10100110_01010111 : OUT <= 1;  //166 / 87 = 1
    16'b10100110_01011000 : OUT <= 1;  //166 / 88 = 1
    16'b10100110_01011001 : OUT <= 1;  //166 / 89 = 1
    16'b10100110_01011010 : OUT <= 1;  //166 / 90 = 1
    16'b10100110_01011011 : OUT <= 1;  //166 / 91 = 1
    16'b10100110_01011100 : OUT <= 1;  //166 / 92 = 1
    16'b10100110_01011101 : OUT <= 1;  //166 / 93 = 1
    16'b10100110_01011110 : OUT <= 1;  //166 / 94 = 1
    16'b10100110_01011111 : OUT <= 1;  //166 / 95 = 1
    16'b10100110_01100000 : OUT <= 1;  //166 / 96 = 1
    16'b10100110_01100001 : OUT <= 1;  //166 / 97 = 1
    16'b10100110_01100010 : OUT <= 1;  //166 / 98 = 1
    16'b10100110_01100011 : OUT <= 1;  //166 / 99 = 1
    16'b10100110_01100100 : OUT <= 1;  //166 / 100 = 1
    16'b10100110_01100101 : OUT <= 1;  //166 / 101 = 1
    16'b10100110_01100110 : OUT <= 1;  //166 / 102 = 1
    16'b10100110_01100111 : OUT <= 1;  //166 / 103 = 1
    16'b10100110_01101000 : OUT <= 1;  //166 / 104 = 1
    16'b10100110_01101001 : OUT <= 1;  //166 / 105 = 1
    16'b10100110_01101010 : OUT <= 1;  //166 / 106 = 1
    16'b10100110_01101011 : OUT <= 1;  //166 / 107 = 1
    16'b10100110_01101100 : OUT <= 1;  //166 / 108 = 1
    16'b10100110_01101101 : OUT <= 1;  //166 / 109 = 1
    16'b10100110_01101110 : OUT <= 1;  //166 / 110 = 1
    16'b10100110_01101111 : OUT <= 1;  //166 / 111 = 1
    16'b10100110_01110000 : OUT <= 1;  //166 / 112 = 1
    16'b10100110_01110001 : OUT <= 1;  //166 / 113 = 1
    16'b10100110_01110010 : OUT <= 1;  //166 / 114 = 1
    16'b10100110_01110011 : OUT <= 1;  //166 / 115 = 1
    16'b10100110_01110100 : OUT <= 1;  //166 / 116 = 1
    16'b10100110_01110101 : OUT <= 1;  //166 / 117 = 1
    16'b10100110_01110110 : OUT <= 1;  //166 / 118 = 1
    16'b10100110_01110111 : OUT <= 1;  //166 / 119 = 1
    16'b10100110_01111000 : OUT <= 1;  //166 / 120 = 1
    16'b10100110_01111001 : OUT <= 1;  //166 / 121 = 1
    16'b10100110_01111010 : OUT <= 1;  //166 / 122 = 1
    16'b10100110_01111011 : OUT <= 1;  //166 / 123 = 1
    16'b10100110_01111100 : OUT <= 1;  //166 / 124 = 1
    16'b10100110_01111101 : OUT <= 1;  //166 / 125 = 1
    16'b10100110_01111110 : OUT <= 1;  //166 / 126 = 1
    16'b10100110_01111111 : OUT <= 1;  //166 / 127 = 1
    16'b10100110_10000000 : OUT <= 1;  //166 / 128 = 1
    16'b10100110_10000001 : OUT <= 1;  //166 / 129 = 1
    16'b10100110_10000010 : OUT <= 1;  //166 / 130 = 1
    16'b10100110_10000011 : OUT <= 1;  //166 / 131 = 1
    16'b10100110_10000100 : OUT <= 1;  //166 / 132 = 1
    16'b10100110_10000101 : OUT <= 1;  //166 / 133 = 1
    16'b10100110_10000110 : OUT <= 1;  //166 / 134 = 1
    16'b10100110_10000111 : OUT <= 1;  //166 / 135 = 1
    16'b10100110_10001000 : OUT <= 1;  //166 / 136 = 1
    16'b10100110_10001001 : OUT <= 1;  //166 / 137 = 1
    16'b10100110_10001010 : OUT <= 1;  //166 / 138 = 1
    16'b10100110_10001011 : OUT <= 1;  //166 / 139 = 1
    16'b10100110_10001100 : OUT <= 1;  //166 / 140 = 1
    16'b10100110_10001101 : OUT <= 1;  //166 / 141 = 1
    16'b10100110_10001110 : OUT <= 1;  //166 / 142 = 1
    16'b10100110_10001111 : OUT <= 1;  //166 / 143 = 1
    16'b10100110_10010000 : OUT <= 1;  //166 / 144 = 1
    16'b10100110_10010001 : OUT <= 1;  //166 / 145 = 1
    16'b10100110_10010010 : OUT <= 1;  //166 / 146 = 1
    16'b10100110_10010011 : OUT <= 1;  //166 / 147 = 1
    16'b10100110_10010100 : OUT <= 1;  //166 / 148 = 1
    16'b10100110_10010101 : OUT <= 1;  //166 / 149 = 1
    16'b10100110_10010110 : OUT <= 1;  //166 / 150 = 1
    16'b10100110_10010111 : OUT <= 1;  //166 / 151 = 1
    16'b10100110_10011000 : OUT <= 1;  //166 / 152 = 1
    16'b10100110_10011001 : OUT <= 1;  //166 / 153 = 1
    16'b10100110_10011010 : OUT <= 1;  //166 / 154 = 1
    16'b10100110_10011011 : OUT <= 1;  //166 / 155 = 1
    16'b10100110_10011100 : OUT <= 1;  //166 / 156 = 1
    16'b10100110_10011101 : OUT <= 1;  //166 / 157 = 1
    16'b10100110_10011110 : OUT <= 1;  //166 / 158 = 1
    16'b10100110_10011111 : OUT <= 1;  //166 / 159 = 1
    16'b10100110_10100000 : OUT <= 1;  //166 / 160 = 1
    16'b10100110_10100001 : OUT <= 1;  //166 / 161 = 1
    16'b10100110_10100010 : OUT <= 1;  //166 / 162 = 1
    16'b10100110_10100011 : OUT <= 1;  //166 / 163 = 1
    16'b10100110_10100100 : OUT <= 1;  //166 / 164 = 1
    16'b10100110_10100101 : OUT <= 1;  //166 / 165 = 1
    16'b10100110_10100110 : OUT <= 1;  //166 / 166 = 1
    16'b10100110_10100111 : OUT <= 0;  //166 / 167 = 0
    16'b10100110_10101000 : OUT <= 0;  //166 / 168 = 0
    16'b10100110_10101001 : OUT <= 0;  //166 / 169 = 0
    16'b10100110_10101010 : OUT <= 0;  //166 / 170 = 0
    16'b10100110_10101011 : OUT <= 0;  //166 / 171 = 0
    16'b10100110_10101100 : OUT <= 0;  //166 / 172 = 0
    16'b10100110_10101101 : OUT <= 0;  //166 / 173 = 0
    16'b10100110_10101110 : OUT <= 0;  //166 / 174 = 0
    16'b10100110_10101111 : OUT <= 0;  //166 / 175 = 0
    16'b10100110_10110000 : OUT <= 0;  //166 / 176 = 0
    16'b10100110_10110001 : OUT <= 0;  //166 / 177 = 0
    16'b10100110_10110010 : OUT <= 0;  //166 / 178 = 0
    16'b10100110_10110011 : OUT <= 0;  //166 / 179 = 0
    16'b10100110_10110100 : OUT <= 0;  //166 / 180 = 0
    16'b10100110_10110101 : OUT <= 0;  //166 / 181 = 0
    16'b10100110_10110110 : OUT <= 0;  //166 / 182 = 0
    16'b10100110_10110111 : OUT <= 0;  //166 / 183 = 0
    16'b10100110_10111000 : OUT <= 0;  //166 / 184 = 0
    16'b10100110_10111001 : OUT <= 0;  //166 / 185 = 0
    16'b10100110_10111010 : OUT <= 0;  //166 / 186 = 0
    16'b10100110_10111011 : OUT <= 0;  //166 / 187 = 0
    16'b10100110_10111100 : OUT <= 0;  //166 / 188 = 0
    16'b10100110_10111101 : OUT <= 0;  //166 / 189 = 0
    16'b10100110_10111110 : OUT <= 0;  //166 / 190 = 0
    16'b10100110_10111111 : OUT <= 0;  //166 / 191 = 0
    16'b10100110_11000000 : OUT <= 0;  //166 / 192 = 0
    16'b10100110_11000001 : OUT <= 0;  //166 / 193 = 0
    16'b10100110_11000010 : OUT <= 0;  //166 / 194 = 0
    16'b10100110_11000011 : OUT <= 0;  //166 / 195 = 0
    16'b10100110_11000100 : OUT <= 0;  //166 / 196 = 0
    16'b10100110_11000101 : OUT <= 0;  //166 / 197 = 0
    16'b10100110_11000110 : OUT <= 0;  //166 / 198 = 0
    16'b10100110_11000111 : OUT <= 0;  //166 / 199 = 0
    16'b10100110_11001000 : OUT <= 0;  //166 / 200 = 0
    16'b10100110_11001001 : OUT <= 0;  //166 / 201 = 0
    16'b10100110_11001010 : OUT <= 0;  //166 / 202 = 0
    16'b10100110_11001011 : OUT <= 0;  //166 / 203 = 0
    16'b10100110_11001100 : OUT <= 0;  //166 / 204 = 0
    16'b10100110_11001101 : OUT <= 0;  //166 / 205 = 0
    16'b10100110_11001110 : OUT <= 0;  //166 / 206 = 0
    16'b10100110_11001111 : OUT <= 0;  //166 / 207 = 0
    16'b10100110_11010000 : OUT <= 0;  //166 / 208 = 0
    16'b10100110_11010001 : OUT <= 0;  //166 / 209 = 0
    16'b10100110_11010010 : OUT <= 0;  //166 / 210 = 0
    16'b10100110_11010011 : OUT <= 0;  //166 / 211 = 0
    16'b10100110_11010100 : OUT <= 0;  //166 / 212 = 0
    16'b10100110_11010101 : OUT <= 0;  //166 / 213 = 0
    16'b10100110_11010110 : OUT <= 0;  //166 / 214 = 0
    16'b10100110_11010111 : OUT <= 0;  //166 / 215 = 0
    16'b10100110_11011000 : OUT <= 0;  //166 / 216 = 0
    16'b10100110_11011001 : OUT <= 0;  //166 / 217 = 0
    16'b10100110_11011010 : OUT <= 0;  //166 / 218 = 0
    16'b10100110_11011011 : OUT <= 0;  //166 / 219 = 0
    16'b10100110_11011100 : OUT <= 0;  //166 / 220 = 0
    16'b10100110_11011101 : OUT <= 0;  //166 / 221 = 0
    16'b10100110_11011110 : OUT <= 0;  //166 / 222 = 0
    16'b10100110_11011111 : OUT <= 0;  //166 / 223 = 0
    16'b10100110_11100000 : OUT <= 0;  //166 / 224 = 0
    16'b10100110_11100001 : OUT <= 0;  //166 / 225 = 0
    16'b10100110_11100010 : OUT <= 0;  //166 / 226 = 0
    16'b10100110_11100011 : OUT <= 0;  //166 / 227 = 0
    16'b10100110_11100100 : OUT <= 0;  //166 / 228 = 0
    16'b10100110_11100101 : OUT <= 0;  //166 / 229 = 0
    16'b10100110_11100110 : OUT <= 0;  //166 / 230 = 0
    16'b10100110_11100111 : OUT <= 0;  //166 / 231 = 0
    16'b10100110_11101000 : OUT <= 0;  //166 / 232 = 0
    16'b10100110_11101001 : OUT <= 0;  //166 / 233 = 0
    16'b10100110_11101010 : OUT <= 0;  //166 / 234 = 0
    16'b10100110_11101011 : OUT <= 0;  //166 / 235 = 0
    16'b10100110_11101100 : OUT <= 0;  //166 / 236 = 0
    16'b10100110_11101101 : OUT <= 0;  //166 / 237 = 0
    16'b10100110_11101110 : OUT <= 0;  //166 / 238 = 0
    16'b10100110_11101111 : OUT <= 0;  //166 / 239 = 0
    16'b10100110_11110000 : OUT <= 0;  //166 / 240 = 0
    16'b10100110_11110001 : OUT <= 0;  //166 / 241 = 0
    16'b10100110_11110010 : OUT <= 0;  //166 / 242 = 0
    16'b10100110_11110011 : OUT <= 0;  //166 / 243 = 0
    16'b10100110_11110100 : OUT <= 0;  //166 / 244 = 0
    16'b10100110_11110101 : OUT <= 0;  //166 / 245 = 0
    16'b10100110_11110110 : OUT <= 0;  //166 / 246 = 0
    16'b10100110_11110111 : OUT <= 0;  //166 / 247 = 0
    16'b10100110_11111000 : OUT <= 0;  //166 / 248 = 0
    16'b10100110_11111001 : OUT <= 0;  //166 / 249 = 0
    16'b10100110_11111010 : OUT <= 0;  //166 / 250 = 0
    16'b10100110_11111011 : OUT <= 0;  //166 / 251 = 0
    16'b10100110_11111100 : OUT <= 0;  //166 / 252 = 0
    16'b10100110_11111101 : OUT <= 0;  //166 / 253 = 0
    16'b10100110_11111110 : OUT <= 0;  //166 / 254 = 0
    16'b10100110_11111111 : OUT <= 0;  //166 / 255 = 0
    16'b10100111_00000000 : OUT <= 0;  //167 / 0 = 0
    16'b10100111_00000001 : OUT <= 167;  //167 / 1 = 167
    16'b10100111_00000010 : OUT <= 83;  //167 / 2 = 83
    16'b10100111_00000011 : OUT <= 55;  //167 / 3 = 55
    16'b10100111_00000100 : OUT <= 41;  //167 / 4 = 41
    16'b10100111_00000101 : OUT <= 33;  //167 / 5 = 33
    16'b10100111_00000110 : OUT <= 27;  //167 / 6 = 27
    16'b10100111_00000111 : OUT <= 23;  //167 / 7 = 23
    16'b10100111_00001000 : OUT <= 20;  //167 / 8 = 20
    16'b10100111_00001001 : OUT <= 18;  //167 / 9 = 18
    16'b10100111_00001010 : OUT <= 16;  //167 / 10 = 16
    16'b10100111_00001011 : OUT <= 15;  //167 / 11 = 15
    16'b10100111_00001100 : OUT <= 13;  //167 / 12 = 13
    16'b10100111_00001101 : OUT <= 12;  //167 / 13 = 12
    16'b10100111_00001110 : OUT <= 11;  //167 / 14 = 11
    16'b10100111_00001111 : OUT <= 11;  //167 / 15 = 11
    16'b10100111_00010000 : OUT <= 10;  //167 / 16 = 10
    16'b10100111_00010001 : OUT <= 9;  //167 / 17 = 9
    16'b10100111_00010010 : OUT <= 9;  //167 / 18 = 9
    16'b10100111_00010011 : OUT <= 8;  //167 / 19 = 8
    16'b10100111_00010100 : OUT <= 8;  //167 / 20 = 8
    16'b10100111_00010101 : OUT <= 7;  //167 / 21 = 7
    16'b10100111_00010110 : OUT <= 7;  //167 / 22 = 7
    16'b10100111_00010111 : OUT <= 7;  //167 / 23 = 7
    16'b10100111_00011000 : OUT <= 6;  //167 / 24 = 6
    16'b10100111_00011001 : OUT <= 6;  //167 / 25 = 6
    16'b10100111_00011010 : OUT <= 6;  //167 / 26 = 6
    16'b10100111_00011011 : OUT <= 6;  //167 / 27 = 6
    16'b10100111_00011100 : OUT <= 5;  //167 / 28 = 5
    16'b10100111_00011101 : OUT <= 5;  //167 / 29 = 5
    16'b10100111_00011110 : OUT <= 5;  //167 / 30 = 5
    16'b10100111_00011111 : OUT <= 5;  //167 / 31 = 5
    16'b10100111_00100000 : OUT <= 5;  //167 / 32 = 5
    16'b10100111_00100001 : OUT <= 5;  //167 / 33 = 5
    16'b10100111_00100010 : OUT <= 4;  //167 / 34 = 4
    16'b10100111_00100011 : OUT <= 4;  //167 / 35 = 4
    16'b10100111_00100100 : OUT <= 4;  //167 / 36 = 4
    16'b10100111_00100101 : OUT <= 4;  //167 / 37 = 4
    16'b10100111_00100110 : OUT <= 4;  //167 / 38 = 4
    16'b10100111_00100111 : OUT <= 4;  //167 / 39 = 4
    16'b10100111_00101000 : OUT <= 4;  //167 / 40 = 4
    16'b10100111_00101001 : OUT <= 4;  //167 / 41 = 4
    16'b10100111_00101010 : OUT <= 3;  //167 / 42 = 3
    16'b10100111_00101011 : OUT <= 3;  //167 / 43 = 3
    16'b10100111_00101100 : OUT <= 3;  //167 / 44 = 3
    16'b10100111_00101101 : OUT <= 3;  //167 / 45 = 3
    16'b10100111_00101110 : OUT <= 3;  //167 / 46 = 3
    16'b10100111_00101111 : OUT <= 3;  //167 / 47 = 3
    16'b10100111_00110000 : OUT <= 3;  //167 / 48 = 3
    16'b10100111_00110001 : OUT <= 3;  //167 / 49 = 3
    16'b10100111_00110010 : OUT <= 3;  //167 / 50 = 3
    16'b10100111_00110011 : OUT <= 3;  //167 / 51 = 3
    16'b10100111_00110100 : OUT <= 3;  //167 / 52 = 3
    16'b10100111_00110101 : OUT <= 3;  //167 / 53 = 3
    16'b10100111_00110110 : OUT <= 3;  //167 / 54 = 3
    16'b10100111_00110111 : OUT <= 3;  //167 / 55 = 3
    16'b10100111_00111000 : OUT <= 2;  //167 / 56 = 2
    16'b10100111_00111001 : OUT <= 2;  //167 / 57 = 2
    16'b10100111_00111010 : OUT <= 2;  //167 / 58 = 2
    16'b10100111_00111011 : OUT <= 2;  //167 / 59 = 2
    16'b10100111_00111100 : OUT <= 2;  //167 / 60 = 2
    16'b10100111_00111101 : OUT <= 2;  //167 / 61 = 2
    16'b10100111_00111110 : OUT <= 2;  //167 / 62 = 2
    16'b10100111_00111111 : OUT <= 2;  //167 / 63 = 2
    16'b10100111_01000000 : OUT <= 2;  //167 / 64 = 2
    16'b10100111_01000001 : OUT <= 2;  //167 / 65 = 2
    16'b10100111_01000010 : OUT <= 2;  //167 / 66 = 2
    16'b10100111_01000011 : OUT <= 2;  //167 / 67 = 2
    16'b10100111_01000100 : OUT <= 2;  //167 / 68 = 2
    16'b10100111_01000101 : OUT <= 2;  //167 / 69 = 2
    16'b10100111_01000110 : OUT <= 2;  //167 / 70 = 2
    16'b10100111_01000111 : OUT <= 2;  //167 / 71 = 2
    16'b10100111_01001000 : OUT <= 2;  //167 / 72 = 2
    16'b10100111_01001001 : OUT <= 2;  //167 / 73 = 2
    16'b10100111_01001010 : OUT <= 2;  //167 / 74 = 2
    16'b10100111_01001011 : OUT <= 2;  //167 / 75 = 2
    16'b10100111_01001100 : OUT <= 2;  //167 / 76 = 2
    16'b10100111_01001101 : OUT <= 2;  //167 / 77 = 2
    16'b10100111_01001110 : OUT <= 2;  //167 / 78 = 2
    16'b10100111_01001111 : OUT <= 2;  //167 / 79 = 2
    16'b10100111_01010000 : OUT <= 2;  //167 / 80 = 2
    16'b10100111_01010001 : OUT <= 2;  //167 / 81 = 2
    16'b10100111_01010010 : OUT <= 2;  //167 / 82 = 2
    16'b10100111_01010011 : OUT <= 2;  //167 / 83 = 2
    16'b10100111_01010100 : OUT <= 1;  //167 / 84 = 1
    16'b10100111_01010101 : OUT <= 1;  //167 / 85 = 1
    16'b10100111_01010110 : OUT <= 1;  //167 / 86 = 1
    16'b10100111_01010111 : OUT <= 1;  //167 / 87 = 1
    16'b10100111_01011000 : OUT <= 1;  //167 / 88 = 1
    16'b10100111_01011001 : OUT <= 1;  //167 / 89 = 1
    16'b10100111_01011010 : OUT <= 1;  //167 / 90 = 1
    16'b10100111_01011011 : OUT <= 1;  //167 / 91 = 1
    16'b10100111_01011100 : OUT <= 1;  //167 / 92 = 1
    16'b10100111_01011101 : OUT <= 1;  //167 / 93 = 1
    16'b10100111_01011110 : OUT <= 1;  //167 / 94 = 1
    16'b10100111_01011111 : OUT <= 1;  //167 / 95 = 1
    16'b10100111_01100000 : OUT <= 1;  //167 / 96 = 1
    16'b10100111_01100001 : OUT <= 1;  //167 / 97 = 1
    16'b10100111_01100010 : OUT <= 1;  //167 / 98 = 1
    16'b10100111_01100011 : OUT <= 1;  //167 / 99 = 1
    16'b10100111_01100100 : OUT <= 1;  //167 / 100 = 1
    16'b10100111_01100101 : OUT <= 1;  //167 / 101 = 1
    16'b10100111_01100110 : OUT <= 1;  //167 / 102 = 1
    16'b10100111_01100111 : OUT <= 1;  //167 / 103 = 1
    16'b10100111_01101000 : OUT <= 1;  //167 / 104 = 1
    16'b10100111_01101001 : OUT <= 1;  //167 / 105 = 1
    16'b10100111_01101010 : OUT <= 1;  //167 / 106 = 1
    16'b10100111_01101011 : OUT <= 1;  //167 / 107 = 1
    16'b10100111_01101100 : OUT <= 1;  //167 / 108 = 1
    16'b10100111_01101101 : OUT <= 1;  //167 / 109 = 1
    16'b10100111_01101110 : OUT <= 1;  //167 / 110 = 1
    16'b10100111_01101111 : OUT <= 1;  //167 / 111 = 1
    16'b10100111_01110000 : OUT <= 1;  //167 / 112 = 1
    16'b10100111_01110001 : OUT <= 1;  //167 / 113 = 1
    16'b10100111_01110010 : OUT <= 1;  //167 / 114 = 1
    16'b10100111_01110011 : OUT <= 1;  //167 / 115 = 1
    16'b10100111_01110100 : OUT <= 1;  //167 / 116 = 1
    16'b10100111_01110101 : OUT <= 1;  //167 / 117 = 1
    16'b10100111_01110110 : OUT <= 1;  //167 / 118 = 1
    16'b10100111_01110111 : OUT <= 1;  //167 / 119 = 1
    16'b10100111_01111000 : OUT <= 1;  //167 / 120 = 1
    16'b10100111_01111001 : OUT <= 1;  //167 / 121 = 1
    16'b10100111_01111010 : OUT <= 1;  //167 / 122 = 1
    16'b10100111_01111011 : OUT <= 1;  //167 / 123 = 1
    16'b10100111_01111100 : OUT <= 1;  //167 / 124 = 1
    16'b10100111_01111101 : OUT <= 1;  //167 / 125 = 1
    16'b10100111_01111110 : OUT <= 1;  //167 / 126 = 1
    16'b10100111_01111111 : OUT <= 1;  //167 / 127 = 1
    16'b10100111_10000000 : OUT <= 1;  //167 / 128 = 1
    16'b10100111_10000001 : OUT <= 1;  //167 / 129 = 1
    16'b10100111_10000010 : OUT <= 1;  //167 / 130 = 1
    16'b10100111_10000011 : OUT <= 1;  //167 / 131 = 1
    16'b10100111_10000100 : OUT <= 1;  //167 / 132 = 1
    16'b10100111_10000101 : OUT <= 1;  //167 / 133 = 1
    16'b10100111_10000110 : OUT <= 1;  //167 / 134 = 1
    16'b10100111_10000111 : OUT <= 1;  //167 / 135 = 1
    16'b10100111_10001000 : OUT <= 1;  //167 / 136 = 1
    16'b10100111_10001001 : OUT <= 1;  //167 / 137 = 1
    16'b10100111_10001010 : OUT <= 1;  //167 / 138 = 1
    16'b10100111_10001011 : OUT <= 1;  //167 / 139 = 1
    16'b10100111_10001100 : OUT <= 1;  //167 / 140 = 1
    16'b10100111_10001101 : OUT <= 1;  //167 / 141 = 1
    16'b10100111_10001110 : OUT <= 1;  //167 / 142 = 1
    16'b10100111_10001111 : OUT <= 1;  //167 / 143 = 1
    16'b10100111_10010000 : OUT <= 1;  //167 / 144 = 1
    16'b10100111_10010001 : OUT <= 1;  //167 / 145 = 1
    16'b10100111_10010010 : OUT <= 1;  //167 / 146 = 1
    16'b10100111_10010011 : OUT <= 1;  //167 / 147 = 1
    16'b10100111_10010100 : OUT <= 1;  //167 / 148 = 1
    16'b10100111_10010101 : OUT <= 1;  //167 / 149 = 1
    16'b10100111_10010110 : OUT <= 1;  //167 / 150 = 1
    16'b10100111_10010111 : OUT <= 1;  //167 / 151 = 1
    16'b10100111_10011000 : OUT <= 1;  //167 / 152 = 1
    16'b10100111_10011001 : OUT <= 1;  //167 / 153 = 1
    16'b10100111_10011010 : OUT <= 1;  //167 / 154 = 1
    16'b10100111_10011011 : OUT <= 1;  //167 / 155 = 1
    16'b10100111_10011100 : OUT <= 1;  //167 / 156 = 1
    16'b10100111_10011101 : OUT <= 1;  //167 / 157 = 1
    16'b10100111_10011110 : OUT <= 1;  //167 / 158 = 1
    16'b10100111_10011111 : OUT <= 1;  //167 / 159 = 1
    16'b10100111_10100000 : OUT <= 1;  //167 / 160 = 1
    16'b10100111_10100001 : OUT <= 1;  //167 / 161 = 1
    16'b10100111_10100010 : OUT <= 1;  //167 / 162 = 1
    16'b10100111_10100011 : OUT <= 1;  //167 / 163 = 1
    16'b10100111_10100100 : OUT <= 1;  //167 / 164 = 1
    16'b10100111_10100101 : OUT <= 1;  //167 / 165 = 1
    16'b10100111_10100110 : OUT <= 1;  //167 / 166 = 1
    16'b10100111_10100111 : OUT <= 1;  //167 / 167 = 1
    16'b10100111_10101000 : OUT <= 0;  //167 / 168 = 0
    16'b10100111_10101001 : OUT <= 0;  //167 / 169 = 0
    16'b10100111_10101010 : OUT <= 0;  //167 / 170 = 0
    16'b10100111_10101011 : OUT <= 0;  //167 / 171 = 0
    16'b10100111_10101100 : OUT <= 0;  //167 / 172 = 0
    16'b10100111_10101101 : OUT <= 0;  //167 / 173 = 0
    16'b10100111_10101110 : OUT <= 0;  //167 / 174 = 0
    16'b10100111_10101111 : OUT <= 0;  //167 / 175 = 0
    16'b10100111_10110000 : OUT <= 0;  //167 / 176 = 0
    16'b10100111_10110001 : OUT <= 0;  //167 / 177 = 0
    16'b10100111_10110010 : OUT <= 0;  //167 / 178 = 0
    16'b10100111_10110011 : OUT <= 0;  //167 / 179 = 0
    16'b10100111_10110100 : OUT <= 0;  //167 / 180 = 0
    16'b10100111_10110101 : OUT <= 0;  //167 / 181 = 0
    16'b10100111_10110110 : OUT <= 0;  //167 / 182 = 0
    16'b10100111_10110111 : OUT <= 0;  //167 / 183 = 0
    16'b10100111_10111000 : OUT <= 0;  //167 / 184 = 0
    16'b10100111_10111001 : OUT <= 0;  //167 / 185 = 0
    16'b10100111_10111010 : OUT <= 0;  //167 / 186 = 0
    16'b10100111_10111011 : OUT <= 0;  //167 / 187 = 0
    16'b10100111_10111100 : OUT <= 0;  //167 / 188 = 0
    16'b10100111_10111101 : OUT <= 0;  //167 / 189 = 0
    16'b10100111_10111110 : OUT <= 0;  //167 / 190 = 0
    16'b10100111_10111111 : OUT <= 0;  //167 / 191 = 0
    16'b10100111_11000000 : OUT <= 0;  //167 / 192 = 0
    16'b10100111_11000001 : OUT <= 0;  //167 / 193 = 0
    16'b10100111_11000010 : OUT <= 0;  //167 / 194 = 0
    16'b10100111_11000011 : OUT <= 0;  //167 / 195 = 0
    16'b10100111_11000100 : OUT <= 0;  //167 / 196 = 0
    16'b10100111_11000101 : OUT <= 0;  //167 / 197 = 0
    16'b10100111_11000110 : OUT <= 0;  //167 / 198 = 0
    16'b10100111_11000111 : OUT <= 0;  //167 / 199 = 0
    16'b10100111_11001000 : OUT <= 0;  //167 / 200 = 0
    16'b10100111_11001001 : OUT <= 0;  //167 / 201 = 0
    16'b10100111_11001010 : OUT <= 0;  //167 / 202 = 0
    16'b10100111_11001011 : OUT <= 0;  //167 / 203 = 0
    16'b10100111_11001100 : OUT <= 0;  //167 / 204 = 0
    16'b10100111_11001101 : OUT <= 0;  //167 / 205 = 0
    16'b10100111_11001110 : OUT <= 0;  //167 / 206 = 0
    16'b10100111_11001111 : OUT <= 0;  //167 / 207 = 0
    16'b10100111_11010000 : OUT <= 0;  //167 / 208 = 0
    16'b10100111_11010001 : OUT <= 0;  //167 / 209 = 0
    16'b10100111_11010010 : OUT <= 0;  //167 / 210 = 0
    16'b10100111_11010011 : OUT <= 0;  //167 / 211 = 0
    16'b10100111_11010100 : OUT <= 0;  //167 / 212 = 0
    16'b10100111_11010101 : OUT <= 0;  //167 / 213 = 0
    16'b10100111_11010110 : OUT <= 0;  //167 / 214 = 0
    16'b10100111_11010111 : OUT <= 0;  //167 / 215 = 0
    16'b10100111_11011000 : OUT <= 0;  //167 / 216 = 0
    16'b10100111_11011001 : OUT <= 0;  //167 / 217 = 0
    16'b10100111_11011010 : OUT <= 0;  //167 / 218 = 0
    16'b10100111_11011011 : OUT <= 0;  //167 / 219 = 0
    16'b10100111_11011100 : OUT <= 0;  //167 / 220 = 0
    16'b10100111_11011101 : OUT <= 0;  //167 / 221 = 0
    16'b10100111_11011110 : OUT <= 0;  //167 / 222 = 0
    16'b10100111_11011111 : OUT <= 0;  //167 / 223 = 0
    16'b10100111_11100000 : OUT <= 0;  //167 / 224 = 0
    16'b10100111_11100001 : OUT <= 0;  //167 / 225 = 0
    16'b10100111_11100010 : OUT <= 0;  //167 / 226 = 0
    16'b10100111_11100011 : OUT <= 0;  //167 / 227 = 0
    16'b10100111_11100100 : OUT <= 0;  //167 / 228 = 0
    16'b10100111_11100101 : OUT <= 0;  //167 / 229 = 0
    16'b10100111_11100110 : OUT <= 0;  //167 / 230 = 0
    16'b10100111_11100111 : OUT <= 0;  //167 / 231 = 0
    16'b10100111_11101000 : OUT <= 0;  //167 / 232 = 0
    16'b10100111_11101001 : OUT <= 0;  //167 / 233 = 0
    16'b10100111_11101010 : OUT <= 0;  //167 / 234 = 0
    16'b10100111_11101011 : OUT <= 0;  //167 / 235 = 0
    16'b10100111_11101100 : OUT <= 0;  //167 / 236 = 0
    16'b10100111_11101101 : OUT <= 0;  //167 / 237 = 0
    16'b10100111_11101110 : OUT <= 0;  //167 / 238 = 0
    16'b10100111_11101111 : OUT <= 0;  //167 / 239 = 0
    16'b10100111_11110000 : OUT <= 0;  //167 / 240 = 0
    16'b10100111_11110001 : OUT <= 0;  //167 / 241 = 0
    16'b10100111_11110010 : OUT <= 0;  //167 / 242 = 0
    16'b10100111_11110011 : OUT <= 0;  //167 / 243 = 0
    16'b10100111_11110100 : OUT <= 0;  //167 / 244 = 0
    16'b10100111_11110101 : OUT <= 0;  //167 / 245 = 0
    16'b10100111_11110110 : OUT <= 0;  //167 / 246 = 0
    16'b10100111_11110111 : OUT <= 0;  //167 / 247 = 0
    16'b10100111_11111000 : OUT <= 0;  //167 / 248 = 0
    16'b10100111_11111001 : OUT <= 0;  //167 / 249 = 0
    16'b10100111_11111010 : OUT <= 0;  //167 / 250 = 0
    16'b10100111_11111011 : OUT <= 0;  //167 / 251 = 0
    16'b10100111_11111100 : OUT <= 0;  //167 / 252 = 0
    16'b10100111_11111101 : OUT <= 0;  //167 / 253 = 0
    16'b10100111_11111110 : OUT <= 0;  //167 / 254 = 0
    16'b10100111_11111111 : OUT <= 0;  //167 / 255 = 0
    16'b10101000_00000000 : OUT <= 0;  //168 / 0 = 0
    16'b10101000_00000001 : OUT <= 168;  //168 / 1 = 168
    16'b10101000_00000010 : OUT <= 84;  //168 / 2 = 84
    16'b10101000_00000011 : OUT <= 56;  //168 / 3 = 56
    16'b10101000_00000100 : OUT <= 42;  //168 / 4 = 42
    16'b10101000_00000101 : OUT <= 33;  //168 / 5 = 33
    16'b10101000_00000110 : OUT <= 28;  //168 / 6 = 28
    16'b10101000_00000111 : OUT <= 24;  //168 / 7 = 24
    16'b10101000_00001000 : OUT <= 21;  //168 / 8 = 21
    16'b10101000_00001001 : OUT <= 18;  //168 / 9 = 18
    16'b10101000_00001010 : OUT <= 16;  //168 / 10 = 16
    16'b10101000_00001011 : OUT <= 15;  //168 / 11 = 15
    16'b10101000_00001100 : OUT <= 14;  //168 / 12 = 14
    16'b10101000_00001101 : OUT <= 12;  //168 / 13 = 12
    16'b10101000_00001110 : OUT <= 12;  //168 / 14 = 12
    16'b10101000_00001111 : OUT <= 11;  //168 / 15 = 11
    16'b10101000_00010000 : OUT <= 10;  //168 / 16 = 10
    16'b10101000_00010001 : OUT <= 9;  //168 / 17 = 9
    16'b10101000_00010010 : OUT <= 9;  //168 / 18 = 9
    16'b10101000_00010011 : OUT <= 8;  //168 / 19 = 8
    16'b10101000_00010100 : OUT <= 8;  //168 / 20 = 8
    16'b10101000_00010101 : OUT <= 8;  //168 / 21 = 8
    16'b10101000_00010110 : OUT <= 7;  //168 / 22 = 7
    16'b10101000_00010111 : OUT <= 7;  //168 / 23 = 7
    16'b10101000_00011000 : OUT <= 7;  //168 / 24 = 7
    16'b10101000_00011001 : OUT <= 6;  //168 / 25 = 6
    16'b10101000_00011010 : OUT <= 6;  //168 / 26 = 6
    16'b10101000_00011011 : OUT <= 6;  //168 / 27 = 6
    16'b10101000_00011100 : OUT <= 6;  //168 / 28 = 6
    16'b10101000_00011101 : OUT <= 5;  //168 / 29 = 5
    16'b10101000_00011110 : OUT <= 5;  //168 / 30 = 5
    16'b10101000_00011111 : OUT <= 5;  //168 / 31 = 5
    16'b10101000_00100000 : OUT <= 5;  //168 / 32 = 5
    16'b10101000_00100001 : OUT <= 5;  //168 / 33 = 5
    16'b10101000_00100010 : OUT <= 4;  //168 / 34 = 4
    16'b10101000_00100011 : OUT <= 4;  //168 / 35 = 4
    16'b10101000_00100100 : OUT <= 4;  //168 / 36 = 4
    16'b10101000_00100101 : OUT <= 4;  //168 / 37 = 4
    16'b10101000_00100110 : OUT <= 4;  //168 / 38 = 4
    16'b10101000_00100111 : OUT <= 4;  //168 / 39 = 4
    16'b10101000_00101000 : OUT <= 4;  //168 / 40 = 4
    16'b10101000_00101001 : OUT <= 4;  //168 / 41 = 4
    16'b10101000_00101010 : OUT <= 4;  //168 / 42 = 4
    16'b10101000_00101011 : OUT <= 3;  //168 / 43 = 3
    16'b10101000_00101100 : OUT <= 3;  //168 / 44 = 3
    16'b10101000_00101101 : OUT <= 3;  //168 / 45 = 3
    16'b10101000_00101110 : OUT <= 3;  //168 / 46 = 3
    16'b10101000_00101111 : OUT <= 3;  //168 / 47 = 3
    16'b10101000_00110000 : OUT <= 3;  //168 / 48 = 3
    16'b10101000_00110001 : OUT <= 3;  //168 / 49 = 3
    16'b10101000_00110010 : OUT <= 3;  //168 / 50 = 3
    16'b10101000_00110011 : OUT <= 3;  //168 / 51 = 3
    16'b10101000_00110100 : OUT <= 3;  //168 / 52 = 3
    16'b10101000_00110101 : OUT <= 3;  //168 / 53 = 3
    16'b10101000_00110110 : OUT <= 3;  //168 / 54 = 3
    16'b10101000_00110111 : OUT <= 3;  //168 / 55 = 3
    16'b10101000_00111000 : OUT <= 3;  //168 / 56 = 3
    16'b10101000_00111001 : OUT <= 2;  //168 / 57 = 2
    16'b10101000_00111010 : OUT <= 2;  //168 / 58 = 2
    16'b10101000_00111011 : OUT <= 2;  //168 / 59 = 2
    16'b10101000_00111100 : OUT <= 2;  //168 / 60 = 2
    16'b10101000_00111101 : OUT <= 2;  //168 / 61 = 2
    16'b10101000_00111110 : OUT <= 2;  //168 / 62 = 2
    16'b10101000_00111111 : OUT <= 2;  //168 / 63 = 2
    16'b10101000_01000000 : OUT <= 2;  //168 / 64 = 2
    16'b10101000_01000001 : OUT <= 2;  //168 / 65 = 2
    16'b10101000_01000010 : OUT <= 2;  //168 / 66 = 2
    16'b10101000_01000011 : OUT <= 2;  //168 / 67 = 2
    16'b10101000_01000100 : OUT <= 2;  //168 / 68 = 2
    16'b10101000_01000101 : OUT <= 2;  //168 / 69 = 2
    16'b10101000_01000110 : OUT <= 2;  //168 / 70 = 2
    16'b10101000_01000111 : OUT <= 2;  //168 / 71 = 2
    16'b10101000_01001000 : OUT <= 2;  //168 / 72 = 2
    16'b10101000_01001001 : OUT <= 2;  //168 / 73 = 2
    16'b10101000_01001010 : OUT <= 2;  //168 / 74 = 2
    16'b10101000_01001011 : OUT <= 2;  //168 / 75 = 2
    16'b10101000_01001100 : OUT <= 2;  //168 / 76 = 2
    16'b10101000_01001101 : OUT <= 2;  //168 / 77 = 2
    16'b10101000_01001110 : OUT <= 2;  //168 / 78 = 2
    16'b10101000_01001111 : OUT <= 2;  //168 / 79 = 2
    16'b10101000_01010000 : OUT <= 2;  //168 / 80 = 2
    16'b10101000_01010001 : OUT <= 2;  //168 / 81 = 2
    16'b10101000_01010010 : OUT <= 2;  //168 / 82 = 2
    16'b10101000_01010011 : OUT <= 2;  //168 / 83 = 2
    16'b10101000_01010100 : OUT <= 2;  //168 / 84 = 2
    16'b10101000_01010101 : OUT <= 1;  //168 / 85 = 1
    16'b10101000_01010110 : OUT <= 1;  //168 / 86 = 1
    16'b10101000_01010111 : OUT <= 1;  //168 / 87 = 1
    16'b10101000_01011000 : OUT <= 1;  //168 / 88 = 1
    16'b10101000_01011001 : OUT <= 1;  //168 / 89 = 1
    16'b10101000_01011010 : OUT <= 1;  //168 / 90 = 1
    16'b10101000_01011011 : OUT <= 1;  //168 / 91 = 1
    16'b10101000_01011100 : OUT <= 1;  //168 / 92 = 1
    16'b10101000_01011101 : OUT <= 1;  //168 / 93 = 1
    16'b10101000_01011110 : OUT <= 1;  //168 / 94 = 1
    16'b10101000_01011111 : OUT <= 1;  //168 / 95 = 1
    16'b10101000_01100000 : OUT <= 1;  //168 / 96 = 1
    16'b10101000_01100001 : OUT <= 1;  //168 / 97 = 1
    16'b10101000_01100010 : OUT <= 1;  //168 / 98 = 1
    16'b10101000_01100011 : OUT <= 1;  //168 / 99 = 1
    16'b10101000_01100100 : OUT <= 1;  //168 / 100 = 1
    16'b10101000_01100101 : OUT <= 1;  //168 / 101 = 1
    16'b10101000_01100110 : OUT <= 1;  //168 / 102 = 1
    16'b10101000_01100111 : OUT <= 1;  //168 / 103 = 1
    16'b10101000_01101000 : OUT <= 1;  //168 / 104 = 1
    16'b10101000_01101001 : OUT <= 1;  //168 / 105 = 1
    16'b10101000_01101010 : OUT <= 1;  //168 / 106 = 1
    16'b10101000_01101011 : OUT <= 1;  //168 / 107 = 1
    16'b10101000_01101100 : OUT <= 1;  //168 / 108 = 1
    16'b10101000_01101101 : OUT <= 1;  //168 / 109 = 1
    16'b10101000_01101110 : OUT <= 1;  //168 / 110 = 1
    16'b10101000_01101111 : OUT <= 1;  //168 / 111 = 1
    16'b10101000_01110000 : OUT <= 1;  //168 / 112 = 1
    16'b10101000_01110001 : OUT <= 1;  //168 / 113 = 1
    16'b10101000_01110010 : OUT <= 1;  //168 / 114 = 1
    16'b10101000_01110011 : OUT <= 1;  //168 / 115 = 1
    16'b10101000_01110100 : OUT <= 1;  //168 / 116 = 1
    16'b10101000_01110101 : OUT <= 1;  //168 / 117 = 1
    16'b10101000_01110110 : OUT <= 1;  //168 / 118 = 1
    16'b10101000_01110111 : OUT <= 1;  //168 / 119 = 1
    16'b10101000_01111000 : OUT <= 1;  //168 / 120 = 1
    16'b10101000_01111001 : OUT <= 1;  //168 / 121 = 1
    16'b10101000_01111010 : OUT <= 1;  //168 / 122 = 1
    16'b10101000_01111011 : OUT <= 1;  //168 / 123 = 1
    16'b10101000_01111100 : OUT <= 1;  //168 / 124 = 1
    16'b10101000_01111101 : OUT <= 1;  //168 / 125 = 1
    16'b10101000_01111110 : OUT <= 1;  //168 / 126 = 1
    16'b10101000_01111111 : OUT <= 1;  //168 / 127 = 1
    16'b10101000_10000000 : OUT <= 1;  //168 / 128 = 1
    16'b10101000_10000001 : OUT <= 1;  //168 / 129 = 1
    16'b10101000_10000010 : OUT <= 1;  //168 / 130 = 1
    16'b10101000_10000011 : OUT <= 1;  //168 / 131 = 1
    16'b10101000_10000100 : OUT <= 1;  //168 / 132 = 1
    16'b10101000_10000101 : OUT <= 1;  //168 / 133 = 1
    16'b10101000_10000110 : OUT <= 1;  //168 / 134 = 1
    16'b10101000_10000111 : OUT <= 1;  //168 / 135 = 1
    16'b10101000_10001000 : OUT <= 1;  //168 / 136 = 1
    16'b10101000_10001001 : OUT <= 1;  //168 / 137 = 1
    16'b10101000_10001010 : OUT <= 1;  //168 / 138 = 1
    16'b10101000_10001011 : OUT <= 1;  //168 / 139 = 1
    16'b10101000_10001100 : OUT <= 1;  //168 / 140 = 1
    16'b10101000_10001101 : OUT <= 1;  //168 / 141 = 1
    16'b10101000_10001110 : OUT <= 1;  //168 / 142 = 1
    16'b10101000_10001111 : OUT <= 1;  //168 / 143 = 1
    16'b10101000_10010000 : OUT <= 1;  //168 / 144 = 1
    16'b10101000_10010001 : OUT <= 1;  //168 / 145 = 1
    16'b10101000_10010010 : OUT <= 1;  //168 / 146 = 1
    16'b10101000_10010011 : OUT <= 1;  //168 / 147 = 1
    16'b10101000_10010100 : OUT <= 1;  //168 / 148 = 1
    16'b10101000_10010101 : OUT <= 1;  //168 / 149 = 1
    16'b10101000_10010110 : OUT <= 1;  //168 / 150 = 1
    16'b10101000_10010111 : OUT <= 1;  //168 / 151 = 1
    16'b10101000_10011000 : OUT <= 1;  //168 / 152 = 1
    16'b10101000_10011001 : OUT <= 1;  //168 / 153 = 1
    16'b10101000_10011010 : OUT <= 1;  //168 / 154 = 1
    16'b10101000_10011011 : OUT <= 1;  //168 / 155 = 1
    16'b10101000_10011100 : OUT <= 1;  //168 / 156 = 1
    16'b10101000_10011101 : OUT <= 1;  //168 / 157 = 1
    16'b10101000_10011110 : OUT <= 1;  //168 / 158 = 1
    16'b10101000_10011111 : OUT <= 1;  //168 / 159 = 1
    16'b10101000_10100000 : OUT <= 1;  //168 / 160 = 1
    16'b10101000_10100001 : OUT <= 1;  //168 / 161 = 1
    16'b10101000_10100010 : OUT <= 1;  //168 / 162 = 1
    16'b10101000_10100011 : OUT <= 1;  //168 / 163 = 1
    16'b10101000_10100100 : OUT <= 1;  //168 / 164 = 1
    16'b10101000_10100101 : OUT <= 1;  //168 / 165 = 1
    16'b10101000_10100110 : OUT <= 1;  //168 / 166 = 1
    16'b10101000_10100111 : OUT <= 1;  //168 / 167 = 1
    16'b10101000_10101000 : OUT <= 1;  //168 / 168 = 1
    16'b10101000_10101001 : OUT <= 0;  //168 / 169 = 0
    16'b10101000_10101010 : OUT <= 0;  //168 / 170 = 0
    16'b10101000_10101011 : OUT <= 0;  //168 / 171 = 0
    16'b10101000_10101100 : OUT <= 0;  //168 / 172 = 0
    16'b10101000_10101101 : OUT <= 0;  //168 / 173 = 0
    16'b10101000_10101110 : OUT <= 0;  //168 / 174 = 0
    16'b10101000_10101111 : OUT <= 0;  //168 / 175 = 0
    16'b10101000_10110000 : OUT <= 0;  //168 / 176 = 0
    16'b10101000_10110001 : OUT <= 0;  //168 / 177 = 0
    16'b10101000_10110010 : OUT <= 0;  //168 / 178 = 0
    16'b10101000_10110011 : OUT <= 0;  //168 / 179 = 0
    16'b10101000_10110100 : OUT <= 0;  //168 / 180 = 0
    16'b10101000_10110101 : OUT <= 0;  //168 / 181 = 0
    16'b10101000_10110110 : OUT <= 0;  //168 / 182 = 0
    16'b10101000_10110111 : OUT <= 0;  //168 / 183 = 0
    16'b10101000_10111000 : OUT <= 0;  //168 / 184 = 0
    16'b10101000_10111001 : OUT <= 0;  //168 / 185 = 0
    16'b10101000_10111010 : OUT <= 0;  //168 / 186 = 0
    16'b10101000_10111011 : OUT <= 0;  //168 / 187 = 0
    16'b10101000_10111100 : OUT <= 0;  //168 / 188 = 0
    16'b10101000_10111101 : OUT <= 0;  //168 / 189 = 0
    16'b10101000_10111110 : OUT <= 0;  //168 / 190 = 0
    16'b10101000_10111111 : OUT <= 0;  //168 / 191 = 0
    16'b10101000_11000000 : OUT <= 0;  //168 / 192 = 0
    16'b10101000_11000001 : OUT <= 0;  //168 / 193 = 0
    16'b10101000_11000010 : OUT <= 0;  //168 / 194 = 0
    16'b10101000_11000011 : OUT <= 0;  //168 / 195 = 0
    16'b10101000_11000100 : OUT <= 0;  //168 / 196 = 0
    16'b10101000_11000101 : OUT <= 0;  //168 / 197 = 0
    16'b10101000_11000110 : OUT <= 0;  //168 / 198 = 0
    16'b10101000_11000111 : OUT <= 0;  //168 / 199 = 0
    16'b10101000_11001000 : OUT <= 0;  //168 / 200 = 0
    16'b10101000_11001001 : OUT <= 0;  //168 / 201 = 0
    16'b10101000_11001010 : OUT <= 0;  //168 / 202 = 0
    16'b10101000_11001011 : OUT <= 0;  //168 / 203 = 0
    16'b10101000_11001100 : OUT <= 0;  //168 / 204 = 0
    16'b10101000_11001101 : OUT <= 0;  //168 / 205 = 0
    16'b10101000_11001110 : OUT <= 0;  //168 / 206 = 0
    16'b10101000_11001111 : OUT <= 0;  //168 / 207 = 0
    16'b10101000_11010000 : OUT <= 0;  //168 / 208 = 0
    16'b10101000_11010001 : OUT <= 0;  //168 / 209 = 0
    16'b10101000_11010010 : OUT <= 0;  //168 / 210 = 0
    16'b10101000_11010011 : OUT <= 0;  //168 / 211 = 0
    16'b10101000_11010100 : OUT <= 0;  //168 / 212 = 0
    16'b10101000_11010101 : OUT <= 0;  //168 / 213 = 0
    16'b10101000_11010110 : OUT <= 0;  //168 / 214 = 0
    16'b10101000_11010111 : OUT <= 0;  //168 / 215 = 0
    16'b10101000_11011000 : OUT <= 0;  //168 / 216 = 0
    16'b10101000_11011001 : OUT <= 0;  //168 / 217 = 0
    16'b10101000_11011010 : OUT <= 0;  //168 / 218 = 0
    16'b10101000_11011011 : OUT <= 0;  //168 / 219 = 0
    16'b10101000_11011100 : OUT <= 0;  //168 / 220 = 0
    16'b10101000_11011101 : OUT <= 0;  //168 / 221 = 0
    16'b10101000_11011110 : OUT <= 0;  //168 / 222 = 0
    16'b10101000_11011111 : OUT <= 0;  //168 / 223 = 0
    16'b10101000_11100000 : OUT <= 0;  //168 / 224 = 0
    16'b10101000_11100001 : OUT <= 0;  //168 / 225 = 0
    16'b10101000_11100010 : OUT <= 0;  //168 / 226 = 0
    16'b10101000_11100011 : OUT <= 0;  //168 / 227 = 0
    16'b10101000_11100100 : OUT <= 0;  //168 / 228 = 0
    16'b10101000_11100101 : OUT <= 0;  //168 / 229 = 0
    16'b10101000_11100110 : OUT <= 0;  //168 / 230 = 0
    16'b10101000_11100111 : OUT <= 0;  //168 / 231 = 0
    16'b10101000_11101000 : OUT <= 0;  //168 / 232 = 0
    16'b10101000_11101001 : OUT <= 0;  //168 / 233 = 0
    16'b10101000_11101010 : OUT <= 0;  //168 / 234 = 0
    16'b10101000_11101011 : OUT <= 0;  //168 / 235 = 0
    16'b10101000_11101100 : OUT <= 0;  //168 / 236 = 0
    16'b10101000_11101101 : OUT <= 0;  //168 / 237 = 0
    16'b10101000_11101110 : OUT <= 0;  //168 / 238 = 0
    16'b10101000_11101111 : OUT <= 0;  //168 / 239 = 0
    16'b10101000_11110000 : OUT <= 0;  //168 / 240 = 0
    16'b10101000_11110001 : OUT <= 0;  //168 / 241 = 0
    16'b10101000_11110010 : OUT <= 0;  //168 / 242 = 0
    16'b10101000_11110011 : OUT <= 0;  //168 / 243 = 0
    16'b10101000_11110100 : OUT <= 0;  //168 / 244 = 0
    16'b10101000_11110101 : OUT <= 0;  //168 / 245 = 0
    16'b10101000_11110110 : OUT <= 0;  //168 / 246 = 0
    16'b10101000_11110111 : OUT <= 0;  //168 / 247 = 0
    16'b10101000_11111000 : OUT <= 0;  //168 / 248 = 0
    16'b10101000_11111001 : OUT <= 0;  //168 / 249 = 0
    16'b10101000_11111010 : OUT <= 0;  //168 / 250 = 0
    16'b10101000_11111011 : OUT <= 0;  //168 / 251 = 0
    16'b10101000_11111100 : OUT <= 0;  //168 / 252 = 0
    16'b10101000_11111101 : OUT <= 0;  //168 / 253 = 0
    16'b10101000_11111110 : OUT <= 0;  //168 / 254 = 0
    16'b10101000_11111111 : OUT <= 0;  //168 / 255 = 0
    16'b10101001_00000000 : OUT <= 0;  //169 / 0 = 0
    16'b10101001_00000001 : OUT <= 169;  //169 / 1 = 169
    16'b10101001_00000010 : OUT <= 84;  //169 / 2 = 84
    16'b10101001_00000011 : OUT <= 56;  //169 / 3 = 56
    16'b10101001_00000100 : OUT <= 42;  //169 / 4 = 42
    16'b10101001_00000101 : OUT <= 33;  //169 / 5 = 33
    16'b10101001_00000110 : OUT <= 28;  //169 / 6 = 28
    16'b10101001_00000111 : OUT <= 24;  //169 / 7 = 24
    16'b10101001_00001000 : OUT <= 21;  //169 / 8 = 21
    16'b10101001_00001001 : OUT <= 18;  //169 / 9 = 18
    16'b10101001_00001010 : OUT <= 16;  //169 / 10 = 16
    16'b10101001_00001011 : OUT <= 15;  //169 / 11 = 15
    16'b10101001_00001100 : OUT <= 14;  //169 / 12 = 14
    16'b10101001_00001101 : OUT <= 13;  //169 / 13 = 13
    16'b10101001_00001110 : OUT <= 12;  //169 / 14 = 12
    16'b10101001_00001111 : OUT <= 11;  //169 / 15 = 11
    16'b10101001_00010000 : OUT <= 10;  //169 / 16 = 10
    16'b10101001_00010001 : OUT <= 9;  //169 / 17 = 9
    16'b10101001_00010010 : OUT <= 9;  //169 / 18 = 9
    16'b10101001_00010011 : OUT <= 8;  //169 / 19 = 8
    16'b10101001_00010100 : OUT <= 8;  //169 / 20 = 8
    16'b10101001_00010101 : OUT <= 8;  //169 / 21 = 8
    16'b10101001_00010110 : OUT <= 7;  //169 / 22 = 7
    16'b10101001_00010111 : OUT <= 7;  //169 / 23 = 7
    16'b10101001_00011000 : OUT <= 7;  //169 / 24 = 7
    16'b10101001_00011001 : OUT <= 6;  //169 / 25 = 6
    16'b10101001_00011010 : OUT <= 6;  //169 / 26 = 6
    16'b10101001_00011011 : OUT <= 6;  //169 / 27 = 6
    16'b10101001_00011100 : OUT <= 6;  //169 / 28 = 6
    16'b10101001_00011101 : OUT <= 5;  //169 / 29 = 5
    16'b10101001_00011110 : OUT <= 5;  //169 / 30 = 5
    16'b10101001_00011111 : OUT <= 5;  //169 / 31 = 5
    16'b10101001_00100000 : OUT <= 5;  //169 / 32 = 5
    16'b10101001_00100001 : OUT <= 5;  //169 / 33 = 5
    16'b10101001_00100010 : OUT <= 4;  //169 / 34 = 4
    16'b10101001_00100011 : OUT <= 4;  //169 / 35 = 4
    16'b10101001_00100100 : OUT <= 4;  //169 / 36 = 4
    16'b10101001_00100101 : OUT <= 4;  //169 / 37 = 4
    16'b10101001_00100110 : OUT <= 4;  //169 / 38 = 4
    16'b10101001_00100111 : OUT <= 4;  //169 / 39 = 4
    16'b10101001_00101000 : OUT <= 4;  //169 / 40 = 4
    16'b10101001_00101001 : OUT <= 4;  //169 / 41 = 4
    16'b10101001_00101010 : OUT <= 4;  //169 / 42 = 4
    16'b10101001_00101011 : OUT <= 3;  //169 / 43 = 3
    16'b10101001_00101100 : OUT <= 3;  //169 / 44 = 3
    16'b10101001_00101101 : OUT <= 3;  //169 / 45 = 3
    16'b10101001_00101110 : OUT <= 3;  //169 / 46 = 3
    16'b10101001_00101111 : OUT <= 3;  //169 / 47 = 3
    16'b10101001_00110000 : OUT <= 3;  //169 / 48 = 3
    16'b10101001_00110001 : OUT <= 3;  //169 / 49 = 3
    16'b10101001_00110010 : OUT <= 3;  //169 / 50 = 3
    16'b10101001_00110011 : OUT <= 3;  //169 / 51 = 3
    16'b10101001_00110100 : OUT <= 3;  //169 / 52 = 3
    16'b10101001_00110101 : OUT <= 3;  //169 / 53 = 3
    16'b10101001_00110110 : OUT <= 3;  //169 / 54 = 3
    16'b10101001_00110111 : OUT <= 3;  //169 / 55 = 3
    16'b10101001_00111000 : OUT <= 3;  //169 / 56 = 3
    16'b10101001_00111001 : OUT <= 2;  //169 / 57 = 2
    16'b10101001_00111010 : OUT <= 2;  //169 / 58 = 2
    16'b10101001_00111011 : OUT <= 2;  //169 / 59 = 2
    16'b10101001_00111100 : OUT <= 2;  //169 / 60 = 2
    16'b10101001_00111101 : OUT <= 2;  //169 / 61 = 2
    16'b10101001_00111110 : OUT <= 2;  //169 / 62 = 2
    16'b10101001_00111111 : OUT <= 2;  //169 / 63 = 2
    16'b10101001_01000000 : OUT <= 2;  //169 / 64 = 2
    16'b10101001_01000001 : OUT <= 2;  //169 / 65 = 2
    16'b10101001_01000010 : OUT <= 2;  //169 / 66 = 2
    16'b10101001_01000011 : OUT <= 2;  //169 / 67 = 2
    16'b10101001_01000100 : OUT <= 2;  //169 / 68 = 2
    16'b10101001_01000101 : OUT <= 2;  //169 / 69 = 2
    16'b10101001_01000110 : OUT <= 2;  //169 / 70 = 2
    16'b10101001_01000111 : OUT <= 2;  //169 / 71 = 2
    16'b10101001_01001000 : OUT <= 2;  //169 / 72 = 2
    16'b10101001_01001001 : OUT <= 2;  //169 / 73 = 2
    16'b10101001_01001010 : OUT <= 2;  //169 / 74 = 2
    16'b10101001_01001011 : OUT <= 2;  //169 / 75 = 2
    16'b10101001_01001100 : OUT <= 2;  //169 / 76 = 2
    16'b10101001_01001101 : OUT <= 2;  //169 / 77 = 2
    16'b10101001_01001110 : OUT <= 2;  //169 / 78 = 2
    16'b10101001_01001111 : OUT <= 2;  //169 / 79 = 2
    16'b10101001_01010000 : OUT <= 2;  //169 / 80 = 2
    16'b10101001_01010001 : OUT <= 2;  //169 / 81 = 2
    16'b10101001_01010010 : OUT <= 2;  //169 / 82 = 2
    16'b10101001_01010011 : OUT <= 2;  //169 / 83 = 2
    16'b10101001_01010100 : OUT <= 2;  //169 / 84 = 2
    16'b10101001_01010101 : OUT <= 1;  //169 / 85 = 1
    16'b10101001_01010110 : OUT <= 1;  //169 / 86 = 1
    16'b10101001_01010111 : OUT <= 1;  //169 / 87 = 1
    16'b10101001_01011000 : OUT <= 1;  //169 / 88 = 1
    16'b10101001_01011001 : OUT <= 1;  //169 / 89 = 1
    16'b10101001_01011010 : OUT <= 1;  //169 / 90 = 1
    16'b10101001_01011011 : OUT <= 1;  //169 / 91 = 1
    16'b10101001_01011100 : OUT <= 1;  //169 / 92 = 1
    16'b10101001_01011101 : OUT <= 1;  //169 / 93 = 1
    16'b10101001_01011110 : OUT <= 1;  //169 / 94 = 1
    16'b10101001_01011111 : OUT <= 1;  //169 / 95 = 1
    16'b10101001_01100000 : OUT <= 1;  //169 / 96 = 1
    16'b10101001_01100001 : OUT <= 1;  //169 / 97 = 1
    16'b10101001_01100010 : OUT <= 1;  //169 / 98 = 1
    16'b10101001_01100011 : OUT <= 1;  //169 / 99 = 1
    16'b10101001_01100100 : OUT <= 1;  //169 / 100 = 1
    16'b10101001_01100101 : OUT <= 1;  //169 / 101 = 1
    16'b10101001_01100110 : OUT <= 1;  //169 / 102 = 1
    16'b10101001_01100111 : OUT <= 1;  //169 / 103 = 1
    16'b10101001_01101000 : OUT <= 1;  //169 / 104 = 1
    16'b10101001_01101001 : OUT <= 1;  //169 / 105 = 1
    16'b10101001_01101010 : OUT <= 1;  //169 / 106 = 1
    16'b10101001_01101011 : OUT <= 1;  //169 / 107 = 1
    16'b10101001_01101100 : OUT <= 1;  //169 / 108 = 1
    16'b10101001_01101101 : OUT <= 1;  //169 / 109 = 1
    16'b10101001_01101110 : OUT <= 1;  //169 / 110 = 1
    16'b10101001_01101111 : OUT <= 1;  //169 / 111 = 1
    16'b10101001_01110000 : OUT <= 1;  //169 / 112 = 1
    16'b10101001_01110001 : OUT <= 1;  //169 / 113 = 1
    16'b10101001_01110010 : OUT <= 1;  //169 / 114 = 1
    16'b10101001_01110011 : OUT <= 1;  //169 / 115 = 1
    16'b10101001_01110100 : OUT <= 1;  //169 / 116 = 1
    16'b10101001_01110101 : OUT <= 1;  //169 / 117 = 1
    16'b10101001_01110110 : OUT <= 1;  //169 / 118 = 1
    16'b10101001_01110111 : OUT <= 1;  //169 / 119 = 1
    16'b10101001_01111000 : OUT <= 1;  //169 / 120 = 1
    16'b10101001_01111001 : OUT <= 1;  //169 / 121 = 1
    16'b10101001_01111010 : OUT <= 1;  //169 / 122 = 1
    16'b10101001_01111011 : OUT <= 1;  //169 / 123 = 1
    16'b10101001_01111100 : OUT <= 1;  //169 / 124 = 1
    16'b10101001_01111101 : OUT <= 1;  //169 / 125 = 1
    16'b10101001_01111110 : OUT <= 1;  //169 / 126 = 1
    16'b10101001_01111111 : OUT <= 1;  //169 / 127 = 1
    16'b10101001_10000000 : OUT <= 1;  //169 / 128 = 1
    16'b10101001_10000001 : OUT <= 1;  //169 / 129 = 1
    16'b10101001_10000010 : OUT <= 1;  //169 / 130 = 1
    16'b10101001_10000011 : OUT <= 1;  //169 / 131 = 1
    16'b10101001_10000100 : OUT <= 1;  //169 / 132 = 1
    16'b10101001_10000101 : OUT <= 1;  //169 / 133 = 1
    16'b10101001_10000110 : OUT <= 1;  //169 / 134 = 1
    16'b10101001_10000111 : OUT <= 1;  //169 / 135 = 1
    16'b10101001_10001000 : OUT <= 1;  //169 / 136 = 1
    16'b10101001_10001001 : OUT <= 1;  //169 / 137 = 1
    16'b10101001_10001010 : OUT <= 1;  //169 / 138 = 1
    16'b10101001_10001011 : OUT <= 1;  //169 / 139 = 1
    16'b10101001_10001100 : OUT <= 1;  //169 / 140 = 1
    16'b10101001_10001101 : OUT <= 1;  //169 / 141 = 1
    16'b10101001_10001110 : OUT <= 1;  //169 / 142 = 1
    16'b10101001_10001111 : OUT <= 1;  //169 / 143 = 1
    16'b10101001_10010000 : OUT <= 1;  //169 / 144 = 1
    16'b10101001_10010001 : OUT <= 1;  //169 / 145 = 1
    16'b10101001_10010010 : OUT <= 1;  //169 / 146 = 1
    16'b10101001_10010011 : OUT <= 1;  //169 / 147 = 1
    16'b10101001_10010100 : OUT <= 1;  //169 / 148 = 1
    16'b10101001_10010101 : OUT <= 1;  //169 / 149 = 1
    16'b10101001_10010110 : OUT <= 1;  //169 / 150 = 1
    16'b10101001_10010111 : OUT <= 1;  //169 / 151 = 1
    16'b10101001_10011000 : OUT <= 1;  //169 / 152 = 1
    16'b10101001_10011001 : OUT <= 1;  //169 / 153 = 1
    16'b10101001_10011010 : OUT <= 1;  //169 / 154 = 1
    16'b10101001_10011011 : OUT <= 1;  //169 / 155 = 1
    16'b10101001_10011100 : OUT <= 1;  //169 / 156 = 1
    16'b10101001_10011101 : OUT <= 1;  //169 / 157 = 1
    16'b10101001_10011110 : OUT <= 1;  //169 / 158 = 1
    16'b10101001_10011111 : OUT <= 1;  //169 / 159 = 1
    16'b10101001_10100000 : OUT <= 1;  //169 / 160 = 1
    16'b10101001_10100001 : OUT <= 1;  //169 / 161 = 1
    16'b10101001_10100010 : OUT <= 1;  //169 / 162 = 1
    16'b10101001_10100011 : OUT <= 1;  //169 / 163 = 1
    16'b10101001_10100100 : OUT <= 1;  //169 / 164 = 1
    16'b10101001_10100101 : OUT <= 1;  //169 / 165 = 1
    16'b10101001_10100110 : OUT <= 1;  //169 / 166 = 1
    16'b10101001_10100111 : OUT <= 1;  //169 / 167 = 1
    16'b10101001_10101000 : OUT <= 1;  //169 / 168 = 1
    16'b10101001_10101001 : OUT <= 1;  //169 / 169 = 1
    16'b10101001_10101010 : OUT <= 0;  //169 / 170 = 0
    16'b10101001_10101011 : OUT <= 0;  //169 / 171 = 0
    16'b10101001_10101100 : OUT <= 0;  //169 / 172 = 0
    16'b10101001_10101101 : OUT <= 0;  //169 / 173 = 0
    16'b10101001_10101110 : OUT <= 0;  //169 / 174 = 0
    16'b10101001_10101111 : OUT <= 0;  //169 / 175 = 0
    16'b10101001_10110000 : OUT <= 0;  //169 / 176 = 0
    16'b10101001_10110001 : OUT <= 0;  //169 / 177 = 0
    16'b10101001_10110010 : OUT <= 0;  //169 / 178 = 0
    16'b10101001_10110011 : OUT <= 0;  //169 / 179 = 0
    16'b10101001_10110100 : OUT <= 0;  //169 / 180 = 0
    16'b10101001_10110101 : OUT <= 0;  //169 / 181 = 0
    16'b10101001_10110110 : OUT <= 0;  //169 / 182 = 0
    16'b10101001_10110111 : OUT <= 0;  //169 / 183 = 0
    16'b10101001_10111000 : OUT <= 0;  //169 / 184 = 0
    16'b10101001_10111001 : OUT <= 0;  //169 / 185 = 0
    16'b10101001_10111010 : OUT <= 0;  //169 / 186 = 0
    16'b10101001_10111011 : OUT <= 0;  //169 / 187 = 0
    16'b10101001_10111100 : OUT <= 0;  //169 / 188 = 0
    16'b10101001_10111101 : OUT <= 0;  //169 / 189 = 0
    16'b10101001_10111110 : OUT <= 0;  //169 / 190 = 0
    16'b10101001_10111111 : OUT <= 0;  //169 / 191 = 0
    16'b10101001_11000000 : OUT <= 0;  //169 / 192 = 0
    16'b10101001_11000001 : OUT <= 0;  //169 / 193 = 0
    16'b10101001_11000010 : OUT <= 0;  //169 / 194 = 0
    16'b10101001_11000011 : OUT <= 0;  //169 / 195 = 0
    16'b10101001_11000100 : OUT <= 0;  //169 / 196 = 0
    16'b10101001_11000101 : OUT <= 0;  //169 / 197 = 0
    16'b10101001_11000110 : OUT <= 0;  //169 / 198 = 0
    16'b10101001_11000111 : OUT <= 0;  //169 / 199 = 0
    16'b10101001_11001000 : OUT <= 0;  //169 / 200 = 0
    16'b10101001_11001001 : OUT <= 0;  //169 / 201 = 0
    16'b10101001_11001010 : OUT <= 0;  //169 / 202 = 0
    16'b10101001_11001011 : OUT <= 0;  //169 / 203 = 0
    16'b10101001_11001100 : OUT <= 0;  //169 / 204 = 0
    16'b10101001_11001101 : OUT <= 0;  //169 / 205 = 0
    16'b10101001_11001110 : OUT <= 0;  //169 / 206 = 0
    16'b10101001_11001111 : OUT <= 0;  //169 / 207 = 0
    16'b10101001_11010000 : OUT <= 0;  //169 / 208 = 0
    16'b10101001_11010001 : OUT <= 0;  //169 / 209 = 0
    16'b10101001_11010010 : OUT <= 0;  //169 / 210 = 0
    16'b10101001_11010011 : OUT <= 0;  //169 / 211 = 0
    16'b10101001_11010100 : OUT <= 0;  //169 / 212 = 0
    16'b10101001_11010101 : OUT <= 0;  //169 / 213 = 0
    16'b10101001_11010110 : OUT <= 0;  //169 / 214 = 0
    16'b10101001_11010111 : OUT <= 0;  //169 / 215 = 0
    16'b10101001_11011000 : OUT <= 0;  //169 / 216 = 0
    16'b10101001_11011001 : OUT <= 0;  //169 / 217 = 0
    16'b10101001_11011010 : OUT <= 0;  //169 / 218 = 0
    16'b10101001_11011011 : OUT <= 0;  //169 / 219 = 0
    16'b10101001_11011100 : OUT <= 0;  //169 / 220 = 0
    16'b10101001_11011101 : OUT <= 0;  //169 / 221 = 0
    16'b10101001_11011110 : OUT <= 0;  //169 / 222 = 0
    16'b10101001_11011111 : OUT <= 0;  //169 / 223 = 0
    16'b10101001_11100000 : OUT <= 0;  //169 / 224 = 0
    16'b10101001_11100001 : OUT <= 0;  //169 / 225 = 0
    16'b10101001_11100010 : OUT <= 0;  //169 / 226 = 0
    16'b10101001_11100011 : OUT <= 0;  //169 / 227 = 0
    16'b10101001_11100100 : OUT <= 0;  //169 / 228 = 0
    16'b10101001_11100101 : OUT <= 0;  //169 / 229 = 0
    16'b10101001_11100110 : OUT <= 0;  //169 / 230 = 0
    16'b10101001_11100111 : OUT <= 0;  //169 / 231 = 0
    16'b10101001_11101000 : OUT <= 0;  //169 / 232 = 0
    16'b10101001_11101001 : OUT <= 0;  //169 / 233 = 0
    16'b10101001_11101010 : OUT <= 0;  //169 / 234 = 0
    16'b10101001_11101011 : OUT <= 0;  //169 / 235 = 0
    16'b10101001_11101100 : OUT <= 0;  //169 / 236 = 0
    16'b10101001_11101101 : OUT <= 0;  //169 / 237 = 0
    16'b10101001_11101110 : OUT <= 0;  //169 / 238 = 0
    16'b10101001_11101111 : OUT <= 0;  //169 / 239 = 0
    16'b10101001_11110000 : OUT <= 0;  //169 / 240 = 0
    16'b10101001_11110001 : OUT <= 0;  //169 / 241 = 0
    16'b10101001_11110010 : OUT <= 0;  //169 / 242 = 0
    16'b10101001_11110011 : OUT <= 0;  //169 / 243 = 0
    16'b10101001_11110100 : OUT <= 0;  //169 / 244 = 0
    16'b10101001_11110101 : OUT <= 0;  //169 / 245 = 0
    16'b10101001_11110110 : OUT <= 0;  //169 / 246 = 0
    16'b10101001_11110111 : OUT <= 0;  //169 / 247 = 0
    16'b10101001_11111000 : OUT <= 0;  //169 / 248 = 0
    16'b10101001_11111001 : OUT <= 0;  //169 / 249 = 0
    16'b10101001_11111010 : OUT <= 0;  //169 / 250 = 0
    16'b10101001_11111011 : OUT <= 0;  //169 / 251 = 0
    16'b10101001_11111100 : OUT <= 0;  //169 / 252 = 0
    16'b10101001_11111101 : OUT <= 0;  //169 / 253 = 0
    16'b10101001_11111110 : OUT <= 0;  //169 / 254 = 0
    16'b10101001_11111111 : OUT <= 0;  //169 / 255 = 0
    16'b10101010_00000000 : OUT <= 0;  //170 / 0 = 0
    16'b10101010_00000001 : OUT <= 170;  //170 / 1 = 170
    16'b10101010_00000010 : OUT <= 85;  //170 / 2 = 85
    16'b10101010_00000011 : OUT <= 56;  //170 / 3 = 56
    16'b10101010_00000100 : OUT <= 42;  //170 / 4 = 42
    16'b10101010_00000101 : OUT <= 34;  //170 / 5 = 34
    16'b10101010_00000110 : OUT <= 28;  //170 / 6 = 28
    16'b10101010_00000111 : OUT <= 24;  //170 / 7 = 24
    16'b10101010_00001000 : OUT <= 21;  //170 / 8 = 21
    16'b10101010_00001001 : OUT <= 18;  //170 / 9 = 18
    16'b10101010_00001010 : OUT <= 17;  //170 / 10 = 17
    16'b10101010_00001011 : OUT <= 15;  //170 / 11 = 15
    16'b10101010_00001100 : OUT <= 14;  //170 / 12 = 14
    16'b10101010_00001101 : OUT <= 13;  //170 / 13 = 13
    16'b10101010_00001110 : OUT <= 12;  //170 / 14 = 12
    16'b10101010_00001111 : OUT <= 11;  //170 / 15 = 11
    16'b10101010_00010000 : OUT <= 10;  //170 / 16 = 10
    16'b10101010_00010001 : OUT <= 10;  //170 / 17 = 10
    16'b10101010_00010010 : OUT <= 9;  //170 / 18 = 9
    16'b10101010_00010011 : OUT <= 8;  //170 / 19 = 8
    16'b10101010_00010100 : OUT <= 8;  //170 / 20 = 8
    16'b10101010_00010101 : OUT <= 8;  //170 / 21 = 8
    16'b10101010_00010110 : OUT <= 7;  //170 / 22 = 7
    16'b10101010_00010111 : OUT <= 7;  //170 / 23 = 7
    16'b10101010_00011000 : OUT <= 7;  //170 / 24 = 7
    16'b10101010_00011001 : OUT <= 6;  //170 / 25 = 6
    16'b10101010_00011010 : OUT <= 6;  //170 / 26 = 6
    16'b10101010_00011011 : OUT <= 6;  //170 / 27 = 6
    16'b10101010_00011100 : OUT <= 6;  //170 / 28 = 6
    16'b10101010_00011101 : OUT <= 5;  //170 / 29 = 5
    16'b10101010_00011110 : OUT <= 5;  //170 / 30 = 5
    16'b10101010_00011111 : OUT <= 5;  //170 / 31 = 5
    16'b10101010_00100000 : OUT <= 5;  //170 / 32 = 5
    16'b10101010_00100001 : OUT <= 5;  //170 / 33 = 5
    16'b10101010_00100010 : OUT <= 5;  //170 / 34 = 5
    16'b10101010_00100011 : OUT <= 4;  //170 / 35 = 4
    16'b10101010_00100100 : OUT <= 4;  //170 / 36 = 4
    16'b10101010_00100101 : OUT <= 4;  //170 / 37 = 4
    16'b10101010_00100110 : OUT <= 4;  //170 / 38 = 4
    16'b10101010_00100111 : OUT <= 4;  //170 / 39 = 4
    16'b10101010_00101000 : OUT <= 4;  //170 / 40 = 4
    16'b10101010_00101001 : OUT <= 4;  //170 / 41 = 4
    16'b10101010_00101010 : OUT <= 4;  //170 / 42 = 4
    16'b10101010_00101011 : OUT <= 3;  //170 / 43 = 3
    16'b10101010_00101100 : OUT <= 3;  //170 / 44 = 3
    16'b10101010_00101101 : OUT <= 3;  //170 / 45 = 3
    16'b10101010_00101110 : OUT <= 3;  //170 / 46 = 3
    16'b10101010_00101111 : OUT <= 3;  //170 / 47 = 3
    16'b10101010_00110000 : OUT <= 3;  //170 / 48 = 3
    16'b10101010_00110001 : OUT <= 3;  //170 / 49 = 3
    16'b10101010_00110010 : OUT <= 3;  //170 / 50 = 3
    16'b10101010_00110011 : OUT <= 3;  //170 / 51 = 3
    16'b10101010_00110100 : OUT <= 3;  //170 / 52 = 3
    16'b10101010_00110101 : OUT <= 3;  //170 / 53 = 3
    16'b10101010_00110110 : OUT <= 3;  //170 / 54 = 3
    16'b10101010_00110111 : OUT <= 3;  //170 / 55 = 3
    16'b10101010_00111000 : OUT <= 3;  //170 / 56 = 3
    16'b10101010_00111001 : OUT <= 2;  //170 / 57 = 2
    16'b10101010_00111010 : OUT <= 2;  //170 / 58 = 2
    16'b10101010_00111011 : OUT <= 2;  //170 / 59 = 2
    16'b10101010_00111100 : OUT <= 2;  //170 / 60 = 2
    16'b10101010_00111101 : OUT <= 2;  //170 / 61 = 2
    16'b10101010_00111110 : OUT <= 2;  //170 / 62 = 2
    16'b10101010_00111111 : OUT <= 2;  //170 / 63 = 2
    16'b10101010_01000000 : OUT <= 2;  //170 / 64 = 2
    16'b10101010_01000001 : OUT <= 2;  //170 / 65 = 2
    16'b10101010_01000010 : OUT <= 2;  //170 / 66 = 2
    16'b10101010_01000011 : OUT <= 2;  //170 / 67 = 2
    16'b10101010_01000100 : OUT <= 2;  //170 / 68 = 2
    16'b10101010_01000101 : OUT <= 2;  //170 / 69 = 2
    16'b10101010_01000110 : OUT <= 2;  //170 / 70 = 2
    16'b10101010_01000111 : OUT <= 2;  //170 / 71 = 2
    16'b10101010_01001000 : OUT <= 2;  //170 / 72 = 2
    16'b10101010_01001001 : OUT <= 2;  //170 / 73 = 2
    16'b10101010_01001010 : OUT <= 2;  //170 / 74 = 2
    16'b10101010_01001011 : OUT <= 2;  //170 / 75 = 2
    16'b10101010_01001100 : OUT <= 2;  //170 / 76 = 2
    16'b10101010_01001101 : OUT <= 2;  //170 / 77 = 2
    16'b10101010_01001110 : OUT <= 2;  //170 / 78 = 2
    16'b10101010_01001111 : OUT <= 2;  //170 / 79 = 2
    16'b10101010_01010000 : OUT <= 2;  //170 / 80 = 2
    16'b10101010_01010001 : OUT <= 2;  //170 / 81 = 2
    16'b10101010_01010010 : OUT <= 2;  //170 / 82 = 2
    16'b10101010_01010011 : OUT <= 2;  //170 / 83 = 2
    16'b10101010_01010100 : OUT <= 2;  //170 / 84 = 2
    16'b10101010_01010101 : OUT <= 2;  //170 / 85 = 2
    16'b10101010_01010110 : OUT <= 1;  //170 / 86 = 1
    16'b10101010_01010111 : OUT <= 1;  //170 / 87 = 1
    16'b10101010_01011000 : OUT <= 1;  //170 / 88 = 1
    16'b10101010_01011001 : OUT <= 1;  //170 / 89 = 1
    16'b10101010_01011010 : OUT <= 1;  //170 / 90 = 1
    16'b10101010_01011011 : OUT <= 1;  //170 / 91 = 1
    16'b10101010_01011100 : OUT <= 1;  //170 / 92 = 1
    16'b10101010_01011101 : OUT <= 1;  //170 / 93 = 1
    16'b10101010_01011110 : OUT <= 1;  //170 / 94 = 1
    16'b10101010_01011111 : OUT <= 1;  //170 / 95 = 1
    16'b10101010_01100000 : OUT <= 1;  //170 / 96 = 1
    16'b10101010_01100001 : OUT <= 1;  //170 / 97 = 1
    16'b10101010_01100010 : OUT <= 1;  //170 / 98 = 1
    16'b10101010_01100011 : OUT <= 1;  //170 / 99 = 1
    16'b10101010_01100100 : OUT <= 1;  //170 / 100 = 1
    16'b10101010_01100101 : OUT <= 1;  //170 / 101 = 1
    16'b10101010_01100110 : OUT <= 1;  //170 / 102 = 1
    16'b10101010_01100111 : OUT <= 1;  //170 / 103 = 1
    16'b10101010_01101000 : OUT <= 1;  //170 / 104 = 1
    16'b10101010_01101001 : OUT <= 1;  //170 / 105 = 1
    16'b10101010_01101010 : OUT <= 1;  //170 / 106 = 1
    16'b10101010_01101011 : OUT <= 1;  //170 / 107 = 1
    16'b10101010_01101100 : OUT <= 1;  //170 / 108 = 1
    16'b10101010_01101101 : OUT <= 1;  //170 / 109 = 1
    16'b10101010_01101110 : OUT <= 1;  //170 / 110 = 1
    16'b10101010_01101111 : OUT <= 1;  //170 / 111 = 1
    16'b10101010_01110000 : OUT <= 1;  //170 / 112 = 1
    16'b10101010_01110001 : OUT <= 1;  //170 / 113 = 1
    16'b10101010_01110010 : OUT <= 1;  //170 / 114 = 1
    16'b10101010_01110011 : OUT <= 1;  //170 / 115 = 1
    16'b10101010_01110100 : OUT <= 1;  //170 / 116 = 1
    16'b10101010_01110101 : OUT <= 1;  //170 / 117 = 1
    16'b10101010_01110110 : OUT <= 1;  //170 / 118 = 1
    16'b10101010_01110111 : OUT <= 1;  //170 / 119 = 1
    16'b10101010_01111000 : OUT <= 1;  //170 / 120 = 1
    16'b10101010_01111001 : OUT <= 1;  //170 / 121 = 1
    16'b10101010_01111010 : OUT <= 1;  //170 / 122 = 1
    16'b10101010_01111011 : OUT <= 1;  //170 / 123 = 1
    16'b10101010_01111100 : OUT <= 1;  //170 / 124 = 1
    16'b10101010_01111101 : OUT <= 1;  //170 / 125 = 1
    16'b10101010_01111110 : OUT <= 1;  //170 / 126 = 1
    16'b10101010_01111111 : OUT <= 1;  //170 / 127 = 1
    16'b10101010_10000000 : OUT <= 1;  //170 / 128 = 1
    16'b10101010_10000001 : OUT <= 1;  //170 / 129 = 1
    16'b10101010_10000010 : OUT <= 1;  //170 / 130 = 1
    16'b10101010_10000011 : OUT <= 1;  //170 / 131 = 1
    16'b10101010_10000100 : OUT <= 1;  //170 / 132 = 1
    16'b10101010_10000101 : OUT <= 1;  //170 / 133 = 1
    16'b10101010_10000110 : OUT <= 1;  //170 / 134 = 1
    16'b10101010_10000111 : OUT <= 1;  //170 / 135 = 1
    16'b10101010_10001000 : OUT <= 1;  //170 / 136 = 1
    16'b10101010_10001001 : OUT <= 1;  //170 / 137 = 1
    16'b10101010_10001010 : OUT <= 1;  //170 / 138 = 1
    16'b10101010_10001011 : OUT <= 1;  //170 / 139 = 1
    16'b10101010_10001100 : OUT <= 1;  //170 / 140 = 1
    16'b10101010_10001101 : OUT <= 1;  //170 / 141 = 1
    16'b10101010_10001110 : OUT <= 1;  //170 / 142 = 1
    16'b10101010_10001111 : OUT <= 1;  //170 / 143 = 1
    16'b10101010_10010000 : OUT <= 1;  //170 / 144 = 1
    16'b10101010_10010001 : OUT <= 1;  //170 / 145 = 1
    16'b10101010_10010010 : OUT <= 1;  //170 / 146 = 1
    16'b10101010_10010011 : OUT <= 1;  //170 / 147 = 1
    16'b10101010_10010100 : OUT <= 1;  //170 / 148 = 1
    16'b10101010_10010101 : OUT <= 1;  //170 / 149 = 1
    16'b10101010_10010110 : OUT <= 1;  //170 / 150 = 1
    16'b10101010_10010111 : OUT <= 1;  //170 / 151 = 1
    16'b10101010_10011000 : OUT <= 1;  //170 / 152 = 1
    16'b10101010_10011001 : OUT <= 1;  //170 / 153 = 1
    16'b10101010_10011010 : OUT <= 1;  //170 / 154 = 1
    16'b10101010_10011011 : OUT <= 1;  //170 / 155 = 1
    16'b10101010_10011100 : OUT <= 1;  //170 / 156 = 1
    16'b10101010_10011101 : OUT <= 1;  //170 / 157 = 1
    16'b10101010_10011110 : OUT <= 1;  //170 / 158 = 1
    16'b10101010_10011111 : OUT <= 1;  //170 / 159 = 1
    16'b10101010_10100000 : OUT <= 1;  //170 / 160 = 1
    16'b10101010_10100001 : OUT <= 1;  //170 / 161 = 1
    16'b10101010_10100010 : OUT <= 1;  //170 / 162 = 1
    16'b10101010_10100011 : OUT <= 1;  //170 / 163 = 1
    16'b10101010_10100100 : OUT <= 1;  //170 / 164 = 1
    16'b10101010_10100101 : OUT <= 1;  //170 / 165 = 1
    16'b10101010_10100110 : OUT <= 1;  //170 / 166 = 1
    16'b10101010_10100111 : OUT <= 1;  //170 / 167 = 1
    16'b10101010_10101000 : OUT <= 1;  //170 / 168 = 1
    16'b10101010_10101001 : OUT <= 1;  //170 / 169 = 1
    16'b10101010_10101010 : OUT <= 1;  //170 / 170 = 1
    16'b10101010_10101011 : OUT <= 0;  //170 / 171 = 0
    16'b10101010_10101100 : OUT <= 0;  //170 / 172 = 0
    16'b10101010_10101101 : OUT <= 0;  //170 / 173 = 0
    16'b10101010_10101110 : OUT <= 0;  //170 / 174 = 0
    16'b10101010_10101111 : OUT <= 0;  //170 / 175 = 0
    16'b10101010_10110000 : OUT <= 0;  //170 / 176 = 0
    16'b10101010_10110001 : OUT <= 0;  //170 / 177 = 0
    16'b10101010_10110010 : OUT <= 0;  //170 / 178 = 0
    16'b10101010_10110011 : OUT <= 0;  //170 / 179 = 0
    16'b10101010_10110100 : OUT <= 0;  //170 / 180 = 0
    16'b10101010_10110101 : OUT <= 0;  //170 / 181 = 0
    16'b10101010_10110110 : OUT <= 0;  //170 / 182 = 0
    16'b10101010_10110111 : OUT <= 0;  //170 / 183 = 0
    16'b10101010_10111000 : OUT <= 0;  //170 / 184 = 0
    16'b10101010_10111001 : OUT <= 0;  //170 / 185 = 0
    16'b10101010_10111010 : OUT <= 0;  //170 / 186 = 0
    16'b10101010_10111011 : OUT <= 0;  //170 / 187 = 0
    16'b10101010_10111100 : OUT <= 0;  //170 / 188 = 0
    16'b10101010_10111101 : OUT <= 0;  //170 / 189 = 0
    16'b10101010_10111110 : OUT <= 0;  //170 / 190 = 0
    16'b10101010_10111111 : OUT <= 0;  //170 / 191 = 0
    16'b10101010_11000000 : OUT <= 0;  //170 / 192 = 0
    16'b10101010_11000001 : OUT <= 0;  //170 / 193 = 0
    16'b10101010_11000010 : OUT <= 0;  //170 / 194 = 0
    16'b10101010_11000011 : OUT <= 0;  //170 / 195 = 0
    16'b10101010_11000100 : OUT <= 0;  //170 / 196 = 0
    16'b10101010_11000101 : OUT <= 0;  //170 / 197 = 0
    16'b10101010_11000110 : OUT <= 0;  //170 / 198 = 0
    16'b10101010_11000111 : OUT <= 0;  //170 / 199 = 0
    16'b10101010_11001000 : OUT <= 0;  //170 / 200 = 0
    16'b10101010_11001001 : OUT <= 0;  //170 / 201 = 0
    16'b10101010_11001010 : OUT <= 0;  //170 / 202 = 0
    16'b10101010_11001011 : OUT <= 0;  //170 / 203 = 0
    16'b10101010_11001100 : OUT <= 0;  //170 / 204 = 0
    16'b10101010_11001101 : OUT <= 0;  //170 / 205 = 0
    16'b10101010_11001110 : OUT <= 0;  //170 / 206 = 0
    16'b10101010_11001111 : OUT <= 0;  //170 / 207 = 0
    16'b10101010_11010000 : OUT <= 0;  //170 / 208 = 0
    16'b10101010_11010001 : OUT <= 0;  //170 / 209 = 0
    16'b10101010_11010010 : OUT <= 0;  //170 / 210 = 0
    16'b10101010_11010011 : OUT <= 0;  //170 / 211 = 0
    16'b10101010_11010100 : OUT <= 0;  //170 / 212 = 0
    16'b10101010_11010101 : OUT <= 0;  //170 / 213 = 0
    16'b10101010_11010110 : OUT <= 0;  //170 / 214 = 0
    16'b10101010_11010111 : OUT <= 0;  //170 / 215 = 0
    16'b10101010_11011000 : OUT <= 0;  //170 / 216 = 0
    16'b10101010_11011001 : OUT <= 0;  //170 / 217 = 0
    16'b10101010_11011010 : OUT <= 0;  //170 / 218 = 0
    16'b10101010_11011011 : OUT <= 0;  //170 / 219 = 0
    16'b10101010_11011100 : OUT <= 0;  //170 / 220 = 0
    16'b10101010_11011101 : OUT <= 0;  //170 / 221 = 0
    16'b10101010_11011110 : OUT <= 0;  //170 / 222 = 0
    16'b10101010_11011111 : OUT <= 0;  //170 / 223 = 0
    16'b10101010_11100000 : OUT <= 0;  //170 / 224 = 0
    16'b10101010_11100001 : OUT <= 0;  //170 / 225 = 0
    16'b10101010_11100010 : OUT <= 0;  //170 / 226 = 0
    16'b10101010_11100011 : OUT <= 0;  //170 / 227 = 0
    16'b10101010_11100100 : OUT <= 0;  //170 / 228 = 0
    16'b10101010_11100101 : OUT <= 0;  //170 / 229 = 0
    16'b10101010_11100110 : OUT <= 0;  //170 / 230 = 0
    16'b10101010_11100111 : OUT <= 0;  //170 / 231 = 0
    16'b10101010_11101000 : OUT <= 0;  //170 / 232 = 0
    16'b10101010_11101001 : OUT <= 0;  //170 / 233 = 0
    16'b10101010_11101010 : OUT <= 0;  //170 / 234 = 0
    16'b10101010_11101011 : OUT <= 0;  //170 / 235 = 0
    16'b10101010_11101100 : OUT <= 0;  //170 / 236 = 0
    16'b10101010_11101101 : OUT <= 0;  //170 / 237 = 0
    16'b10101010_11101110 : OUT <= 0;  //170 / 238 = 0
    16'b10101010_11101111 : OUT <= 0;  //170 / 239 = 0
    16'b10101010_11110000 : OUT <= 0;  //170 / 240 = 0
    16'b10101010_11110001 : OUT <= 0;  //170 / 241 = 0
    16'b10101010_11110010 : OUT <= 0;  //170 / 242 = 0
    16'b10101010_11110011 : OUT <= 0;  //170 / 243 = 0
    16'b10101010_11110100 : OUT <= 0;  //170 / 244 = 0
    16'b10101010_11110101 : OUT <= 0;  //170 / 245 = 0
    16'b10101010_11110110 : OUT <= 0;  //170 / 246 = 0
    16'b10101010_11110111 : OUT <= 0;  //170 / 247 = 0
    16'b10101010_11111000 : OUT <= 0;  //170 / 248 = 0
    16'b10101010_11111001 : OUT <= 0;  //170 / 249 = 0
    16'b10101010_11111010 : OUT <= 0;  //170 / 250 = 0
    16'b10101010_11111011 : OUT <= 0;  //170 / 251 = 0
    16'b10101010_11111100 : OUT <= 0;  //170 / 252 = 0
    16'b10101010_11111101 : OUT <= 0;  //170 / 253 = 0
    16'b10101010_11111110 : OUT <= 0;  //170 / 254 = 0
    16'b10101010_11111111 : OUT <= 0;  //170 / 255 = 0
    16'b10101011_00000000 : OUT <= 0;  //171 / 0 = 0
    16'b10101011_00000001 : OUT <= 171;  //171 / 1 = 171
    16'b10101011_00000010 : OUT <= 85;  //171 / 2 = 85
    16'b10101011_00000011 : OUT <= 57;  //171 / 3 = 57
    16'b10101011_00000100 : OUT <= 42;  //171 / 4 = 42
    16'b10101011_00000101 : OUT <= 34;  //171 / 5 = 34
    16'b10101011_00000110 : OUT <= 28;  //171 / 6 = 28
    16'b10101011_00000111 : OUT <= 24;  //171 / 7 = 24
    16'b10101011_00001000 : OUT <= 21;  //171 / 8 = 21
    16'b10101011_00001001 : OUT <= 19;  //171 / 9 = 19
    16'b10101011_00001010 : OUT <= 17;  //171 / 10 = 17
    16'b10101011_00001011 : OUT <= 15;  //171 / 11 = 15
    16'b10101011_00001100 : OUT <= 14;  //171 / 12 = 14
    16'b10101011_00001101 : OUT <= 13;  //171 / 13 = 13
    16'b10101011_00001110 : OUT <= 12;  //171 / 14 = 12
    16'b10101011_00001111 : OUT <= 11;  //171 / 15 = 11
    16'b10101011_00010000 : OUT <= 10;  //171 / 16 = 10
    16'b10101011_00010001 : OUT <= 10;  //171 / 17 = 10
    16'b10101011_00010010 : OUT <= 9;  //171 / 18 = 9
    16'b10101011_00010011 : OUT <= 9;  //171 / 19 = 9
    16'b10101011_00010100 : OUT <= 8;  //171 / 20 = 8
    16'b10101011_00010101 : OUT <= 8;  //171 / 21 = 8
    16'b10101011_00010110 : OUT <= 7;  //171 / 22 = 7
    16'b10101011_00010111 : OUT <= 7;  //171 / 23 = 7
    16'b10101011_00011000 : OUT <= 7;  //171 / 24 = 7
    16'b10101011_00011001 : OUT <= 6;  //171 / 25 = 6
    16'b10101011_00011010 : OUT <= 6;  //171 / 26 = 6
    16'b10101011_00011011 : OUT <= 6;  //171 / 27 = 6
    16'b10101011_00011100 : OUT <= 6;  //171 / 28 = 6
    16'b10101011_00011101 : OUT <= 5;  //171 / 29 = 5
    16'b10101011_00011110 : OUT <= 5;  //171 / 30 = 5
    16'b10101011_00011111 : OUT <= 5;  //171 / 31 = 5
    16'b10101011_00100000 : OUT <= 5;  //171 / 32 = 5
    16'b10101011_00100001 : OUT <= 5;  //171 / 33 = 5
    16'b10101011_00100010 : OUT <= 5;  //171 / 34 = 5
    16'b10101011_00100011 : OUT <= 4;  //171 / 35 = 4
    16'b10101011_00100100 : OUT <= 4;  //171 / 36 = 4
    16'b10101011_00100101 : OUT <= 4;  //171 / 37 = 4
    16'b10101011_00100110 : OUT <= 4;  //171 / 38 = 4
    16'b10101011_00100111 : OUT <= 4;  //171 / 39 = 4
    16'b10101011_00101000 : OUT <= 4;  //171 / 40 = 4
    16'b10101011_00101001 : OUT <= 4;  //171 / 41 = 4
    16'b10101011_00101010 : OUT <= 4;  //171 / 42 = 4
    16'b10101011_00101011 : OUT <= 3;  //171 / 43 = 3
    16'b10101011_00101100 : OUT <= 3;  //171 / 44 = 3
    16'b10101011_00101101 : OUT <= 3;  //171 / 45 = 3
    16'b10101011_00101110 : OUT <= 3;  //171 / 46 = 3
    16'b10101011_00101111 : OUT <= 3;  //171 / 47 = 3
    16'b10101011_00110000 : OUT <= 3;  //171 / 48 = 3
    16'b10101011_00110001 : OUT <= 3;  //171 / 49 = 3
    16'b10101011_00110010 : OUT <= 3;  //171 / 50 = 3
    16'b10101011_00110011 : OUT <= 3;  //171 / 51 = 3
    16'b10101011_00110100 : OUT <= 3;  //171 / 52 = 3
    16'b10101011_00110101 : OUT <= 3;  //171 / 53 = 3
    16'b10101011_00110110 : OUT <= 3;  //171 / 54 = 3
    16'b10101011_00110111 : OUT <= 3;  //171 / 55 = 3
    16'b10101011_00111000 : OUT <= 3;  //171 / 56 = 3
    16'b10101011_00111001 : OUT <= 3;  //171 / 57 = 3
    16'b10101011_00111010 : OUT <= 2;  //171 / 58 = 2
    16'b10101011_00111011 : OUT <= 2;  //171 / 59 = 2
    16'b10101011_00111100 : OUT <= 2;  //171 / 60 = 2
    16'b10101011_00111101 : OUT <= 2;  //171 / 61 = 2
    16'b10101011_00111110 : OUT <= 2;  //171 / 62 = 2
    16'b10101011_00111111 : OUT <= 2;  //171 / 63 = 2
    16'b10101011_01000000 : OUT <= 2;  //171 / 64 = 2
    16'b10101011_01000001 : OUT <= 2;  //171 / 65 = 2
    16'b10101011_01000010 : OUT <= 2;  //171 / 66 = 2
    16'b10101011_01000011 : OUT <= 2;  //171 / 67 = 2
    16'b10101011_01000100 : OUT <= 2;  //171 / 68 = 2
    16'b10101011_01000101 : OUT <= 2;  //171 / 69 = 2
    16'b10101011_01000110 : OUT <= 2;  //171 / 70 = 2
    16'b10101011_01000111 : OUT <= 2;  //171 / 71 = 2
    16'b10101011_01001000 : OUT <= 2;  //171 / 72 = 2
    16'b10101011_01001001 : OUT <= 2;  //171 / 73 = 2
    16'b10101011_01001010 : OUT <= 2;  //171 / 74 = 2
    16'b10101011_01001011 : OUT <= 2;  //171 / 75 = 2
    16'b10101011_01001100 : OUT <= 2;  //171 / 76 = 2
    16'b10101011_01001101 : OUT <= 2;  //171 / 77 = 2
    16'b10101011_01001110 : OUT <= 2;  //171 / 78 = 2
    16'b10101011_01001111 : OUT <= 2;  //171 / 79 = 2
    16'b10101011_01010000 : OUT <= 2;  //171 / 80 = 2
    16'b10101011_01010001 : OUT <= 2;  //171 / 81 = 2
    16'b10101011_01010010 : OUT <= 2;  //171 / 82 = 2
    16'b10101011_01010011 : OUT <= 2;  //171 / 83 = 2
    16'b10101011_01010100 : OUT <= 2;  //171 / 84 = 2
    16'b10101011_01010101 : OUT <= 2;  //171 / 85 = 2
    16'b10101011_01010110 : OUT <= 1;  //171 / 86 = 1
    16'b10101011_01010111 : OUT <= 1;  //171 / 87 = 1
    16'b10101011_01011000 : OUT <= 1;  //171 / 88 = 1
    16'b10101011_01011001 : OUT <= 1;  //171 / 89 = 1
    16'b10101011_01011010 : OUT <= 1;  //171 / 90 = 1
    16'b10101011_01011011 : OUT <= 1;  //171 / 91 = 1
    16'b10101011_01011100 : OUT <= 1;  //171 / 92 = 1
    16'b10101011_01011101 : OUT <= 1;  //171 / 93 = 1
    16'b10101011_01011110 : OUT <= 1;  //171 / 94 = 1
    16'b10101011_01011111 : OUT <= 1;  //171 / 95 = 1
    16'b10101011_01100000 : OUT <= 1;  //171 / 96 = 1
    16'b10101011_01100001 : OUT <= 1;  //171 / 97 = 1
    16'b10101011_01100010 : OUT <= 1;  //171 / 98 = 1
    16'b10101011_01100011 : OUT <= 1;  //171 / 99 = 1
    16'b10101011_01100100 : OUT <= 1;  //171 / 100 = 1
    16'b10101011_01100101 : OUT <= 1;  //171 / 101 = 1
    16'b10101011_01100110 : OUT <= 1;  //171 / 102 = 1
    16'b10101011_01100111 : OUT <= 1;  //171 / 103 = 1
    16'b10101011_01101000 : OUT <= 1;  //171 / 104 = 1
    16'b10101011_01101001 : OUT <= 1;  //171 / 105 = 1
    16'b10101011_01101010 : OUT <= 1;  //171 / 106 = 1
    16'b10101011_01101011 : OUT <= 1;  //171 / 107 = 1
    16'b10101011_01101100 : OUT <= 1;  //171 / 108 = 1
    16'b10101011_01101101 : OUT <= 1;  //171 / 109 = 1
    16'b10101011_01101110 : OUT <= 1;  //171 / 110 = 1
    16'b10101011_01101111 : OUT <= 1;  //171 / 111 = 1
    16'b10101011_01110000 : OUT <= 1;  //171 / 112 = 1
    16'b10101011_01110001 : OUT <= 1;  //171 / 113 = 1
    16'b10101011_01110010 : OUT <= 1;  //171 / 114 = 1
    16'b10101011_01110011 : OUT <= 1;  //171 / 115 = 1
    16'b10101011_01110100 : OUT <= 1;  //171 / 116 = 1
    16'b10101011_01110101 : OUT <= 1;  //171 / 117 = 1
    16'b10101011_01110110 : OUT <= 1;  //171 / 118 = 1
    16'b10101011_01110111 : OUT <= 1;  //171 / 119 = 1
    16'b10101011_01111000 : OUT <= 1;  //171 / 120 = 1
    16'b10101011_01111001 : OUT <= 1;  //171 / 121 = 1
    16'b10101011_01111010 : OUT <= 1;  //171 / 122 = 1
    16'b10101011_01111011 : OUT <= 1;  //171 / 123 = 1
    16'b10101011_01111100 : OUT <= 1;  //171 / 124 = 1
    16'b10101011_01111101 : OUT <= 1;  //171 / 125 = 1
    16'b10101011_01111110 : OUT <= 1;  //171 / 126 = 1
    16'b10101011_01111111 : OUT <= 1;  //171 / 127 = 1
    16'b10101011_10000000 : OUT <= 1;  //171 / 128 = 1
    16'b10101011_10000001 : OUT <= 1;  //171 / 129 = 1
    16'b10101011_10000010 : OUT <= 1;  //171 / 130 = 1
    16'b10101011_10000011 : OUT <= 1;  //171 / 131 = 1
    16'b10101011_10000100 : OUT <= 1;  //171 / 132 = 1
    16'b10101011_10000101 : OUT <= 1;  //171 / 133 = 1
    16'b10101011_10000110 : OUT <= 1;  //171 / 134 = 1
    16'b10101011_10000111 : OUT <= 1;  //171 / 135 = 1
    16'b10101011_10001000 : OUT <= 1;  //171 / 136 = 1
    16'b10101011_10001001 : OUT <= 1;  //171 / 137 = 1
    16'b10101011_10001010 : OUT <= 1;  //171 / 138 = 1
    16'b10101011_10001011 : OUT <= 1;  //171 / 139 = 1
    16'b10101011_10001100 : OUT <= 1;  //171 / 140 = 1
    16'b10101011_10001101 : OUT <= 1;  //171 / 141 = 1
    16'b10101011_10001110 : OUT <= 1;  //171 / 142 = 1
    16'b10101011_10001111 : OUT <= 1;  //171 / 143 = 1
    16'b10101011_10010000 : OUT <= 1;  //171 / 144 = 1
    16'b10101011_10010001 : OUT <= 1;  //171 / 145 = 1
    16'b10101011_10010010 : OUT <= 1;  //171 / 146 = 1
    16'b10101011_10010011 : OUT <= 1;  //171 / 147 = 1
    16'b10101011_10010100 : OUT <= 1;  //171 / 148 = 1
    16'b10101011_10010101 : OUT <= 1;  //171 / 149 = 1
    16'b10101011_10010110 : OUT <= 1;  //171 / 150 = 1
    16'b10101011_10010111 : OUT <= 1;  //171 / 151 = 1
    16'b10101011_10011000 : OUT <= 1;  //171 / 152 = 1
    16'b10101011_10011001 : OUT <= 1;  //171 / 153 = 1
    16'b10101011_10011010 : OUT <= 1;  //171 / 154 = 1
    16'b10101011_10011011 : OUT <= 1;  //171 / 155 = 1
    16'b10101011_10011100 : OUT <= 1;  //171 / 156 = 1
    16'b10101011_10011101 : OUT <= 1;  //171 / 157 = 1
    16'b10101011_10011110 : OUT <= 1;  //171 / 158 = 1
    16'b10101011_10011111 : OUT <= 1;  //171 / 159 = 1
    16'b10101011_10100000 : OUT <= 1;  //171 / 160 = 1
    16'b10101011_10100001 : OUT <= 1;  //171 / 161 = 1
    16'b10101011_10100010 : OUT <= 1;  //171 / 162 = 1
    16'b10101011_10100011 : OUT <= 1;  //171 / 163 = 1
    16'b10101011_10100100 : OUT <= 1;  //171 / 164 = 1
    16'b10101011_10100101 : OUT <= 1;  //171 / 165 = 1
    16'b10101011_10100110 : OUT <= 1;  //171 / 166 = 1
    16'b10101011_10100111 : OUT <= 1;  //171 / 167 = 1
    16'b10101011_10101000 : OUT <= 1;  //171 / 168 = 1
    16'b10101011_10101001 : OUT <= 1;  //171 / 169 = 1
    16'b10101011_10101010 : OUT <= 1;  //171 / 170 = 1
    16'b10101011_10101011 : OUT <= 1;  //171 / 171 = 1
    16'b10101011_10101100 : OUT <= 0;  //171 / 172 = 0
    16'b10101011_10101101 : OUT <= 0;  //171 / 173 = 0
    16'b10101011_10101110 : OUT <= 0;  //171 / 174 = 0
    16'b10101011_10101111 : OUT <= 0;  //171 / 175 = 0
    16'b10101011_10110000 : OUT <= 0;  //171 / 176 = 0
    16'b10101011_10110001 : OUT <= 0;  //171 / 177 = 0
    16'b10101011_10110010 : OUT <= 0;  //171 / 178 = 0
    16'b10101011_10110011 : OUT <= 0;  //171 / 179 = 0
    16'b10101011_10110100 : OUT <= 0;  //171 / 180 = 0
    16'b10101011_10110101 : OUT <= 0;  //171 / 181 = 0
    16'b10101011_10110110 : OUT <= 0;  //171 / 182 = 0
    16'b10101011_10110111 : OUT <= 0;  //171 / 183 = 0
    16'b10101011_10111000 : OUT <= 0;  //171 / 184 = 0
    16'b10101011_10111001 : OUT <= 0;  //171 / 185 = 0
    16'b10101011_10111010 : OUT <= 0;  //171 / 186 = 0
    16'b10101011_10111011 : OUT <= 0;  //171 / 187 = 0
    16'b10101011_10111100 : OUT <= 0;  //171 / 188 = 0
    16'b10101011_10111101 : OUT <= 0;  //171 / 189 = 0
    16'b10101011_10111110 : OUT <= 0;  //171 / 190 = 0
    16'b10101011_10111111 : OUT <= 0;  //171 / 191 = 0
    16'b10101011_11000000 : OUT <= 0;  //171 / 192 = 0
    16'b10101011_11000001 : OUT <= 0;  //171 / 193 = 0
    16'b10101011_11000010 : OUT <= 0;  //171 / 194 = 0
    16'b10101011_11000011 : OUT <= 0;  //171 / 195 = 0
    16'b10101011_11000100 : OUT <= 0;  //171 / 196 = 0
    16'b10101011_11000101 : OUT <= 0;  //171 / 197 = 0
    16'b10101011_11000110 : OUT <= 0;  //171 / 198 = 0
    16'b10101011_11000111 : OUT <= 0;  //171 / 199 = 0
    16'b10101011_11001000 : OUT <= 0;  //171 / 200 = 0
    16'b10101011_11001001 : OUT <= 0;  //171 / 201 = 0
    16'b10101011_11001010 : OUT <= 0;  //171 / 202 = 0
    16'b10101011_11001011 : OUT <= 0;  //171 / 203 = 0
    16'b10101011_11001100 : OUT <= 0;  //171 / 204 = 0
    16'b10101011_11001101 : OUT <= 0;  //171 / 205 = 0
    16'b10101011_11001110 : OUT <= 0;  //171 / 206 = 0
    16'b10101011_11001111 : OUT <= 0;  //171 / 207 = 0
    16'b10101011_11010000 : OUT <= 0;  //171 / 208 = 0
    16'b10101011_11010001 : OUT <= 0;  //171 / 209 = 0
    16'b10101011_11010010 : OUT <= 0;  //171 / 210 = 0
    16'b10101011_11010011 : OUT <= 0;  //171 / 211 = 0
    16'b10101011_11010100 : OUT <= 0;  //171 / 212 = 0
    16'b10101011_11010101 : OUT <= 0;  //171 / 213 = 0
    16'b10101011_11010110 : OUT <= 0;  //171 / 214 = 0
    16'b10101011_11010111 : OUT <= 0;  //171 / 215 = 0
    16'b10101011_11011000 : OUT <= 0;  //171 / 216 = 0
    16'b10101011_11011001 : OUT <= 0;  //171 / 217 = 0
    16'b10101011_11011010 : OUT <= 0;  //171 / 218 = 0
    16'b10101011_11011011 : OUT <= 0;  //171 / 219 = 0
    16'b10101011_11011100 : OUT <= 0;  //171 / 220 = 0
    16'b10101011_11011101 : OUT <= 0;  //171 / 221 = 0
    16'b10101011_11011110 : OUT <= 0;  //171 / 222 = 0
    16'b10101011_11011111 : OUT <= 0;  //171 / 223 = 0
    16'b10101011_11100000 : OUT <= 0;  //171 / 224 = 0
    16'b10101011_11100001 : OUT <= 0;  //171 / 225 = 0
    16'b10101011_11100010 : OUT <= 0;  //171 / 226 = 0
    16'b10101011_11100011 : OUT <= 0;  //171 / 227 = 0
    16'b10101011_11100100 : OUT <= 0;  //171 / 228 = 0
    16'b10101011_11100101 : OUT <= 0;  //171 / 229 = 0
    16'b10101011_11100110 : OUT <= 0;  //171 / 230 = 0
    16'b10101011_11100111 : OUT <= 0;  //171 / 231 = 0
    16'b10101011_11101000 : OUT <= 0;  //171 / 232 = 0
    16'b10101011_11101001 : OUT <= 0;  //171 / 233 = 0
    16'b10101011_11101010 : OUT <= 0;  //171 / 234 = 0
    16'b10101011_11101011 : OUT <= 0;  //171 / 235 = 0
    16'b10101011_11101100 : OUT <= 0;  //171 / 236 = 0
    16'b10101011_11101101 : OUT <= 0;  //171 / 237 = 0
    16'b10101011_11101110 : OUT <= 0;  //171 / 238 = 0
    16'b10101011_11101111 : OUT <= 0;  //171 / 239 = 0
    16'b10101011_11110000 : OUT <= 0;  //171 / 240 = 0
    16'b10101011_11110001 : OUT <= 0;  //171 / 241 = 0
    16'b10101011_11110010 : OUT <= 0;  //171 / 242 = 0
    16'b10101011_11110011 : OUT <= 0;  //171 / 243 = 0
    16'b10101011_11110100 : OUT <= 0;  //171 / 244 = 0
    16'b10101011_11110101 : OUT <= 0;  //171 / 245 = 0
    16'b10101011_11110110 : OUT <= 0;  //171 / 246 = 0
    16'b10101011_11110111 : OUT <= 0;  //171 / 247 = 0
    16'b10101011_11111000 : OUT <= 0;  //171 / 248 = 0
    16'b10101011_11111001 : OUT <= 0;  //171 / 249 = 0
    16'b10101011_11111010 : OUT <= 0;  //171 / 250 = 0
    16'b10101011_11111011 : OUT <= 0;  //171 / 251 = 0
    16'b10101011_11111100 : OUT <= 0;  //171 / 252 = 0
    16'b10101011_11111101 : OUT <= 0;  //171 / 253 = 0
    16'b10101011_11111110 : OUT <= 0;  //171 / 254 = 0
    16'b10101011_11111111 : OUT <= 0;  //171 / 255 = 0
    16'b10101100_00000000 : OUT <= 0;  //172 / 0 = 0
    16'b10101100_00000001 : OUT <= 172;  //172 / 1 = 172
    16'b10101100_00000010 : OUT <= 86;  //172 / 2 = 86
    16'b10101100_00000011 : OUT <= 57;  //172 / 3 = 57
    16'b10101100_00000100 : OUT <= 43;  //172 / 4 = 43
    16'b10101100_00000101 : OUT <= 34;  //172 / 5 = 34
    16'b10101100_00000110 : OUT <= 28;  //172 / 6 = 28
    16'b10101100_00000111 : OUT <= 24;  //172 / 7 = 24
    16'b10101100_00001000 : OUT <= 21;  //172 / 8 = 21
    16'b10101100_00001001 : OUT <= 19;  //172 / 9 = 19
    16'b10101100_00001010 : OUT <= 17;  //172 / 10 = 17
    16'b10101100_00001011 : OUT <= 15;  //172 / 11 = 15
    16'b10101100_00001100 : OUT <= 14;  //172 / 12 = 14
    16'b10101100_00001101 : OUT <= 13;  //172 / 13 = 13
    16'b10101100_00001110 : OUT <= 12;  //172 / 14 = 12
    16'b10101100_00001111 : OUT <= 11;  //172 / 15 = 11
    16'b10101100_00010000 : OUT <= 10;  //172 / 16 = 10
    16'b10101100_00010001 : OUT <= 10;  //172 / 17 = 10
    16'b10101100_00010010 : OUT <= 9;  //172 / 18 = 9
    16'b10101100_00010011 : OUT <= 9;  //172 / 19 = 9
    16'b10101100_00010100 : OUT <= 8;  //172 / 20 = 8
    16'b10101100_00010101 : OUT <= 8;  //172 / 21 = 8
    16'b10101100_00010110 : OUT <= 7;  //172 / 22 = 7
    16'b10101100_00010111 : OUT <= 7;  //172 / 23 = 7
    16'b10101100_00011000 : OUT <= 7;  //172 / 24 = 7
    16'b10101100_00011001 : OUT <= 6;  //172 / 25 = 6
    16'b10101100_00011010 : OUT <= 6;  //172 / 26 = 6
    16'b10101100_00011011 : OUT <= 6;  //172 / 27 = 6
    16'b10101100_00011100 : OUT <= 6;  //172 / 28 = 6
    16'b10101100_00011101 : OUT <= 5;  //172 / 29 = 5
    16'b10101100_00011110 : OUT <= 5;  //172 / 30 = 5
    16'b10101100_00011111 : OUT <= 5;  //172 / 31 = 5
    16'b10101100_00100000 : OUT <= 5;  //172 / 32 = 5
    16'b10101100_00100001 : OUT <= 5;  //172 / 33 = 5
    16'b10101100_00100010 : OUT <= 5;  //172 / 34 = 5
    16'b10101100_00100011 : OUT <= 4;  //172 / 35 = 4
    16'b10101100_00100100 : OUT <= 4;  //172 / 36 = 4
    16'b10101100_00100101 : OUT <= 4;  //172 / 37 = 4
    16'b10101100_00100110 : OUT <= 4;  //172 / 38 = 4
    16'b10101100_00100111 : OUT <= 4;  //172 / 39 = 4
    16'b10101100_00101000 : OUT <= 4;  //172 / 40 = 4
    16'b10101100_00101001 : OUT <= 4;  //172 / 41 = 4
    16'b10101100_00101010 : OUT <= 4;  //172 / 42 = 4
    16'b10101100_00101011 : OUT <= 4;  //172 / 43 = 4
    16'b10101100_00101100 : OUT <= 3;  //172 / 44 = 3
    16'b10101100_00101101 : OUT <= 3;  //172 / 45 = 3
    16'b10101100_00101110 : OUT <= 3;  //172 / 46 = 3
    16'b10101100_00101111 : OUT <= 3;  //172 / 47 = 3
    16'b10101100_00110000 : OUT <= 3;  //172 / 48 = 3
    16'b10101100_00110001 : OUT <= 3;  //172 / 49 = 3
    16'b10101100_00110010 : OUT <= 3;  //172 / 50 = 3
    16'b10101100_00110011 : OUT <= 3;  //172 / 51 = 3
    16'b10101100_00110100 : OUT <= 3;  //172 / 52 = 3
    16'b10101100_00110101 : OUT <= 3;  //172 / 53 = 3
    16'b10101100_00110110 : OUT <= 3;  //172 / 54 = 3
    16'b10101100_00110111 : OUT <= 3;  //172 / 55 = 3
    16'b10101100_00111000 : OUT <= 3;  //172 / 56 = 3
    16'b10101100_00111001 : OUT <= 3;  //172 / 57 = 3
    16'b10101100_00111010 : OUT <= 2;  //172 / 58 = 2
    16'b10101100_00111011 : OUT <= 2;  //172 / 59 = 2
    16'b10101100_00111100 : OUT <= 2;  //172 / 60 = 2
    16'b10101100_00111101 : OUT <= 2;  //172 / 61 = 2
    16'b10101100_00111110 : OUT <= 2;  //172 / 62 = 2
    16'b10101100_00111111 : OUT <= 2;  //172 / 63 = 2
    16'b10101100_01000000 : OUT <= 2;  //172 / 64 = 2
    16'b10101100_01000001 : OUT <= 2;  //172 / 65 = 2
    16'b10101100_01000010 : OUT <= 2;  //172 / 66 = 2
    16'b10101100_01000011 : OUT <= 2;  //172 / 67 = 2
    16'b10101100_01000100 : OUT <= 2;  //172 / 68 = 2
    16'b10101100_01000101 : OUT <= 2;  //172 / 69 = 2
    16'b10101100_01000110 : OUT <= 2;  //172 / 70 = 2
    16'b10101100_01000111 : OUT <= 2;  //172 / 71 = 2
    16'b10101100_01001000 : OUT <= 2;  //172 / 72 = 2
    16'b10101100_01001001 : OUT <= 2;  //172 / 73 = 2
    16'b10101100_01001010 : OUT <= 2;  //172 / 74 = 2
    16'b10101100_01001011 : OUT <= 2;  //172 / 75 = 2
    16'b10101100_01001100 : OUT <= 2;  //172 / 76 = 2
    16'b10101100_01001101 : OUT <= 2;  //172 / 77 = 2
    16'b10101100_01001110 : OUT <= 2;  //172 / 78 = 2
    16'b10101100_01001111 : OUT <= 2;  //172 / 79 = 2
    16'b10101100_01010000 : OUT <= 2;  //172 / 80 = 2
    16'b10101100_01010001 : OUT <= 2;  //172 / 81 = 2
    16'b10101100_01010010 : OUT <= 2;  //172 / 82 = 2
    16'b10101100_01010011 : OUT <= 2;  //172 / 83 = 2
    16'b10101100_01010100 : OUT <= 2;  //172 / 84 = 2
    16'b10101100_01010101 : OUT <= 2;  //172 / 85 = 2
    16'b10101100_01010110 : OUT <= 2;  //172 / 86 = 2
    16'b10101100_01010111 : OUT <= 1;  //172 / 87 = 1
    16'b10101100_01011000 : OUT <= 1;  //172 / 88 = 1
    16'b10101100_01011001 : OUT <= 1;  //172 / 89 = 1
    16'b10101100_01011010 : OUT <= 1;  //172 / 90 = 1
    16'b10101100_01011011 : OUT <= 1;  //172 / 91 = 1
    16'b10101100_01011100 : OUT <= 1;  //172 / 92 = 1
    16'b10101100_01011101 : OUT <= 1;  //172 / 93 = 1
    16'b10101100_01011110 : OUT <= 1;  //172 / 94 = 1
    16'b10101100_01011111 : OUT <= 1;  //172 / 95 = 1
    16'b10101100_01100000 : OUT <= 1;  //172 / 96 = 1
    16'b10101100_01100001 : OUT <= 1;  //172 / 97 = 1
    16'b10101100_01100010 : OUT <= 1;  //172 / 98 = 1
    16'b10101100_01100011 : OUT <= 1;  //172 / 99 = 1
    16'b10101100_01100100 : OUT <= 1;  //172 / 100 = 1
    16'b10101100_01100101 : OUT <= 1;  //172 / 101 = 1
    16'b10101100_01100110 : OUT <= 1;  //172 / 102 = 1
    16'b10101100_01100111 : OUT <= 1;  //172 / 103 = 1
    16'b10101100_01101000 : OUT <= 1;  //172 / 104 = 1
    16'b10101100_01101001 : OUT <= 1;  //172 / 105 = 1
    16'b10101100_01101010 : OUT <= 1;  //172 / 106 = 1
    16'b10101100_01101011 : OUT <= 1;  //172 / 107 = 1
    16'b10101100_01101100 : OUT <= 1;  //172 / 108 = 1
    16'b10101100_01101101 : OUT <= 1;  //172 / 109 = 1
    16'b10101100_01101110 : OUT <= 1;  //172 / 110 = 1
    16'b10101100_01101111 : OUT <= 1;  //172 / 111 = 1
    16'b10101100_01110000 : OUT <= 1;  //172 / 112 = 1
    16'b10101100_01110001 : OUT <= 1;  //172 / 113 = 1
    16'b10101100_01110010 : OUT <= 1;  //172 / 114 = 1
    16'b10101100_01110011 : OUT <= 1;  //172 / 115 = 1
    16'b10101100_01110100 : OUT <= 1;  //172 / 116 = 1
    16'b10101100_01110101 : OUT <= 1;  //172 / 117 = 1
    16'b10101100_01110110 : OUT <= 1;  //172 / 118 = 1
    16'b10101100_01110111 : OUT <= 1;  //172 / 119 = 1
    16'b10101100_01111000 : OUT <= 1;  //172 / 120 = 1
    16'b10101100_01111001 : OUT <= 1;  //172 / 121 = 1
    16'b10101100_01111010 : OUT <= 1;  //172 / 122 = 1
    16'b10101100_01111011 : OUT <= 1;  //172 / 123 = 1
    16'b10101100_01111100 : OUT <= 1;  //172 / 124 = 1
    16'b10101100_01111101 : OUT <= 1;  //172 / 125 = 1
    16'b10101100_01111110 : OUT <= 1;  //172 / 126 = 1
    16'b10101100_01111111 : OUT <= 1;  //172 / 127 = 1
    16'b10101100_10000000 : OUT <= 1;  //172 / 128 = 1
    16'b10101100_10000001 : OUT <= 1;  //172 / 129 = 1
    16'b10101100_10000010 : OUT <= 1;  //172 / 130 = 1
    16'b10101100_10000011 : OUT <= 1;  //172 / 131 = 1
    16'b10101100_10000100 : OUT <= 1;  //172 / 132 = 1
    16'b10101100_10000101 : OUT <= 1;  //172 / 133 = 1
    16'b10101100_10000110 : OUT <= 1;  //172 / 134 = 1
    16'b10101100_10000111 : OUT <= 1;  //172 / 135 = 1
    16'b10101100_10001000 : OUT <= 1;  //172 / 136 = 1
    16'b10101100_10001001 : OUT <= 1;  //172 / 137 = 1
    16'b10101100_10001010 : OUT <= 1;  //172 / 138 = 1
    16'b10101100_10001011 : OUT <= 1;  //172 / 139 = 1
    16'b10101100_10001100 : OUT <= 1;  //172 / 140 = 1
    16'b10101100_10001101 : OUT <= 1;  //172 / 141 = 1
    16'b10101100_10001110 : OUT <= 1;  //172 / 142 = 1
    16'b10101100_10001111 : OUT <= 1;  //172 / 143 = 1
    16'b10101100_10010000 : OUT <= 1;  //172 / 144 = 1
    16'b10101100_10010001 : OUT <= 1;  //172 / 145 = 1
    16'b10101100_10010010 : OUT <= 1;  //172 / 146 = 1
    16'b10101100_10010011 : OUT <= 1;  //172 / 147 = 1
    16'b10101100_10010100 : OUT <= 1;  //172 / 148 = 1
    16'b10101100_10010101 : OUT <= 1;  //172 / 149 = 1
    16'b10101100_10010110 : OUT <= 1;  //172 / 150 = 1
    16'b10101100_10010111 : OUT <= 1;  //172 / 151 = 1
    16'b10101100_10011000 : OUT <= 1;  //172 / 152 = 1
    16'b10101100_10011001 : OUT <= 1;  //172 / 153 = 1
    16'b10101100_10011010 : OUT <= 1;  //172 / 154 = 1
    16'b10101100_10011011 : OUT <= 1;  //172 / 155 = 1
    16'b10101100_10011100 : OUT <= 1;  //172 / 156 = 1
    16'b10101100_10011101 : OUT <= 1;  //172 / 157 = 1
    16'b10101100_10011110 : OUT <= 1;  //172 / 158 = 1
    16'b10101100_10011111 : OUT <= 1;  //172 / 159 = 1
    16'b10101100_10100000 : OUT <= 1;  //172 / 160 = 1
    16'b10101100_10100001 : OUT <= 1;  //172 / 161 = 1
    16'b10101100_10100010 : OUT <= 1;  //172 / 162 = 1
    16'b10101100_10100011 : OUT <= 1;  //172 / 163 = 1
    16'b10101100_10100100 : OUT <= 1;  //172 / 164 = 1
    16'b10101100_10100101 : OUT <= 1;  //172 / 165 = 1
    16'b10101100_10100110 : OUT <= 1;  //172 / 166 = 1
    16'b10101100_10100111 : OUT <= 1;  //172 / 167 = 1
    16'b10101100_10101000 : OUT <= 1;  //172 / 168 = 1
    16'b10101100_10101001 : OUT <= 1;  //172 / 169 = 1
    16'b10101100_10101010 : OUT <= 1;  //172 / 170 = 1
    16'b10101100_10101011 : OUT <= 1;  //172 / 171 = 1
    16'b10101100_10101100 : OUT <= 1;  //172 / 172 = 1
    16'b10101100_10101101 : OUT <= 0;  //172 / 173 = 0
    16'b10101100_10101110 : OUT <= 0;  //172 / 174 = 0
    16'b10101100_10101111 : OUT <= 0;  //172 / 175 = 0
    16'b10101100_10110000 : OUT <= 0;  //172 / 176 = 0
    16'b10101100_10110001 : OUT <= 0;  //172 / 177 = 0
    16'b10101100_10110010 : OUT <= 0;  //172 / 178 = 0
    16'b10101100_10110011 : OUT <= 0;  //172 / 179 = 0
    16'b10101100_10110100 : OUT <= 0;  //172 / 180 = 0
    16'b10101100_10110101 : OUT <= 0;  //172 / 181 = 0
    16'b10101100_10110110 : OUT <= 0;  //172 / 182 = 0
    16'b10101100_10110111 : OUT <= 0;  //172 / 183 = 0
    16'b10101100_10111000 : OUT <= 0;  //172 / 184 = 0
    16'b10101100_10111001 : OUT <= 0;  //172 / 185 = 0
    16'b10101100_10111010 : OUT <= 0;  //172 / 186 = 0
    16'b10101100_10111011 : OUT <= 0;  //172 / 187 = 0
    16'b10101100_10111100 : OUT <= 0;  //172 / 188 = 0
    16'b10101100_10111101 : OUT <= 0;  //172 / 189 = 0
    16'b10101100_10111110 : OUT <= 0;  //172 / 190 = 0
    16'b10101100_10111111 : OUT <= 0;  //172 / 191 = 0
    16'b10101100_11000000 : OUT <= 0;  //172 / 192 = 0
    16'b10101100_11000001 : OUT <= 0;  //172 / 193 = 0
    16'b10101100_11000010 : OUT <= 0;  //172 / 194 = 0
    16'b10101100_11000011 : OUT <= 0;  //172 / 195 = 0
    16'b10101100_11000100 : OUT <= 0;  //172 / 196 = 0
    16'b10101100_11000101 : OUT <= 0;  //172 / 197 = 0
    16'b10101100_11000110 : OUT <= 0;  //172 / 198 = 0
    16'b10101100_11000111 : OUT <= 0;  //172 / 199 = 0
    16'b10101100_11001000 : OUT <= 0;  //172 / 200 = 0
    16'b10101100_11001001 : OUT <= 0;  //172 / 201 = 0
    16'b10101100_11001010 : OUT <= 0;  //172 / 202 = 0
    16'b10101100_11001011 : OUT <= 0;  //172 / 203 = 0
    16'b10101100_11001100 : OUT <= 0;  //172 / 204 = 0
    16'b10101100_11001101 : OUT <= 0;  //172 / 205 = 0
    16'b10101100_11001110 : OUT <= 0;  //172 / 206 = 0
    16'b10101100_11001111 : OUT <= 0;  //172 / 207 = 0
    16'b10101100_11010000 : OUT <= 0;  //172 / 208 = 0
    16'b10101100_11010001 : OUT <= 0;  //172 / 209 = 0
    16'b10101100_11010010 : OUT <= 0;  //172 / 210 = 0
    16'b10101100_11010011 : OUT <= 0;  //172 / 211 = 0
    16'b10101100_11010100 : OUT <= 0;  //172 / 212 = 0
    16'b10101100_11010101 : OUT <= 0;  //172 / 213 = 0
    16'b10101100_11010110 : OUT <= 0;  //172 / 214 = 0
    16'b10101100_11010111 : OUT <= 0;  //172 / 215 = 0
    16'b10101100_11011000 : OUT <= 0;  //172 / 216 = 0
    16'b10101100_11011001 : OUT <= 0;  //172 / 217 = 0
    16'b10101100_11011010 : OUT <= 0;  //172 / 218 = 0
    16'b10101100_11011011 : OUT <= 0;  //172 / 219 = 0
    16'b10101100_11011100 : OUT <= 0;  //172 / 220 = 0
    16'b10101100_11011101 : OUT <= 0;  //172 / 221 = 0
    16'b10101100_11011110 : OUT <= 0;  //172 / 222 = 0
    16'b10101100_11011111 : OUT <= 0;  //172 / 223 = 0
    16'b10101100_11100000 : OUT <= 0;  //172 / 224 = 0
    16'b10101100_11100001 : OUT <= 0;  //172 / 225 = 0
    16'b10101100_11100010 : OUT <= 0;  //172 / 226 = 0
    16'b10101100_11100011 : OUT <= 0;  //172 / 227 = 0
    16'b10101100_11100100 : OUT <= 0;  //172 / 228 = 0
    16'b10101100_11100101 : OUT <= 0;  //172 / 229 = 0
    16'b10101100_11100110 : OUT <= 0;  //172 / 230 = 0
    16'b10101100_11100111 : OUT <= 0;  //172 / 231 = 0
    16'b10101100_11101000 : OUT <= 0;  //172 / 232 = 0
    16'b10101100_11101001 : OUT <= 0;  //172 / 233 = 0
    16'b10101100_11101010 : OUT <= 0;  //172 / 234 = 0
    16'b10101100_11101011 : OUT <= 0;  //172 / 235 = 0
    16'b10101100_11101100 : OUT <= 0;  //172 / 236 = 0
    16'b10101100_11101101 : OUT <= 0;  //172 / 237 = 0
    16'b10101100_11101110 : OUT <= 0;  //172 / 238 = 0
    16'b10101100_11101111 : OUT <= 0;  //172 / 239 = 0
    16'b10101100_11110000 : OUT <= 0;  //172 / 240 = 0
    16'b10101100_11110001 : OUT <= 0;  //172 / 241 = 0
    16'b10101100_11110010 : OUT <= 0;  //172 / 242 = 0
    16'b10101100_11110011 : OUT <= 0;  //172 / 243 = 0
    16'b10101100_11110100 : OUT <= 0;  //172 / 244 = 0
    16'b10101100_11110101 : OUT <= 0;  //172 / 245 = 0
    16'b10101100_11110110 : OUT <= 0;  //172 / 246 = 0
    16'b10101100_11110111 : OUT <= 0;  //172 / 247 = 0
    16'b10101100_11111000 : OUT <= 0;  //172 / 248 = 0
    16'b10101100_11111001 : OUT <= 0;  //172 / 249 = 0
    16'b10101100_11111010 : OUT <= 0;  //172 / 250 = 0
    16'b10101100_11111011 : OUT <= 0;  //172 / 251 = 0
    16'b10101100_11111100 : OUT <= 0;  //172 / 252 = 0
    16'b10101100_11111101 : OUT <= 0;  //172 / 253 = 0
    16'b10101100_11111110 : OUT <= 0;  //172 / 254 = 0
    16'b10101100_11111111 : OUT <= 0;  //172 / 255 = 0
    16'b10101101_00000000 : OUT <= 0;  //173 / 0 = 0
    16'b10101101_00000001 : OUT <= 173;  //173 / 1 = 173
    16'b10101101_00000010 : OUT <= 86;  //173 / 2 = 86
    16'b10101101_00000011 : OUT <= 57;  //173 / 3 = 57
    16'b10101101_00000100 : OUT <= 43;  //173 / 4 = 43
    16'b10101101_00000101 : OUT <= 34;  //173 / 5 = 34
    16'b10101101_00000110 : OUT <= 28;  //173 / 6 = 28
    16'b10101101_00000111 : OUT <= 24;  //173 / 7 = 24
    16'b10101101_00001000 : OUT <= 21;  //173 / 8 = 21
    16'b10101101_00001001 : OUT <= 19;  //173 / 9 = 19
    16'b10101101_00001010 : OUT <= 17;  //173 / 10 = 17
    16'b10101101_00001011 : OUT <= 15;  //173 / 11 = 15
    16'b10101101_00001100 : OUT <= 14;  //173 / 12 = 14
    16'b10101101_00001101 : OUT <= 13;  //173 / 13 = 13
    16'b10101101_00001110 : OUT <= 12;  //173 / 14 = 12
    16'b10101101_00001111 : OUT <= 11;  //173 / 15 = 11
    16'b10101101_00010000 : OUT <= 10;  //173 / 16 = 10
    16'b10101101_00010001 : OUT <= 10;  //173 / 17 = 10
    16'b10101101_00010010 : OUT <= 9;  //173 / 18 = 9
    16'b10101101_00010011 : OUT <= 9;  //173 / 19 = 9
    16'b10101101_00010100 : OUT <= 8;  //173 / 20 = 8
    16'b10101101_00010101 : OUT <= 8;  //173 / 21 = 8
    16'b10101101_00010110 : OUT <= 7;  //173 / 22 = 7
    16'b10101101_00010111 : OUT <= 7;  //173 / 23 = 7
    16'b10101101_00011000 : OUT <= 7;  //173 / 24 = 7
    16'b10101101_00011001 : OUT <= 6;  //173 / 25 = 6
    16'b10101101_00011010 : OUT <= 6;  //173 / 26 = 6
    16'b10101101_00011011 : OUT <= 6;  //173 / 27 = 6
    16'b10101101_00011100 : OUT <= 6;  //173 / 28 = 6
    16'b10101101_00011101 : OUT <= 5;  //173 / 29 = 5
    16'b10101101_00011110 : OUT <= 5;  //173 / 30 = 5
    16'b10101101_00011111 : OUT <= 5;  //173 / 31 = 5
    16'b10101101_00100000 : OUT <= 5;  //173 / 32 = 5
    16'b10101101_00100001 : OUT <= 5;  //173 / 33 = 5
    16'b10101101_00100010 : OUT <= 5;  //173 / 34 = 5
    16'b10101101_00100011 : OUT <= 4;  //173 / 35 = 4
    16'b10101101_00100100 : OUT <= 4;  //173 / 36 = 4
    16'b10101101_00100101 : OUT <= 4;  //173 / 37 = 4
    16'b10101101_00100110 : OUT <= 4;  //173 / 38 = 4
    16'b10101101_00100111 : OUT <= 4;  //173 / 39 = 4
    16'b10101101_00101000 : OUT <= 4;  //173 / 40 = 4
    16'b10101101_00101001 : OUT <= 4;  //173 / 41 = 4
    16'b10101101_00101010 : OUT <= 4;  //173 / 42 = 4
    16'b10101101_00101011 : OUT <= 4;  //173 / 43 = 4
    16'b10101101_00101100 : OUT <= 3;  //173 / 44 = 3
    16'b10101101_00101101 : OUT <= 3;  //173 / 45 = 3
    16'b10101101_00101110 : OUT <= 3;  //173 / 46 = 3
    16'b10101101_00101111 : OUT <= 3;  //173 / 47 = 3
    16'b10101101_00110000 : OUT <= 3;  //173 / 48 = 3
    16'b10101101_00110001 : OUT <= 3;  //173 / 49 = 3
    16'b10101101_00110010 : OUT <= 3;  //173 / 50 = 3
    16'b10101101_00110011 : OUT <= 3;  //173 / 51 = 3
    16'b10101101_00110100 : OUT <= 3;  //173 / 52 = 3
    16'b10101101_00110101 : OUT <= 3;  //173 / 53 = 3
    16'b10101101_00110110 : OUT <= 3;  //173 / 54 = 3
    16'b10101101_00110111 : OUT <= 3;  //173 / 55 = 3
    16'b10101101_00111000 : OUT <= 3;  //173 / 56 = 3
    16'b10101101_00111001 : OUT <= 3;  //173 / 57 = 3
    16'b10101101_00111010 : OUT <= 2;  //173 / 58 = 2
    16'b10101101_00111011 : OUT <= 2;  //173 / 59 = 2
    16'b10101101_00111100 : OUT <= 2;  //173 / 60 = 2
    16'b10101101_00111101 : OUT <= 2;  //173 / 61 = 2
    16'b10101101_00111110 : OUT <= 2;  //173 / 62 = 2
    16'b10101101_00111111 : OUT <= 2;  //173 / 63 = 2
    16'b10101101_01000000 : OUT <= 2;  //173 / 64 = 2
    16'b10101101_01000001 : OUT <= 2;  //173 / 65 = 2
    16'b10101101_01000010 : OUT <= 2;  //173 / 66 = 2
    16'b10101101_01000011 : OUT <= 2;  //173 / 67 = 2
    16'b10101101_01000100 : OUT <= 2;  //173 / 68 = 2
    16'b10101101_01000101 : OUT <= 2;  //173 / 69 = 2
    16'b10101101_01000110 : OUT <= 2;  //173 / 70 = 2
    16'b10101101_01000111 : OUT <= 2;  //173 / 71 = 2
    16'b10101101_01001000 : OUT <= 2;  //173 / 72 = 2
    16'b10101101_01001001 : OUT <= 2;  //173 / 73 = 2
    16'b10101101_01001010 : OUT <= 2;  //173 / 74 = 2
    16'b10101101_01001011 : OUT <= 2;  //173 / 75 = 2
    16'b10101101_01001100 : OUT <= 2;  //173 / 76 = 2
    16'b10101101_01001101 : OUT <= 2;  //173 / 77 = 2
    16'b10101101_01001110 : OUT <= 2;  //173 / 78 = 2
    16'b10101101_01001111 : OUT <= 2;  //173 / 79 = 2
    16'b10101101_01010000 : OUT <= 2;  //173 / 80 = 2
    16'b10101101_01010001 : OUT <= 2;  //173 / 81 = 2
    16'b10101101_01010010 : OUT <= 2;  //173 / 82 = 2
    16'b10101101_01010011 : OUT <= 2;  //173 / 83 = 2
    16'b10101101_01010100 : OUT <= 2;  //173 / 84 = 2
    16'b10101101_01010101 : OUT <= 2;  //173 / 85 = 2
    16'b10101101_01010110 : OUT <= 2;  //173 / 86 = 2
    16'b10101101_01010111 : OUT <= 1;  //173 / 87 = 1
    16'b10101101_01011000 : OUT <= 1;  //173 / 88 = 1
    16'b10101101_01011001 : OUT <= 1;  //173 / 89 = 1
    16'b10101101_01011010 : OUT <= 1;  //173 / 90 = 1
    16'b10101101_01011011 : OUT <= 1;  //173 / 91 = 1
    16'b10101101_01011100 : OUT <= 1;  //173 / 92 = 1
    16'b10101101_01011101 : OUT <= 1;  //173 / 93 = 1
    16'b10101101_01011110 : OUT <= 1;  //173 / 94 = 1
    16'b10101101_01011111 : OUT <= 1;  //173 / 95 = 1
    16'b10101101_01100000 : OUT <= 1;  //173 / 96 = 1
    16'b10101101_01100001 : OUT <= 1;  //173 / 97 = 1
    16'b10101101_01100010 : OUT <= 1;  //173 / 98 = 1
    16'b10101101_01100011 : OUT <= 1;  //173 / 99 = 1
    16'b10101101_01100100 : OUT <= 1;  //173 / 100 = 1
    16'b10101101_01100101 : OUT <= 1;  //173 / 101 = 1
    16'b10101101_01100110 : OUT <= 1;  //173 / 102 = 1
    16'b10101101_01100111 : OUT <= 1;  //173 / 103 = 1
    16'b10101101_01101000 : OUT <= 1;  //173 / 104 = 1
    16'b10101101_01101001 : OUT <= 1;  //173 / 105 = 1
    16'b10101101_01101010 : OUT <= 1;  //173 / 106 = 1
    16'b10101101_01101011 : OUT <= 1;  //173 / 107 = 1
    16'b10101101_01101100 : OUT <= 1;  //173 / 108 = 1
    16'b10101101_01101101 : OUT <= 1;  //173 / 109 = 1
    16'b10101101_01101110 : OUT <= 1;  //173 / 110 = 1
    16'b10101101_01101111 : OUT <= 1;  //173 / 111 = 1
    16'b10101101_01110000 : OUT <= 1;  //173 / 112 = 1
    16'b10101101_01110001 : OUT <= 1;  //173 / 113 = 1
    16'b10101101_01110010 : OUT <= 1;  //173 / 114 = 1
    16'b10101101_01110011 : OUT <= 1;  //173 / 115 = 1
    16'b10101101_01110100 : OUT <= 1;  //173 / 116 = 1
    16'b10101101_01110101 : OUT <= 1;  //173 / 117 = 1
    16'b10101101_01110110 : OUT <= 1;  //173 / 118 = 1
    16'b10101101_01110111 : OUT <= 1;  //173 / 119 = 1
    16'b10101101_01111000 : OUT <= 1;  //173 / 120 = 1
    16'b10101101_01111001 : OUT <= 1;  //173 / 121 = 1
    16'b10101101_01111010 : OUT <= 1;  //173 / 122 = 1
    16'b10101101_01111011 : OUT <= 1;  //173 / 123 = 1
    16'b10101101_01111100 : OUT <= 1;  //173 / 124 = 1
    16'b10101101_01111101 : OUT <= 1;  //173 / 125 = 1
    16'b10101101_01111110 : OUT <= 1;  //173 / 126 = 1
    16'b10101101_01111111 : OUT <= 1;  //173 / 127 = 1
    16'b10101101_10000000 : OUT <= 1;  //173 / 128 = 1
    16'b10101101_10000001 : OUT <= 1;  //173 / 129 = 1
    16'b10101101_10000010 : OUT <= 1;  //173 / 130 = 1
    16'b10101101_10000011 : OUT <= 1;  //173 / 131 = 1
    16'b10101101_10000100 : OUT <= 1;  //173 / 132 = 1
    16'b10101101_10000101 : OUT <= 1;  //173 / 133 = 1
    16'b10101101_10000110 : OUT <= 1;  //173 / 134 = 1
    16'b10101101_10000111 : OUT <= 1;  //173 / 135 = 1
    16'b10101101_10001000 : OUT <= 1;  //173 / 136 = 1
    16'b10101101_10001001 : OUT <= 1;  //173 / 137 = 1
    16'b10101101_10001010 : OUT <= 1;  //173 / 138 = 1
    16'b10101101_10001011 : OUT <= 1;  //173 / 139 = 1
    16'b10101101_10001100 : OUT <= 1;  //173 / 140 = 1
    16'b10101101_10001101 : OUT <= 1;  //173 / 141 = 1
    16'b10101101_10001110 : OUT <= 1;  //173 / 142 = 1
    16'b10101101_10001111 : OUT <= 1;  //173 / 143 = 1
    16'b10101101_10010000 : OUT <= 1;  //173 / 144 = 1
    16'b10101101_10010001 : OUT <= 1;  //173 / 145 = 1
    16'b10101101_10010010 : OUT <= 1;  //173 / 146 = 1
    16'b10101101_10010011 : OUT <= 1;  //173 / 147 = 1
    16'b10101101_10010100 : OUT <= 1;  //173 / 148 = 1
    16'b10101101_10010101 : OUT <= 1;  //173 / 149 = 1
    16'b10101101_10010110 : OUT <= 1;  //173 / 150 = 1
    16'b10101101_10010111 : OUT <= 1;  //173 / 151 = 1
    16'b10101101_10011000 : OUT <= 1;  //173 / 152 = 1
    16'b10101101_10011001 : OUT <= 1;  //173 / 153 = 1
    16'b10101101_10011010 : OUT <= 1;  //173 / 154 = 1
    16'b10101101_10011011 : OUT <= 1;  //173 / 155 = 1
    16'b10101101_10011100 : OUT <= 1;  //173 / 156 = 1
    16'b10101101_10011101 : OUT <= 1;  //173 / 157 = 1
    16'b10101101_10011110 : OUT <= 1;  //173 / 158 = 1
    16'b10101101_10011111 : OUT <= 1;  //173 / 159 = 1
    16'b10101101_10100000 : OUT <= 1;  //173 / 160 = 1
    16'b10101101_10100001 : OUT <= 1;  //173 / 161 = 1
    16'b10101101_10100010 : OUT <= 1;  //173 / 162 = 1
    16'b10101101_10100011 : OUT <= 1;  //173 / 163 = 1
    16'b10101101_10100100 : OUT <= 1;  //173 / 164 = 1
    16'b10101101_10100101 : OUT <= 1;  //173 / 165 = 1
    16'b10101101_10100110 : OUT <= 1;  //173 / 166 = 1
    16'b10101101_10100111 : OUT <= 1;  //173 / 167 = 1
    16'b10101101_10101000 : OUT <= 1;  //173 / 168 = 1
    16'b10101101_10101001 : OUT <= 1;  //173 / 169 = 1
    16'b10101101_10101010 : OUT <= 1;  //173 / 170 = 1
    16'b10101101_10101011 : OUT <= 1;  //173 / 171 = 1
    16'b10101101_10101100 : OUT <= 1;  //173 / 172 = 1
    16'b10101101_10101101 : OUT <= 1;  //173 / 173 = 1
    16'b10101101_10101110 : OUT <= 0;  //173 / 174 = 0
    16'b10101101_10101111 : OUT <= 0;  //173 / 175 = 0
    16'b10101101_10110000 : OUT <= 0;  //173 / 176 = 0
    16'b10101101_10110001 : OUT <= 0;  //173 / 177 = 0
    16'b10101101_10110010 : OUT <= 0;  //173 / 178 = 0
    16'b10101101_10110011 : OUT <= 0;  //173 / 179 = 0
    16'b10101101_10110100 : OUT <= 0;  //173 / 180 = 0
    16'b10101101_10110101 : OUT <= 0;  //173 / 181 = 0
    16'b10101101_10110110 : OUT <= 0;  //173 / 182 = 0
    16'b10101101_10110111 : OUT <= 0;  //173 / 183 = 0
    16'b10101101_10111000 : OUT <= 0;  //173 / 184 = 0
    16'b10101101_10111001 : OUT <= 0;  //173 / 185 = 0
    16'b10101101_10111010 : OUT <= 0;  //173 / 186 = 0
    16'b10101101_10111011 : OUT <= 0;  //173 / 187 = 0
    16'b10101101_10111100 : OUT <= 0;  //173 / 188 = 0
    16'b10101101_10111101 : OUT <= 0;  //173 / 189 = 0
    16'b10101101_10111110 : OUT <= 0;  //173 / 190 = 0
    16'b10101101_10111111 : OUT <= 0;  //173 / 191 = 0
    16'b10101101_11000000 : OUT <= 0;  //173 / 192 = 0
    16'b10101101_11000001 : OUT <= 0;  //173 / 193 = 0
    16'b10101101_11000010 : OUT <= 0;  //173 / 194 = 0
    16'b10101101_11000011 : OUT <= 0;  //173 / 195 = 0
    16'b10101101_11000100 : OUT <= 0;  //173 / 196 = 0
    16'b10101101_11000101 : OUT <= 0;  //173 / 197 = 0
    16'b10101101_11000110 : OUT <= 0;  //173 / 198 = 0
    16'b10101101_11000111 : OUT <= 0;  //173 / 199 = 0
    16'b10101101_11001000 : OUT <= 0;  //173 / 200 = 0
    16'b10101101_11001001 : OUT <= 0;  //173 / 201 = 0
    16'b10101101_11001010 : OUT <= 0;  //173 / 202 = 0
    16'b10101101_11001011 : OUT <= 0;  //173 / 203 = 0
    16'b10101101_11001100 : OUT <= 0;  //173 / 204 = 0
    16'b10101101_11001101 : OUT <= 0;  //173 / 205 = 0
    16'b10101101_11001110 : OUT <= 0;  //173 / 206 = 0
    16'b10101101_11001111 : OUT <= 0;  //173 / 207 = 0
    16'b10101101_11010000 : OUT <= 0;  //173 / 208 = 0
    16'b10101101_11010001 : OUT <= 0;  //173 / 209 = 0
    16'b10101101_11010010 : OUT <= 0;  //173 / 210 = 0
    16'b10101101_11010011 : OUT <= 0;  //173 / 211 = 0
    16'b10101101_11010100 : OUT <= 0;  //173 / 212 = 0
    16'b10101101_11010101 : OUT <= 0;  //173 / 213 = 0
    16'b10101101_11010110 : OUT <= 0;  //173 / 214 = 0
    16'b10101101_11010111 : OUT <= 0;  //173 / 215 = 0
    16'b10101101_11011000 : OUT <= 0;  //173 / 216 = 0
    16'b10101101_11011001 : OUT <= 0;  //173 / 217 = 0
    16'b10101101_11011010 : OUT <= 0;  //173 / 218 = 0
    16'b10101101_11011011 : OUT <= 0;  //173 / 219 = 0
    16'b10101101_11011100 : OUT <= 0;  //173 / 220 = 0
    16'b10101101_11011101 : OUT <= 0;  //173 / 221 = 0
    16'b10101101_11011110 : OUT <= 0;  //173 / 222 = 0
    16'b10101101_11011111 : OUT <= 0;  //173 / 223 = 0
    16'b10101101_11100000 : OUT <= 0;  //173 / 224 = 0
    16'b10101101_11100001 : OUT <= 0;  //173 / 225 = 0
    16'b10101101_11100010 : OUT <= 0;  //173 / 226 = 0
    16'b10101101_11100011 : OUT <= 0;  //173 / 227 = 0
    16'b10101101_11100100 : OUT <= 0;  //173 / 228 = 0
    16'b10101101_11100101 : OUT <= 0;  //173 / 229 = 0
    16'b10101101_11100110 : OUT <= 0;  //173 / 230 = 0
    16'b10101101_11100111 : OUT <= 0;  //173 / 231 = 0
    16'b10101101_11101000 : OUT <= 0;  //173 / 232 = 0
    16'b10101101_11101001 : OUT <= 0;  //173 / 233 = 0
    16'b10101101_11101010 : OUT <= 0;  //173 / 234 = 0
    16'b10101101_11101011 : OUT <= 0;  //173 / 235 = 0
    16'b10101101_11101100 : OUT <= 0;  //173 / 236 = 0
    16'b10101101_11101101 : OUT <= 0;  //173 / 237 = 0
    16'b10101101_11101110 : OUT <= 0;  //173 / 238 = 0
    16'b10101101_11101111 : OUT <= 0;  //173 / 239 = 0
    16'b10101101_11110000 : OUT <= 0;  //173 / 240 = 0
    16'b10101101_11110001 : OUT <= 0;  //173 / 241 = 0
    16'b10101101_11110010 : OUT <= 0;  //173 / 242 = 0
    16'b10101101_11110011 : OUT <= 0;  //173 / 243 = 0
    16'b10101101_11110100 : OUT <= 0;  //173 / 244 = 0
    16'b10101101_11110101 : OUT <= 0;  //173 / 245 = 0
    16'b10101101_11110110 : OUT <= 0;  //173 / 246 = 0
    16'b10101101_11110111 : OUT <= 0;  //173 / 247 = 0
    16'b10101101_11111000 : OUT <= 0;  //173 / 248 = 0
    16'b10101101_11111001 : OUT <= 0;  //173 / 249 = 0
    16'b10101101_11111010 : OUT <= 0;  //173 / 250 = 0
    16'b10101101_11111011 : OUT <= 0;  //173 / 251 = 0
    16'b10101101_11111100 : OUT <= 0;  //173 / 252 = 0
    16'b10101101_11111101 : OUT <= 0;  //173 / 253 = 0
    16'b10101101_11111110 : OUT <= 0;  //173 / 254 = 0
    16'b10101101_11111111 : OUT <= 0;  //173 / 255 = 0
    16'b10101110_00000000 : OUT <= 0;  //174 / 0 = 0
    16'b10101110_00000001 : OUT <= 174;  //174 / 1 = 174
    16'b10101110_00000010 : OUT <= 87;  //174 / 2 = 87
    16'b10101110_00000011 : OUT <= 58;  //174 / 3 = 58
    16'b10101110_00000100 : OUT <= 43;  //174 / 4 = 43
    16'b10101110_00000101 : OUT <= 34;  //174 / 5 = 34
    16'b10101110_00000110 : OUT <= 29;  //174 / 6 = 29
    16'b10101110_00000111 : OUT <= 24;  //174 / 7 = 24
    16'b10101110_00001000 : OUT <= 21;  //174 / 8 = 21
    16'b10101110_00001001 : OUT <= 19;  //174 / 9 = 19
    16'b10101110_00001010 : OUT <= 17;  //174 / 10 = 17
    16'b10101110_00001011 : OUT <= 15;  //174 / 11 = 15
    16'b10101110_00001100 : OUT <= 14;  //174 / 12 = 14
    16'b10101110_00001101 : OUT <= 13;  //174 / 13 = 13
    16'b10101110_00001110 : OUT <= 12;  //174 / 14 = 12
    16'b10101110_00001111 : OUT <= 11;  //174 / 15 = 11
    16'b10101110_00010000 : OUT <= 10;  //174 / 16 = 10
    16'b10101110_00010001 : OUT <= 10;  //174 / 17 = 10
    16'b10101110_00010010 : OUT <= 9;  //174 / 18 = 9
    16'b10101110_00010011 : OUT <= 9;  //174 / 19 = 9
    16'b10101110_00010100 : OUT <= 8;  //174 / 20 = 8
    16'b10101110_00010101 : OUT <= 8;  //174 / 21 = 8
    16'b10101110_00010110 : OUT <= 7;  //174 / 22 = 7
    16'b10101110_00010111 : OUT <= 7;  //174 / 23 = 7
    16'b10101110_00011000 : OUT <= 7;  //174 / 24 = 7
    16'b10101110_00011001 : OUT <= 6;  //174 / 25 = 6
    16'b10101110_00011010 : OUT <= 6;  //174 / 26 = 6
    16'b10101110_00011011 : OUT <= 6;  //174 / 27 = 6
    16'b10101110_00011100 : OUT <= 6;  //174 / 28 = 6
    16'b10101110_00011101 : OUT <= 6;  //174 / 29 = 6
    16'b10101110_00011110 : OUT <= 5;  //174 / 30 = 5
    16'b10101110_00011111 : OUT <= 5;  //174 / 31 = 5
    16'b10101110_00100000 : OUT <= 5;  //174 / 32 = 5
    16'b10101110_00100001 : OUT <= 5;  //174 / 33 = 5
    16'b10101110_00100010 : OUT <= 5;  //174 / 34 = 5
    16'b10101110_00100011 : OUT <= 4;  //174 / 35 = 4
    16'b10101110_00100100 : OUT <= 4;  //174 / 36 = 4
    16'b10101110_00100101 : OUT <= 4;  //174 / 37 = 4
    16'b10101110_00100110 : OUT <= 4;  //174 / 38 = 4
    16'b10101110_00100111 : OUT <= 4;  //174 / 39 = 4
    16'b10101110_00101000 : OUT <= 4;  //174 / 40 = 4
    16'b10101110_00101001 : OUT <= 4;  //174 / 41 = 4
    16'b10101110_00101010 : OUT <= 4;  //174 / 42 = 4
    16'b10101110_00101011 : OUT <= 4;  //174 / 43 = 4
    16'b10101110_00101100 : OUT <= 3;  //174 / 44 = 3
    16'b10101110_00101101 : OUT <= 3;  //174 / 45 = 3
    16'b10101110_00101110 : OUT <= 3;  //174 / 46 = 3
    16'b10101110_00101111 : OUT <= 3;  //174 / 47 = 3
    16'b10101110_00110000 : OUT <= 3;  //174 / 48 = 3
    16'b10101110_00110001 : OUT <= 3;  //174 / 49 = 3
    16'b10101110_00110010 : OUT <= 3;  //174 / 50 = 3
    16'b10101110_00110011 : OUT <= 3;  //174 / 51 = 3
    16'b10101110_00110100 : OUT <= 3;  //174 / 52 = 3
    16'b10101110_00110101 : OUT <= 3;  //174 / 53 = 3
    16'b10101110_00110110 : OUT <= 3;  //174 / 54 = 3
    16'b10101110_00110111 : OUT <= 3;  //174 / 55 = 3
    16'b10101110_00111000 : OUT <= 3;  //174 / 56 = 3
    16'b10101110_00111001 : OUT <= 3;  //174 / 57 = 3
    16'b10101110_00111010 : OUT <= 3;  //174 / 58 = 3
    16'b10101110_00111011 : OUT <= 2;  //174 / 59 = 2
    16'b10101110_00111100 : OUT <= 2;  //174 / 60 = 2
    16'b10101110_00111101 : OUT <= 2;  //174 / 61 = 2
    16'b10101110_00111110 : OUT <= 2;  //174 / 62 = 2
    16'b10101110_00111111 : OUT <= 2;  //174 / 63 = 2
    16'b10101110_01000000 : OUT <= 2;  //174 / 64 = 2
    16'b10101110_01000001 : OUT <= 2;  //174 / 65 = 2
    16'b10101110_01000010 : OUT <= 2;  //174 / 66 = 2
    16'b10101110_01000011 : OUT <= 2;  //174 / 67 = 2
    16'b10101110_01000100 : OUT <= 2;  //174 / 68 = 2
    16'b10101110_01000101 : OUT <= 2;  //174 / 69 = 2
    16'b10101110_01000110 : OUT <= 2;  //174 / 70 = 2
    16'b10101110_01000111 : OUT <= 2;  //174 / 71 = 2
    16'b10101110_01001000 : OUT <= 2;  //174 / 72 = 2
    16'b10101110_01001001 : OUT <= 2;  //174 / 73 = 2
    16'b10101110_01001010 : OUT <= 2;  //174 / 74 = 2
    16'b10101110_01001011 : OUT <= 2;  //174 / 75 = 2
    16'b10101110_01001100 : OUT <= 2;  //174 / 76 = 2
    16'b10101110_01001101 : OUT <= 2;  //174 / 77 = 2
    16'b10101110_01001110 : OUT <= 2;  //174 / 78 = 2
    16'b10101110_01001111 : OUT <= 2;  //174 / 79 = 2
    16'b10101110_01010000 : OUT <= 2;  //174 / 80 = 2
    16'b10101110_01010001 : OUT <= 2;  //174 / 81 = 2
    16'b10101110_01010010 : OUT <= 2;  //174 / 82 = 2
    16'b10101110_01010011 : OUT <= 2;  //174 / 83 = 2
    16'b10101110_01010100 : OUT <= 2;  //174 / 84 = 2
    16'b10101110_01010101 : OUT <= 2;  //174 / 85 = 2
    16'b10101110_01010110 : OUT <= 2;  //174 / 86 = 2
    16'b10101110_01010111 : OUT <= 2;  //174 / 87 = 2
    16'b10101110_01011000 : OUT <= 1;  //174 / 88 = 1
    16'b10101110_01011001 : OUT <= 1;  //174 / 89 = 1
    16'b10101110_01011010 : OUT <= 1;  //174 / 90 = 1
    16'b10101110_01011011 : OUT <= 1;  //174 / 91 = 1
    16'b10101110_01011100 : OUT <= 1;  //174 / 92 = 1
    16'b10101110_01011101 : OUT <= 1;  //174 / 93 = 1
    16'b10101110_01011110 : OUT <= 1;  //174 / 94 = 1
    16'b10101110_01011111 : OUT <= 1;  //174 / 95 = 1
    16'b10101110_01100000 : OUT <= 1;  //174 / 96 = 1
    16'b10101110_01100001 : OUT <= 1;  //174 / 97 = 1
    16'b10101110_01100010 : OUT <= 1;  //174 / 98 = 1
    16'b10101110_01100011 : OUT <= 1;  //174 / 99 = 1
    16'b10101110_01100100 : OUT <= 1;  //174 / 100 = 1
    16'b10101110_01100101 : OUT <= 1;  //174 / 101 = 1
    16'b10101110_01100110 : OUT <= 1;  //174 / 102 = 1
    16'b10101110_01100111 : OUT <= 1;  //174 / 103 = 1
    16'b10101110_01101000 : OUT <= 1;  //174 / 104 = 1
    16'b10101110_01101001 : OUT <= 1;  //174 / 105 = 1
    16'b10101110_01101010 : OUT <= 1;  //174 / 106 = 1
    16'b10101110_01101011 : OUT <= 1;  //174 / 107 = 1
    16'b10101110_01101100 : OUT <= 1;  //174 / 108 = 1
    16'b10101110_01101101 : OUT <= 1;  //174 / 109 = 1
    16'b10101110_01101110 : OUT <= 1;  //174 / 110 = 1
    16'b10101110_01101111 : OUT <= 1;  //174 / 111 = 1
    16'b10101110_01110000 : OUT <= 1;  //174 / 112 = 1
    16'b10101110_01110001 : OUT <= 1;  //174 / 113 = 1
    16'b10101110_01110010 : OUT <= 1;  //174 / 114 = 1
    16'b10101110_01110011 : OUT <= 1;  //174 / 115 = 1
    16'b10101110_01110100 : OUT <= 1;  //174 / 116 = 1
    16'b10101110_01110101 : OUT <= 1;  //174 / 117 = 1
    16'b10101110_01110110 : OUT <= 1;  //174 / 118 = 1
    16'b10101110_01110111 : OUT <= 1;  //174 / 119 = 1
    16'b10101110_01111000 : OUT <= 1;  //174 / 120 = 1
    16'b10101110_01111001 : OUT <= 1;  //174 / 121 = 1
    16'b10101110_01111010 : OUT <= 1;  //174 / 122 = 1
    16'b10101110_01111011 : OUT <= 1;  //174 / 123 = 1
    16'b10101110_01111100 : OUT <= 1;  //174 / 124 = 1
    16'b10101110_01111101 : OUT <= 1;  //174 / 125 = 1
    16'b10101110_01111110 : OUT <= 1;  //174 / 126 = 1
    16'b10101110_01111111 : OUT <= 1;  //174 / 127 = 1
    16'b10101110_10000000 : OUT <= 1;  //174 / 128 = 1
    16'b10101110_10000001 : OUT <= 1;  //174 / 129 = 1
    16'b10101110_10000010 : OUT <= 1;  //174 / 130 = 1
    16'b10101110_10000011 : OUT <= 1;  //174 / 131 = 1
    16'b10101110_10000100 : OUT <= 1;  //174 / 132 = 1
    16'b10101110_10000101 : OUT <= 1;  //174 / 133 = 1
    16'b10101110_10000110 : OUT <= 1;  //174 / 134 = 1
    16'b10101110_10000111 : OUT <= 1;  //174 / 135 = 1
    16'b10101110_10001000 : OUT <= 1;  //174 / 136 = 1
    16'b10101110_10001001 : OUT <= 1;  //174 / 137 = 1
    16'b10101110_10001010 : OUT <= 1;  //174 / 138 = 1
    16'b10101110_10001011 : OUT <= 1;  //174 / 139 = 1
    16'b10101110_10001100 : OUT <= 1;  //174 / 140 = 1
    16'b10101110_10001101 : OUT <= 1;  //174 / 141 = 1
    16'b10101110_10001110 : OUT <= 1;  //174 / 142 = 1
    16'b10101110_10001111 : OUT <= 1;  //174 / 143 = 1
    16'b10101110_10010000 : OUT <= 1;  //174 / 144 = 1
    16'b10101110_10010001 : OUT <= 1;  //174 / 145 = 1
    16'b10101110_10010010 : OUT <= 1;  //174 / 146 = 1
    16'b10101110_10010011 : OUT <= 1;  //174 / 147 = 1
    16'b10101110_10010100 : OUT <= 1;  //174 / 148 = 1
    16'b10101110_10010101 : OUT <= 1;  //174 / 149 = 1
    16'b10101110_10010110 : OUT <= 1;  //174 / 150 = 1
    16'b10101110_10010111 : OUT <= 1;  //174 / 151 = 1
    16'b10101110_10011000 : OUT <= 1;  //174 / 152 = 1
    16'b10101110_10011001 : OUT <= 1;  //174 / 153 = 1
    16'b10101110_10011010 : OUT <= 1;  //174 / 154 = 1
    16'b10101110_10011011 : OUT <= 1;  //174 / 155 = 1
    16'b10101110_10011100 : OUT <= 1;  //174 / 156 = 1
    16'b10101110_10011101 : OUT <= 1;  //174 / 157 = 1
    16'b10101110_10011110 : OUT <= 1;  //174 / 158 = 1
    16'b10101110_10011111 : OUT <= 1;  //174 / 159 = 1
    16'b10101110_10100000 : OUT <= 1;  //174 / 160 = 1
    16'b10101110_10100001 : OUT <= 1;  //174 / 161 = 1
    16'b10101110_10100010 : OUT <= 1;  //174 / 162 = 1
    16'b10101110_10100011 : OUT <= 1;  //174 / 163 = 1
    16'b10101110_10100100 : OUT <= 1;  //174 / 164 = 1
    16'b10101110_10100101 : OUT <= 1;  //174 / 165 = 1
    16'b10101110_10100110 : OUT <= 1;  //174 / 166 = 1
    16'b10101110_10100111 : OUT <= 1;  //174 / 167 = 1
    16'b10101110_10101000 : OUT <= 1;  //174 / 168 = 1
    16'b10101110_10101001 : OUT <= 1;  //174 / 169 = 1
    16'b10101110_10101010 : OUT <= 1;  //174 / 170 = 1
    16'b10101110_10101011 : OUT <= 1;  //174 / 171 = 1
    16'b10101110_10101100 : OUT <= 1;  //174 / 172 = 1
    16'b10101110_10101101 : OUT <= 1;  //174 / 173 = 1
    16'b10101110_10101110 : OUT <= 1;  //174 / 174 = 1
    16'b10101110_10101111 : OUT <= 0;  //174 / 175 = 0
    16'b10101110_10110000 : OUT <= 0;  //174 / 176 = 0
    16'b10101110_10110001 : OUT <= 0;  //174 / 177 = 0
    16'b10101110_10110010 : OUT <= 0;  //174 / 178 = 0
    16'b10101110_10110011 : OUT <= 0;  //174 / 179 = 0
    16'b10101110_10110100 : OUT <= 0;  //174 / 180 = 0
    16'b10101110_10110101 : OUT <= 0;  //174 / 181 = 0
    16'b10101110_10110110 : OUT <= 0;  //174 / 182 = 0
    16'b10101110_10110111 : OUT <= 0;  //174 / 183 = 0
    16'b10101110_10111000 : OUT <= 0;  //174 / 184 = 0
    16'b10101110_10111001 : OUT <= 0;  //174 / 185 = 0
    16'b10101110_10111010 : OUT <= 0;  //174 / 186 = 0
    16'b10101110_10111011 : OUT <= 0;  //174 / 187 = 0
    16'b10101110_10111100 : OUT <= 0;  //174 / 188 = 0
    16'b10101110_10111101 : OUT <= 0;  //174 / 189 = 0
    16'b10101110_10111110 : OUT <= 0;  //174 / 190 = 0
    16'b10101110_10111111 : OUT <= 0;  //174 / 191 = 0
    16'b10101110_11000000 : OUT <= 0;  //174 / 192 = 0
    16'b10101110_11000001 : OUT <= 0;  //174 / 193 = 0
    16'b10101110_11000010 : OUT <= 0;  //174 / 194 = 0
    16'b10101110_11000011 : OUT <= 0;  //174 / 195 = 0
    16'b10101110_11000100 : OUT <= 0;  //174 / 196 = 0
    16'b10101110_11000101 : OUT <= 0;  //174 / 197 = 0
    16'b10101110_11000110 : OUT <= 0;  //174 / 198 = 0
    16'b10101110_11000111 : OUT <= 0;  //174 / 199 = 0
    16'b10101110_11001000 : OUT <= 0;  //174 / 200 = 0
    16'b10101110_11001001 : OUT <= 0;  //174 / 201 = 0
    16'b10101110_11001010 : OUT <= 0;  //174 / 202 = 0
    16'b10101110_11001011 : OUT <= 0;  //174 / 203 = 0
    16'b10101110_11001100 : OUT <= 0;  //174 / 204 = 0
    16'b10101110_11001101 : OUT <= 0;  //174 / 205 = 0
    16'b10101110_11001110 : OUT <= 0;  //174 / 206 = 0
    16'b10101110_11001111 : OUT <= 0;  //174 / 207 = 0
    16'b10101110_11010000 : OUT <= 0;  //174 / 208 = 0
    16'b10101110_11010001 : OUT <= 0;  //174 / 209 = 0
    16'b10101110_11010010 : OUT <= 0;  //174 / 210 = 0
    16'b10101110_11010011 : OUT <= 0;  //174 / 211 = 0
    16'b10101110_11010100 : OUT <= 0;  //174 / 212 = 0
    16'b10101110_11010101 : OUT <= 0;  //174 / 213 = 0
    16'b10101110_11010110 : OUT <= 0;  //174 / 214 = 0
    16'b10101110_11010111 : OUT <= 0;  //174 / 215 = 0
    16'b10101110_11011000 : OUT <= 0;  //174 / 216 = 0
    16'b10101110_11011001 : OUT <= 0;  //174 / 217 = 0
    16'b10101110_11011010 : OUT <= 0;  //174 / 218 = 0
    16'b10101110_11011011 : OUT <= 0;  //174 / 219 = 0
    16'b10101110_11011100 : OUT <= 0;  //174 / 220 = 0
    16'b10101110_11011101 : OUT <= 0;  //174 / 221 = 0
    16'b10101110_11011110 : OUT <= 0;  //174 / 222 = 0
    16'b10101110_11011111 : OUT <= 0;  //174 / 223 = 0
    16'b10101110_11100000 : OUT <= 0;  //174 / 224 = 0
    16'b10101110_11100001 : OUT <= 0;  //174 / 225 = 0
    16'b10101110_11100010 : OUT <= 0;  //174 / 226 = 0
    16'b10101110_11100011 : OUT <= 0;  //174 / 227 = 0
    16'b10101110_11100100 : OUT <= 0;  //174 / 228 = 0
    16'b10101110_11100101 : OUT <= 0;  //174 / 229 = 0
    16'b10101110_11100110 : OUT <= 0;  //174 / 230 = 0
    16'b10101110_11100111 : OUT <= 0;  //174 / 231 = 0
    16'b10101110_11101000 : OUT <= 0;  //174 / 232 = 0
    16'b10101110_11101001 : OUT <= 0;  //174 / 233 = 0
    16'b10101110_11101010 : OUT <= 0;  //174 / 234 = 0
    16'b10101110_11101011 : OUT <= 0;  //174 / 235 = 0
    16'b10101110_11101100 : OUT <= 0;  //174 / 236 = 0
    16'b10101110_11101101 : OUT <= 0;  //174 / 237 = 0
    16'b10101110_11101110 : OUT <= 0;  //174 / 238 = 0
    16'b10101110_11101111 : OUT <= 0;  //174 / 239 = 0
    16'b10101110_11110000 : OUT <= 0;  //174 / 240 = 0
    16'b10101110_11110001 : OUT <= 0;  //174 / 241 = 0
    16'b10101110_11110010 : OUT <= 0;  //174 / 242 = 0
    16'b10101110_11110011 : OUT <= 0;  //174 / 243 = 0
    16'b10101110_11110100 : OUT <= 0;  //174 / 244 = 0
    16'b10101110_11110101 : OUT <= 0;  //174 / 245 = 0
    16'b10101110_11110110 : OUT <= 0;  //174 / 246 = 0
    16'b10101110_11110111 : OUT <= 0;  //174 / 247 = 0
    16'b10101110_11111000 : OUT <= 0;  //174 / 248 = 0
    16'b10101110_11111001 : OUT <= 0;  //174 / 249 = 0
    16'b10101110_11111010 : OUT <= 0;  //174 / 250 = 0
    16'b10101110_11111011 : OUT <= 0;  //174 / 251 = 0
    16'b10101110_11111100 : OUT <= 0;  //174 / 252 = 0
    16'b10101110_11111101 : OUT <= 0;  //174 / 253 = 0
    16'b10101110_11111110 : OUT <= 0;  //174 / 254 = 0
    16'b10101110_11111111 : OUT <= 0;  //174 / 255 = 0
    16'b10101111_00000000 : OUT <= 0;  //175 / 0 = 0
    16'b10101111_00000001 : OUT <= 175;  //175 / 1 = 175
    16'b10101111_00000010 : OUT <= 87;  //175 / 2 = 87
    16'b10101111_00000011 : OUT <= 58;  //175 / 3 = 58
    16'b10101111_00000100 : OUT <= 43;  //175 / 4 = 43
    16'b10101111_00000101 : OUT <= 35;  //175 / 5 = 35
    16'b10101111_00000110 : OUT <= 29;  //175 / 6 = 29
    16'b10101111_00000111 : OUT <= 25;  //175 / 7 = 25
    16'b10101111_00001000 : OUT <= 21;  //175 / 8 = 21
    16'b10101111_00001001 : OUT <= 19;  //175 / 9 = 19
    16'b10101111_00001010 : OUT <= 17;  //175 / 10 = 17
    16'b10101111_00001011 : OUT <= 15;  //175 / 11 = 15
    16'b10101111_00001100 : OUT <= 14;  //175 / 12 = 14
    16'b10101111_00001101 : OUT <= 13;  //175 / 13 = 13
    16'b10101111_00001110 : OUT <= 12;  //175 / 14 = 12
    16'b10101111_00001111 : OUT <= 11;  //175 / 15 = 11
    16'b10101111_00010000 : OUT <= 10;  //175 / 16 = 10
    16'b10101111_00010001 : OUT <= 10;  //175 / 17 = 10
    16'b10101111_00010010 : OUT <= 9;  //175 / 18 = 9
    16'b10101111_00010011 : OUT <= 9;  //175 / 19 = 9
    16'b10101111_00010100 : OUT <= 8;  //175 / 20 = 8
    16'b10101111_00010101 : OUT <= 8;  //175 / 21 = 8
    16'b10101111_00010110 : OUT <= 7;  //175 / 22 = 7
    16'b10101111_00010111 : OUT <= 7;  //175 / 23 = 7
    16'b10101111_00011000 : OUT <= 7;  //175 / 24 = 7
    16'b10101111_00011001 : OUT <= 7;  //175 / 25 = 7
    16'b10101111_00011010 : OUT <= 6;  //175 / 26 = 6
    16'b10101111_00011011 : OUT <= 6;  //175 / 27 = 6
    16'b10101111_00011100 : OUT <= 6;  //175 / 28 = 6
    16'b10101111_00011101 : OUT <= 6;  //175 / 29 = 6
    16'b10101111_00011110 : OUT <= 5;  //175 / 30 = 5
    16'b10101111_00011111 : OUT <= 5;  //175 / 31 = 5
    16'b10101111_00100000 : OUT <= 5;  //175 / 32 = 5
    16'b10101111_00100001 : OUT <= 5;  //175 / 33 = 5
    16'b10101111_00100010 : OUT <= 5;  //175 / 34 = 5
    16'b10101111_00100011 : OUT <= 5;  //175 / 35 = 5
    16'b10101111_00100100 : OUT <= 4;  //175 / 36 = 4
    16'b10101111_00100101 : OUT <= 4;  //175 / 37 = 4
    16'b10101111_00100110 : OUT <= 4;  //175 / 38 = 4
    16'b10101111_00100111 : OUT <= 4;  //175 / 39 = 4
    16'b10101111_00101000 : OUT <= 4;  //175 / 40 = 4
    16'b10101111_00101001 : OUT <= 4;  //175 / 41 = 4
    16'b10101111_00101010 : OUT <= 4;  //175 / 42 = 4
    16'b10101111_00101011 : OUT <= 4;  //175 / 43 = 4
    16'b10101111_00101100 : OUT <= 3;  //175 / 44 = 3
    16'b10101111_00101101 : OUT <= 3;  //175 / 45 = 3
    16'b10101111_00101110 : OUT <= 3;  //175 / 46 = 3
    16'b10101111_00101111 : OUT <= 3;  //175 / 47 = 3
    16'b10101111_00110000 : OUT <= 3;  //175 / 48 = 3
    16'b10101111_00110001 : OUT <= 3;  //175 / 49 = 3
    16'b10101111_00110010 : OUT <= 3;  //175 / 50 = 3
    16'b10101111_00110011 : OUT <= 3;  //175 / 51 = 3
    16'b10101111_00110100 : OUT <= 3;  //175 / 52 = 3
    16'b10101111_00110101 : OUT <= 3;  //175 / 53 = 3
    16'b10101111_00110110 : OUT <= 3;  //175 / 54 = 3
    16'b10101111_00110111 : OUT <= 3;  //175 / 55 = 3
    16'b10101111_00111000 : OUT <= 3;  //175 / 56 = 3
    16'b10101111_00111001 : OUT <= 3;  //175 / 57 = 3
    16'b10101111_00111010 : OUT <= 3;  //175 / 58 = 3
    16'b10101111_00111011 : OUT <= 2;  //175 / 59 = 2
    16'b10101111_00111100 : OUT <= 2;  //175 / 60 = 2
    16'b10101111_00111101 : OUT <= 2;  //175 / 61 = 2
    16'b10101111_00111110 : OUT <= 2;  //175 / 62 = 2
    16'b10101111_00111111 : OUT <= 2;  //175 / 63 = 2
    16'b10101111_01000000 : OUT <= 2;  //175 / 64 = 2
    16'b10101111_01000001 : OUT <= 2;  //175 / 65 = 2
    16'b10101111_01000010 : OUT <= 2;  //175 / 66 = 2
    16'b10101111_01000011 : OUT <= 2;  //175 / 67 = 2
    16'b10101111_01000100 : OUT <= 2;  //175 / 68 = 2
    16'b10101111_01000101 : OUT <= 2;  //175 / 69 = 2
    16'b10101111_01000110 : OUT <= 2;  //175 / 70 = 2
    16'b10101111_01000111 : OUT <= 2;  //175 / 71 = 2
    16'b10101111_01001000 : OUT <= 2;  //175 / 72 = 2
    16'b10101111_01001001 : OUT <= 2;  //175 / 73 = 2
    16'b10101111_01001010 : OUT <= 2;  //175 / 74 = 2
    16'b10101111_01001011 : OUT <= 2;  //175 / 75 = 2
    16'b10101111_01001100 : OUT <= 2;  //175 / 76 = 2
    16'b10101111_01001101 : OUT <= 2;  //175 / 77 = 2
    16'b10101111_01001110 : OUT <= 2;  //175 / 78 = 2
    16'b10101111_01001111 : OUT <= 2;  //175 / 79 = 2
    16'b10101111_01010000 : OUT <= 2;  //175 / 80 = 2
    16'b10101111_01010001 : OUT <= 2;  //175 / 81 = 2
    16'b10101111_01010010 : OUT <= 2;  //175 / 82 = 2
    16'b10101111_01010011 : OUT <= 2;  //175 / 83 = 2
    16'b10101111_01010100 : OUT <= 2;  //175 / 84 = 2
    16'b10101111_01010101 : OUT <= 2;  //175 / 85 = 2
    16'b10101111_01010110 : OUT <= 2;  //175 / 86 = 2
    16'b10101111_01010111 : OUT <= 2;  //175 / 87 = 2
    16'b10101111_01011000 : OUT <= 1;  //175 / 88 = 1
    16'b10101111_01011001 : OUT <= 1;  //175 / 89 = 1
    16'b10101111_01011010 : OUT <= 1;  //175 / 90 = 1
    16'b10101111_01011011 : OUT <= 1;  //175 / 91 = 1
    16'b10101111_01011100 : OUT <= 1;  //175 / 92 = 1
    16'b10101111_01011101 : OUT <= 1;  //175 / 93 = 1
    16'b10101111_01011110 : OUT <= 1;  //175 / 94 = 1
    16'b10101111_01011111 : OUT <= 1;  //175 / 95 = 1
    16'b10101111_01100000 : OUT <= 1;  //175 / 96 = 1
    16'b10101111_01100001 : OUT <= 1;  //175 / 97 = 1
    16'b10101111_01100010 : OUT <= 1;  //175 / 98 = 1
    16'b10101111_01100011 : OUT <= 1;  //175 / 99 = 1
    16'b10101111_01100100 : OUT <= 1;  //175 / 100 = 1
    16'b10101111_01100101 : OUT <= 1;  //175 / 101 = 1
    16'b10101111_01100110 : OUT <= 1;  //175 / 102 = 1
    16'b10101111_01100111 : OUT <= 1;  //175 / 103 = 1
    16'b10101111_01101000 : OUT <= 1;  //175 / 104 = 1
    16'b10101111_01101001 : OUT <= 1;  //175 / 105 = 1
    16'b10101111_01101010 : OUT <= 1;  //175 / 106 = 1
    16'b10101111_01101011 : OUT <= 1;  //175 / 107 = 1
    16'b10101111_01101100 : OUT <= 1;  //175 / 108 = 1
    16'b10101111_01101101 : OUT <= 1;  //175 / 109 = 1
    16'b10101111_01101110 : OUT <= 1;  //175 / 110 = 1
    16'b10101111_01101111 : OUT <= 1;  //175 / 111 = 1
    16'b10101111_01110000 : OUT <= 1;  //175 / 112 = 1
    16'b10101111_01110001 : OUT <= 1;  //175 / 113 = 1
    16'b10101111_01110010 : OUT <= 1;  //175 / 114 = 1
    16'b10101111_01110011 : OUT <= 1;  //175 / 115 = 1
    16'b10101111_01110100 : OUT <= 1;  //175 / 116 = 1
    16'b10101111_01110101 : OUT <= 1;  //175 / 117 = 1
    16'b10101111_01110110 : OUT <= 1;  //175 / 118 = 1
    16'b10101111_01110111 : OUT <= 1;  //175 / 119 = 1
    16'b10101111_01111000 : OUT <= 1;  //175 / 120 = 1
    16'b10101111_01111001 : OUT <= 1;  //175 / 121 = 1
    16'b10101111_01111010 : OUT <= 1;  //175 / 122 = 1
    16'b10101111_01111011 : OUT <= 1;  //175 / 123 = 1
    16'b10101111_01111100 : OUT <= 1;  //175 / 124 = 1
    16'b10101111_01111101 : OUT <= 1;  //175 / 125 = 1
    16'b10101111_01111110 : OUT <= 1;  //175 / 126 = 1
    16'b10101111_01111111 : OUT <= 1;  //175 / 127 = 1
    16'b10101111_10000000 : OUT <= 1;  //175 / 128 = 1
    16'b10101111_10000001 : OUT <= 1;  //175 / 129 = 1
    16'b10101111_10000010 : OUT <= 1;  //175 / 130 = 1
    16'b10101111_10000011 : OUT <= 1;  //175 / 131 = 1
    16'b10101111_10000100 : OUT <= 1;  //175 / 132 = 1
    16'b10101111_10000101 : OUT <= 1;  //175 / 133 = 1
    16'b10101111_10000110 : OUT <= 1;  //175 / 134 = 1
    16'b10101111_10000111 : OUT <= 1;  //175 / 135 = 1
    16'b10101111_10001000 : OUT <= 1;  //175 / 136 = 1
    16'b10101111_10001001 : OUT <= 1;  //175 / 137 = 1
    16'b10101111_10001010 : OUT <= 1;  //175 / 138 = 1
    16'b10101111_10001011 : OUT <= 1;  //175 / 139 = 1
    16'b10101111_10001100 : OUT <= 1;  //175 / 140 = 1
    16'b10101111_10001101 : OUT <= 1;  //175 / 141 = 1
    16'b10101111_10001110 : OUT <= 1;  //175 / 142 = 1
    16'b10101111_10001111 : OUT <= 1;  //175 / 143 = 1
    16'b10101111_10010000 : OUT <= 1;  //175 / 144 = 1
    16'b10101111_10010001 : OUT <= 1;  //175 / 145 = 1
    16'b10101111_10010010 : OUT <= 1;  //175 / 146 = 1
    16'b10101111_10010011 : OUT <= 1;  //175 / 147 = 1
    16'b10101111_10010100 : OUT <= 1;  //175 / 148 = 1
    16'b10101111_10010101 : OUT <= 1;  //175 / 149 = 1
    16'b10101111_10010110 : OUT <= 1;  //175 / 150 = 1
    16'b10101111_10010111 : OUT <= 1;  //175 / 151 = 1
    16'b10101111_10011000 : OUT <= 1;  //175 / 152 = 1
    16'b10101111_10011001 : OUT <= 1;  //175 / 153 = 1
    16'b10101111_10011010 : OUT <= 1;  //175 / 154 = 1
    16'b10101111_10011011 : OUT <= 1;  //175 / 155 = 1
    16'b10101111_10011100 : OUT <= 1;  //175 / 156 = 1
    16'b10101111_10011101 : OUT <= 1;  //175 / 157 = 1
    16'b10101111_10011110 : OUT <= 1;  //175 / 158 = 1
    16'b10101111_10011111 : OUT <= 1;  //175 / 159 = 1
    16'b10101111_10100000 : OUT <= 1;  //175 / 160 = 1
    16'b10101111_10100001 : OUT <= 1;  //175 / 161 = 1
    16'b10101111_10100010 : OUT <= 1;  //175 / 162 = 1
    16'b10101111_10100011 : OUT <= 1;  //175 / 163 = 1
    16'b10101111_10100100 : OUT <= 1;  //175 / 164 = 1
    16'b10101111_10100101 : OUT <= 1;  //175 / 165 = 1
    16'b10101111_10100110 : OUT <= 1;  //175 / 166 = 1
    16'b10101111_10100111 : OUT <= 1;  //175 / 167 = 1
    16'b10101111_10101000 : OUT <= 1;  //175 / 168 = 1
    16'b10101111_10101001 : OUT <= 1;  //175 / 169 = 1
    16'b10101111_10101010 : OUT <= 1;  //175 / 170 = 1
    16'b10101111_10101011 : OUT <= 1;  //175 / 171 = 1
    16'b10101111_10101100 : OUT <= 1;  //175 / 172 = 1
    16'b10101111_10101101 : OUT <= 1;  //175 / 173 = 1
    16'b10101111_10101110 : OUT <= 1;  //175 / 174 = 1
    16'b10101111_10101111 : OUT <= 1;  //175 / 175 = 1
    16'b10101111_10110000 : OUT <= 0;  //175 / 176 = 0
    16'b10101111_10110001 : OUT <= 0;  //175 / 177 = 0
    16'b10101111_10110010 : OUT <= 0;  //175 / 178 = 0
    16'b10101111_10110011 : OUT <= 0;  //175 / 179 = 0
    16'b10101111_10110100 : OUT <= 0;  //175 / 180 = 0
    16'b10101111_10110101 : OUT <= 0;  //175 / 181 = 0
    16'b10101111_10110110 : OUT <= 0;  //175 / 182 = 0
    16'b10101111_10110111 : OUT <= 0;  //175 / 183 = 0
    16'b10101111_10111000 : OUT <= 0;  //175 / 184 = 0
    16'b10101111_10111001 : OUT <= 0;  //175 / 185 = 0
    16'b10101111_10111010 : OUT <= 0;  //175 / 186 = 0
    16'b10101111_10111011 : OUT <= 0;  //175 / 187 = 0
    16'b10101111_10111100 : OUT <= 0;  //175 / 188 = 0
    16'b10101111_10111101 : OUT <= 0;  //175 / 189 = 0
    16'b10101111_10111110 : OUT <= 0;  //175 / 190 = 0
    16'b10101111_10111111 : OUT <= 0;  //175 / 191 = 0
    16'b10101111_11000000 : OUT <= 0;  //175 / 192 = 0
    16'b10101111_11000001 : OUT <= 0;  //175 / 193 = 0
    16'b10101111_11000010 : OUT <= 0;  //175 / 194 = 0
    16'b10101111_11000011 : OUT <= 0;  //175 / 195 = 0
    16'b10101111_11000100 : OUT <= 0;  //175 / 196 = 0
    16'b10101111_11000101 : OUT <= 0;  //175 / 197 = 0
    16'b10101111_11000110 : OUT <= 0;  //175 / 198 = 0
    16'b10101111_11000111 : OUT <= 0;  //175 / 199 = 0
    16'b10101111_11001000 : OUT <= 0;  //175 / 200 = 0
    16'b10101111_11001001 : OUT <= 0;  //175 / 201 = 0
    16'b10101111_11001010 : OUT <= 0;  //175 / 202 = 0
    16'b10101111_11001011 : OUT <= 0;  //175 / 203 = 0
    16'b10101111_11001100 : OUT <= 0;  //175 / 204 = 0
    16'b10101111_11001101 : OUT <= 0;  //175 / 205 = 0
    16'b10101111_11001110 : OUT <= 0;  //175 / 206 = 0
    16'b10101111_11001111 : OUT <= 0;  //175 / 207 = 0
    16'b10101111_11010000 : OUT <= 0;  //175 / 208 = 0
    16'b10101111_11010001 : OUT <= 0;  //175 / 209 = 0
    16'b10101111_11010010 : OUT <= 0;  //175 / 210 = 0
    16'b10101111_11010011 : OUT <= 0;  //175 / 211 = 0
    16'b10101111_11010100 : OUT <= 0;  //175 / 212 = 0
    16'b10101111_11010101 : OUT <= 0;  //175 / 213 = 0
    16'b10101111_11010110 : OUT <= 0;  //175 / 214 = 0
    16'b10101111_11010111 : OUT <= 0;  //175 / 215 = 0
    16'b10101111_11011000 : OUT <= 0;  //175 / 216 = 0
    16'b10101111_11011001 : OUT <= 0;  //175 / 217 = 0
    16'b10101111_11011010 : OUT <= 0;  //175 / 218 = 0
    16'b10101111_11011011 : OUT <= 0;  //175 / 219 = 0
    16'b10101111_11011100 : OUT <= 0;  //175 / 220 = 0
    16'b10101111_11011101 : OUT <= 0;  //175 / 221 = 0
    16'b10101111_11011110 : OUT <= 0;  //175 / 222 = 0
    16'b10101111_11011111 : OUT <= 0;  //175 / 223 = 0
    16'b10101111_11100000 : OUT <= 0;  //175 / 224 = 0
    16'b10101111_11100001 : OUT <= 0;  //175 / 225 = 0
    16'b10101111_11100010 : OUT <= 0;  //175 / 226 = 0
    16'b10101111_11100011 : OUT <= 0;  //175 / 227 = 0
    16'b10101111_11100100 : OUT <= 0;  //175 / 228 = 0
    16'b10101111_11100101 : OUT <= 0;  //175 / 229 = 0
    16'b10101111_11100110 : OUT <= 0;  //175 / 230 = 0
    16'b10101111_11100111 : OUT <= 0;  //175 / 231 = 0
    16'b10101111_11101000 : OUT <= 0;  //175 / 232 = 0
    16'b10101111_11101001 : OUT <= 0;  //175 / 233 = 0
    16'b10101111_11101010 : OUT <= 0;  //175 / 234 = 0
    16'b10101111_11101011 : OUT <= 0;  //175 / 235 = 0
    16'b10101111_11101100 : OUT <= 0;  //175 / 236 = 0
    16'b10101111_11101101 : OUT <= 0;  //175 / 237 = 0
    16'b10101111_11101110 : OUT <= 0;  //175 / 238 = 0
    16'b10101111_11101111 : OUT <= 0;  //175 / 239 = 0
    16'b10101111_11110000 : OUT <= 0;  //175 / 240 = 0
    16'b10101111_11110001 : OUT <= 0;  //175 / 241 = 0
    16'b10101111_11110010 : OUT <= 0;  //175 / 242 = 0
    16'b10101111_11110011 : OUT <= 0;  //175 / 243 = 0
    16'b10101111_11110100 : OUT <= 0;  //175 / 244 = 0
    16'b10101111_11110101 : OUT <= 0;  //175 / 245 = 0
    16'b10101111_11110110 : OUT <= 0;  //175 / 246 = 0
    16'b10101111_11110111 : OUT <= 0;  //175 / 247 = 0
    16'b10101111_11111000 : OUT <= 0;  //175 / 248 = 0
    16'b10101111_11111001 : OUT <= 0;  //175 / 249 = 0
    16'b10101111_11111010 : OUT <= 0;  //175 / 250 = 0
    16'b10101111_11111011 : OUT <= 0;  //175 / 251 = 0
    16'b10101111_11111100 : OUT <= 0;  //175 / 252 = 0
    16'b10101111_11111101 : OUT <= 0;  //175 / 253 = 0
    16'b10101111_11111110 : OUT <= 0;  //175 / 254 = 0
    16'b10101111_11111111 : OUT <= 0;  //175 / 255 = 0
    16'b10110000_00000000 : OUT <= 0;  //176 / 0 = 0
    16'b10110000_00000001 : OUT <= 176;  //176 / 1 = 176
    16'b10110000_00000010 : OUT <= 88;  //176 / 2 = 88
    16'b10110000_00000011 : OUT <= 58;  //176 / 3 = 58
    16'b10110000_00000100 : OUT <= 44;  //176 / 4 = 44
    16'b10110000_00000101 : OUT <= 35;  //176 / 5 = 35
    16'b10110000_00000110 : OUT <= 29;  //176 / 6 = 29
    16'b10110000_00000111 : OUT <= 25;  //176 / 7 = 25
    16'b10110000_00001000 : OUT <= 22;  //176 / 8 = 22
    16'b10110000_00001001 : OUT <= 19;  //176 / 9 = 19
    16'b10110000_00001010 : OUT <= 17;  //176 / 10 = 17
    16'b10110000_00001011 : OUT <= 16;  //176 / 11 = 16
    16'b10110000_00001100 : OUT <= 14;  //176 / 12 = 14
    16'b10110000_00001101 : OUT <= 13;  //176 / 13 = 13
    16'b10110000_00001110 : OUT <= 12;  //176 / 14 = 12
    16'b10110000_00001111 : OUT <= 11;  //176 / 15 = 11
    16'b10110000_00010000 : OUT <= 11;  //176 / 16 = 11
    16'b10110000_00010001 : OUT <= 10;  //176 / 17 = 10
    16'b10110000_00010010 : OUT <= 9;  //176 / 18 = 9
    16'b10110000_00010011 : OUT <= 9;  //176 / 19 = 9
    16'b10110000_00010100 : OUT <= 8;  //176 / 20 = 8
    16'b10110000_00010101 : OUT <= 8;  //176 / 21 = 8
    16'b10110000_00010110 : OUT <= 8;  //176 / 22 = 8
    16'b10110000_00010111 : OUT <= 7;  //176 / 23 = 7
    16'b10110000_00011000 : OUT <= 7;  //176 / 24 = 7
    16'b10110000_00011001 : OUT <= 7;  //176 / 25 = 7
    16'b10110000_00011010 : OUT <= 6;  //176 / 26 = 6
    16'b10110000_00011011 : OUT <= 6;  //176 / 27 = 6
    16'b10110000_00011100 : OUT <= 6;  //176 / 28 = 6
    16'b10110000_00011101 : OUT <= 6;  //176 / 29 = 6
    16'b10110000_00011110 : OUT <= 5;  //176 / 30 = 5
    16'b10110000_00011111 : OUT <= 5;  //176 / 31 = 5
    16'b10110000_00100000 : OUT <= 5;  //176 / 32 = 5
    16'b10110000_00100001 : OUT <= 5;  //176 / 33 = 5
    16'b10110000_00100010 : OUT <= 5;  //176 / 34 = 5
    16'b10110000_00100011 : OUT <= 5;  //176 / 35 = 5
    16'b10110000_00100100 : OUT <= 4;  //176 / 36 = 4
    16'b10110000_00100101 : OUT <= 4;  //176 / 37 = 4
    16'b10110000_00100110 : OUT <= 4;  //176 / 38 = 4
    16'b10110000_00100111 : OUT <= 4;  //176 / 39 = 4
    16'b10110000_00101000 : OUT <= 4;  //176 / 40 = 4
    16'b10110000_00101001 : OUT <= 4;  //176 / 41 = 4
    16'b10110000_00101010 : OUT <= 4;  //176 / 42 = 4
    16'b10110000_00101011 : OUT <= 4;  //176 / 43 = 4
    16'b10110000_00101100 : OUT <= 4;  //176 / 44 = 4
    16'b10110000_00101101 : OUT <= 3;  //176 / 45 = 3
    16'b10110000_00101110 : OUT <= 3;  //176 / 46 = 3
    16'b10110000_00101111 : OUT <= 3;  //176 / 47 = 3
    16'b10110000_00110000 : OUT <= 3;  //176 / 48 = 3
    16'b10110000_00110001 : OUT <= 3;  //176 / 49 = 3
    16'b10110000_00110010 : OUT <= 3;  //176 / 50 = 3
    16'b10110000_00110011 : OUT <= 3;  //176 / 51 = 3
    16'b10110000_00110100 : OUT <= 3;  //176 / 52 = 3
    16'b10110000_00110101 : OUT <= 3;  //176 / 53 = 3
    16'b10110000_00110110 : OUT <= 3;  //176 / 54 = 3
    16'b10110000_00110111 : OUT <= 3;  //176 / 55 = 3
    16'b10110000_00111000 : OUT <= 3;  //176 / 56 = 3
    16'b10110000_00111001 : OUT <= 3;  //176 / 57 = 3
    16'b10110000_00111010 : OUT <= 3;  //176 / 58 = 3
    16'b10110000_00111011 : OUT <= 2;  //176 / 59 = 2
    16'b10110000_00111100 : OUT <= 2;  //176 / 60 = 2
    16'b10110000_00111101 : OUT <= 2;  //176 / 61 = 2
    16'b10110000_00111110 : OUT <= 2;  //176 / 62 = 2
    16'b10110000_00111111 : OUT <= 2;  //176 / 63 = 2
    16'b10110000_01000000 : OUT <= 2;  //176 / 64 = 2
    16'b10110000_01000001 : OUT <= 2;  //176 / 65 = 2
    16'b10110000_01000010 : OUT <= 2;  //176 / 66 = 2
    16'b10110000_01000011 : OUT <= 2;  //176 / 67 = 2
    16'b10110000_01000100 : OUT <= 2;  //176 / 68 = 2
    16'b10110000_01000101 : OUT <= 2;  //176 / 69 = 2
    16'b10110000_01000110 : OUT <= 2;  //176 / 70 = 2
    16'b10110000_01000111 : OUT <= 2;  //176 / 71 = 2
    16'b10110000_01001000 : OUT <= 2;  //176 / 72 = 2
    16'b10110000_01001001 : OUT <= 2;  //176 / 73 = 2
    16'b10110000_01001010 : OUT <= 2;  //176 / 74 = 2
    16'b10110000_01001011 : OUT <= 2;  //176 / 75 = 2
    16'b10110000_01001100 : OUT <= 2;  //176 / 76 = 2
    16'b10110000_01001101 : OUT <= 2;  //176 / 77 = 2
    16'b10110000_01001110 : OUT <= 2;  //176 / 78 = 2
    16'b10110000_01001111 : OUT <= 2;  //176 / 79 = 2
    16'b10110000_01010000 : OUT <= 2;  //176 / 80 = 2
    16'b10110000_01010001 : OUT <= 2;  //176 / 81 = 2
    16'b10110000_01010010 : OUT <= 2;  //176 / 82 = 2
    16'b10110000_01010011 : OUT <= 2;  //176 / 83 = 2
    16'b10110000_01010100 : OUT <= 2;  //176 / 84 = 2
    16'b10110000_01010101 : OUT <= 2;  //176 / 85 = 2
    16'b10110000_01010110 : OUT <= 2;  //176 / 86 = 2
    16'b10110000_01010111 : OUT <= 2;  //176 / 87 = 2
    16'b10110000_01011000 : OUT <= 2;  //176 / 88 = 2
    16'b10110000_01011001 : OUT <= 1;  //176 / 89 = 1
    16'b10110000_01011010 : OUT <= 1;  //176 / 90 = 1
    16'b10110000_01011011 : OUT <= 1;  //176 / 91 = 1
    16'b10110000_01011100 : OUT <= 1;  //176 / 92 = 1
    16'b10110000_01011101 : OUT <= 1;  //176 / 93 = 1
    16'b10110000_01011110 : OUT <= 1;  //176 / 94 = 1
    16'b10110000_01011111 : OUT <= 1;  //176 / 95 = 1
    16'b10110000_01100000 : OUT <= 1;  //176 / 96 = 1
    16'b10110000_01100001 : OUT <= 1;  //176 / 97 = 1
    16'b10110000_01100010 : OUT <= 1;  //176 / 98 = 1
    16'b10110000_01100011 : OUT <= 1;  //176 / 99 = 1
    16'b10110000_01100100 : OUT <= 1;  //176 / 100 = 1
    16'b10110000_01100101 : OUT <= 1;  //176 / 101 = 1
    16'b10110000_01100110 : OUT <= 1;  //176 / 102 = 1
    16'b10110000_01100111 : OUT <= 1;  //176 / 103 = 1
    16'b10110000_01101000 : OUT <= 1;  //176 / 104 = 1
    16'b10110000_01101001 : OUT <= 1;  //176 / 105 = 1
    16'b10110000_01101010 : OUT <= 1;  //176 / 106 = 1
    16'b10110000_01101011 : OUT <= 1;  //176 / 107 = 1
    16'b10110000_01101100 : OUT <= 1;  //176 / 108 = 1
    16'b10110000_01101101 : OUT <= 1;  //176 / 109 = 1
    16'b10110000_01101110 : OUT <= 1;  //176 / 110 = 1
    16'b10110000_01101111 : OUT <= 1;  //176 / 111 = 1
    16'b10110000_01110000 : OUT <= 1;  //176 / 112 = 1
    16'b10110000_01110001 : OUT <= 1;  //176 / 113 = 1
    16'b10110000_01110010 : OUT <= 1;  //176 / 114 = 1
    16'b10110000_01110011 : OUT <= 1;  //176 / 115 = 1
    16'b10110000_01110100 : OUT <= 1;  //176 / 116 = 1
    16'b10110000_01110101 : OUT <= 1;  //176 / 117 = 1
    16'b10110000_01110110 : OUT <= 1;  //176 / 118 = 1
    16'b10110000_01110111 : OUT <= 1;  //176 / 119 = 1
    16'b10110000_01111000 : OUT <= 1;  //176 / 120 = 1
    16'b10110000_01111001 : OUT <= 1;  //176 / 121 = 1
    16'b10110000_01111010 : OUT <= 1;  //176 / 122 = 1
    16'b10110000_01111011 : OUT <= 1;  //176 / 123 = 1
    16'b10110000_01111100 : OUT <= 1;  //176 / 124 = 1
    16'b10110000_01111101 : OUT <= 1;  //176 / 125 = 1
    16'b10110000_01111110 : OUT <= 1;  //176 / 126 = 1
    16'b10110000_01111111 : OUT <= 1;  //176 / 127 = 1
    16'b10110000_10000000 : OUT <= 1;  //176 / 128 = 1
    16'b10110000_10000001 : OUT <= 1;  //176 / 129 = 1
    16'b10110000_10000010 : OUT <= 1;  //176 / 130 = 1
    16'b10110000_10000011 : OUT <= 1;  //176 / 131 = 1
    16'b10110000_10000100 : OUT <= 1;  //176 / 132 = 1
    16'b10110000_10000101 : OUT <= 1;  //176 / 133 = 1
    16'b10110000_10000110 : OUT <= 1;  //176 / 134 = 1
    16'b10110000_10000111 : OUT <= 1;  //176 / 135 = 1
    16'b10110000_10001000 : OUT <= 1;  //176 / 136 = 1
    16'b10110000_10001001 : OUT <= 1;  //176 / 137 = 1
    16'b10110000_10001010 : OUT <= 1;  //176 / 138 = 1
    16'b10110000_10001011 : OUT <= 1;  //176 / 139 = 1
    16'b10110000_10001100 : OUT <= 1;  //176 / 140 = 1
    16'b10110000_10001101 : OUT <= 1;  //176 / 141 = 1
    16'b10110000_10001110 : OUT <= 1;  //176 / 142 = 1
    16'b10110000_10001111 : OUT <= 1;  //176 / 143 = 1
    16'b10110000_10010000 : OUT <= 1;  //176 / 144 = 1
    16'b10110000_10010001 : OUT <= 1;  //176 / 145 = 1
    16'b10110000_10010010 : OUT <= 1;  //176 / 146 = 1
    16'b10110000_10010011 : OUT <= 1;  //176 / 147 = 1
    16'b10110000_10010100 : OUT <= 1;  //176 / 148 = 1
    16'b10110000_10010101 : OUT <= 1;  //176 / 149 = 1
    16'b10110000_10010110 : OUT <= 1;  //176 / 150 = 1
    16'b10110000_10010111 : OUT <= 1;  //176 / 151 = 1
    16'b10110000_10011000 : OUT <= 1;  //176 / 152 = 1
    16'b10110000_10011001 : OUT <= 1;  //176 / 153 = 1
    16'b10110000_10011010 : OUT <= 1;  //176 / 154 = 1
    16'b10110000_10011011 : OUT <= 1;  //176 / 155 = 1
    16'b10110000_10011100 : OUT <= 1;  //176 / 156 = 1
    16'b10110000_10011101 : OUT <= 1;  //176 / 157 = 1
    16'b10110000_10011110 : OUT <= 1;  //176 / 158 = 1
    16'b10110000_10011111 : OUT <= 1;  //176 / 159 = 1
    16'b10110000_10100000 : OUT <= 1;  //176 / 160 = 1
    16'b10110000_10100001 : OUT <= 1;  //176 / 161 = 1
    16'b10110000_10100010 : OUT <= 1;  //176 / 162 = 1
    16'b10110000_10100011 : OUT <= 1;  //176 / 163 = 1
    16'b10110000_10100100 : OUT <= 1;  //176 / 164 = 1
    16'b10110000_10100101 : OUT <= 1;  //176 / 165 = 1
    16'b10110000_10100110 : OUT <= 1;  //176 / 166 = 1
    16'b10110000_10100111 : OUT <= 1;  //176 / 167 = 1
    16'b10110000_10101000 : OUT <= 1;  //176 / 168 = 1
    16'b10110000_10101001 : OUT <= 1;  //176 / 169 = 1
    16'b10110000_10101010 : OUT <= 1;  //176 / 170 = 1
    16'b10110000_10101011 : OUT <= 1;  //176 / 171 = 1
    16'b10110000_10101100 : OUT <= 1;  //176 / 172 = 1
    16'b10110000_10101101 : OUT <= 1;  //176 / 173 = 1
    16'b10110000_10101110 : OUT <= 1;  //176 / 174 = 1
    16'b10110000_10101111 : OUT <= 1;  //176 / 175 = 1
    16'b10110000_10110000 : OUT <= 1;  //176 / 176 = 1
    16'b10110000_10110001 : OUT <= 0;  //176 / 177 = 0
    16'b10110000_10110010 : OUT <= 0;  //176 / 178 = 0
    16'b10110000_10110011 : OUT <= 0;  //176 / 179 = 0
    16'b10110000_10110100 : OUT <= 0;  //176 / 180 = 0
    16'b10110000_10110101 : OUT <= 0;  //176 / 181 = 0
    16'b10110000_10110110 : OUT <= 0;  //176 / 182 = 0
    16'b10110000_10110111 : OUT <= 0;  //176 / 183 = 0
    16'b10110000_10111000 : OUT <= 0;  //176 / 184 = 0
    16'b10110000_10111001 : OUT <= 0;  //176 / 185 = 0
    16'b10110000_10111010 : OUT <= 0;  //176 / 186 = 0
    16'b10110000_10111011 : OUT <= 0;  //176 / 187 = 0
    16'b10110000_10111100 : OUT <= 0;  //176 / 188 = 0
    16'b10110000_10111101 : OUT <= 0;  //176 / 189 = 0
    16'b10110000_10111110 : OUT <= 0;  //176 / 190 = 0
    16'b10110000_10111111 : OUT <= 0;  //176 / 191 = 0
    16'b10110000_11000000 : OUT <= 0;  //176 / 192 = 0
    16'b10110000_11000001 : OUT <= 0;  //176 / 193 = 0
    16'b10110000_11000010 : OUT <= 0;  //176 / 194 = 0
    16'b10110000_11000011 : OUT <= 0;  //176 / 195 = 0
    16'b10110000_11000100 : OUT <= 0;  //176 / 196 = 0
    16'b10110000_11000101 : OUT <= 0;  //176 / 197 = 0
    16'b10110000_11000110 : OUT <= 0;  //176 / 198 = 0
    16'b10110000_11000111 : OUT <= 0;  //176 / 199 = 0
    16'b10110000_11001000 : OUT <= 0;  //176 / 200 = 0
    16'b10110000_11001001 : OUT <= 0;  //176 / 201 = 0
    16'b10110000_11001010 : OUT <= 0;  //176 / 202 = 0
    16'b10110000_11001011 : OUT <= 0;  //176 / 203 = 0
    16'b10110000_11001100 : OUT <= 0;  //176 / 204 = 0
    16'b10110000_11001101 : OUT <= 0;  //176 / 205 = 0
    16'b10110000_11001110 : OUT <= 0;  //176 / 206 = 0
    16'b10110000_11001111 : OUT <= 0;  //176 / 207 = 0
    16'b10110000_11010000 : OUT <= 0;  //176 / 208 = 0
    16'b10110000_11010001 : OUT <= 0;  //176 / 209 = 0
    16'b10110000_11010010 : OUT <= 0;  //176 / 210 = 0
    16'b10110000_11010011 : OUT <= 0;  //176 / 211 = 0
    16'b10110000_11010100 : OUT <= 0;  //176 / 212 = 0
    16'b10110000_11010101 : OUT <= 0;  //176 / 213 = 0
    16'b10110000_11010110 : OUT <= 0;  //176 / 214 = 0
    16'b10110000_11010111 : OUT <= 0;  //176 / 215 = 0
    16'b10110000_11011000 : OUT <= 0;  //176 / 216 = 0
    16'b10110000_11011001 : OUT <= 0;  //176 / 217 = 0
    16'b10110000_11011010 : OUT <= 0;  //176 / 218 = 0
    16'b10110000_11011011 : OUT <= 0;  //176 / 219 = 0
    16'b10110000_11011100 : OUT <= 0;  //176 / 220 = 0
    16'b10110000_11011101 : OUT <= 0;  //176 / 221 = 0
    16'b10110000_11011110 : OUT <= 0;  //176 / 222 = 0
    16'b10110000_11011111 : OUT <= 0;  //176 / 223 = 0
    16'b10110000_11100000 : OUT <= 0;  //176 / 224 = 0
    16'b10110000_11100001 : OUT <= 0;  //176 / 225 = 0
    16'b10110000_11100010 : OUT <= 0;  //176 / 226 = 0
    16'b10110000_11100011 : OUT <= 0;  //176 / 227 = 0
    16'b10110000_11100100 : OUT <= 0;  //176 / 228 = 0
    16'b10110000_11100101 : OUT <= 0;  //176 / 229 = 0
    16'b10110000_11100110 : OUT <= 0;  //176 / 230 = 0
    16'b10110000_11100111 : OUT <= 0;  //176 / 231 = 0
    16'b10110000_11101000 : OUT <= 0;  //176 / 232 = 0
    16'b10110000_11101001 : OUT <= 0;  //176 / 233 = 0
    16'b10110000_11101010 : OUT <= 0;  //176 / 234 = 0
    16'b10110000_11101011 : OUT <= 0;  //176 / 235 = 0
    16'b10110000_11101100 : OUT <= 0;  //176 / 236 = 0
    16'b10110000_11101101 : OUT <= 0;  //176 / 237 = 0
    16'b10110000_11101110 : OUT <= 0;  //176 / 238 = 0
    16'b10110000_11101111 : OUT <= 0;  //176 / 239 = 0
    16'b10110000_11110000 : OUT <= 0;  //176 / 240 = 0
    16'b10110000_11110001 : OUT <= 0;  //176 / 241 = 0
    16'b10110000_11110010 : OUT <= 0;  //176 / 242 = 0
    16'b10110000_11110011 : OUT <= 0;  //176 / 243 = 0
    16'b10110000_11110100 : OUT <= 0;  //176 / 244 = 0
    16'b10110000_11110101 : OUT <= 0;  //176 / 245 = 0
    16'b10110000_11110110 : OUT <= 0;  //176 / 246 = 0
    16'b10110000_11110111 : OUT <= 0;  //176 / 247 = 0
    16'b10110000_11111000 : OUT <= 0;  //176 / 248 = 0
    16'b10110000_11111001 : OUT <= 0;  //176 / 249 = 0
    16'b10110000_11111010 : OUT <= 0;  //176 / 250 = 0
    16'b10110000_11111011 : OUT <= 0;  //176 / 251 = 0
    16'b10110000_11111100 : OUT <= 0;  //176 / 252 = 0
    16'b10110000_11111101 : OUT <= 0;  //176 / 253 = 0
    16'b10110000_11111110 : OUT <= 0;  //176 / 254 = 0
    16'b10110000_11111111 : OUT <= 0;  //176 / 255 = 0
    16'b10110001_00000000 : OUT <= 0;  //177 / 0 = 0
    16'b10110001_00000001 : OUT <= 177;  //177 / 1 = 177
    16'b10110001_00000010 : OUT <= 88;  //177 / 2 = 88
    16'b10110001_00000011 : OUT <= 59;  //177 / 3 = 59
    16'b10110001_00000100 : OUT <= 44;  //177 / 4 = 44
    16'b10110001_00000101 : OUT <= 35;  //177 / 5 = 35
    16'b10110001_00000110 : OUT <= 29;  //177 / 6 = 29
    16'b10110001_00000111 : OUT <= 25;  //177 / 7 = 25
    16'b10110001_00001000 : OUT <= 22;  //177 / 8 = 22
    16'b10110001_00001001 : OUT <= 19;  //177 / 9 = 19
    16'b10110001_00001010 : OUT <= 17;  //177 / 10 = 17
    16'b10110001_00001011 : OUT <= 16;  //177 / 11 = 16
    16'b10110001_00001100 : OUT <= 14;  //177 / 12 = 14
    16'b10110001_00001101 : OUT <= 13;  //177 / 13 = 13
    16'b10110001_00001110 : OUT <= 12;  //177 / 14 = 12
    16'b10110001_00001111 : OUT <= 11;  //177 / 15 = 11
    16'b10110001_00010000 : OUT <= 11;  //177 / 16 = 11
    16'b10110001_00010001 : OUT <= 10;  //177 / 17 = 10
    16'b10110001_00010010 : OUT <= 9;  //177 / 18 = 9
    16'b10110001_00010011 : OUT <= 9;  //177 / 19 = 9
    16'b10110001_00010100 : OUT <= 8;  //177 / 20 = 8
    16'b10110001_00010101 : OUT <= 8;  //177 / 21 = 8
    16'b10110001_00010110 : OUT <= 8;  //177 / 22 = 8
    16'b10110001_00010111 : OUT <= 7;  //177 / 23 = 7
    16'b10110001_00011000 : OUT <= 7;  //177 / 24 = 7
    16'b10110001_00011001 : OUT <= 7;  //177 / 25 = 7
    16'b10110001_00011010 : OUT <= 6;  //177 / 26 = 6
    16'b10110001_00011011 : OUT <= 6;  //177 / 27 = 6
    16'b10110001_00011100 : OUT <= 6;  //177 / 28 = 6
    16'b10110001_00011101 : OUT <= 6;  //177 / 29 = 6
    16'b10110001_00011110 : OUT <= 5;  //177 / 30 = 5
    16'b10110001_00011111 : OUT <= 5;  //177 / 31 = 5
    16'b10110001_00100000 : OUT <= 5;  //177 / 32 = 5
    16'b10110001_00100001 : OUT <= 5;  //177 / 33 = 5
    16'b10110001_00100010 : OUT <= 5;  //177 / 34 = 5
    16'b10110001_00100011 : OUT <= 5;  //177 / 35 = 5
    16'b10110001_00100100 : OUT <= 4;  //177 / 36 = 4
    16'b10110001_00100101 : OUT <= 4;  //177 / 37 = 4
    16'b10110001_00100110 : OUT <= 4;  //177 / 38 = 4
    16'b10110001_00100111 : OUT <= 4;  //177 / 39 = 4
    16'b10110001_00101000 : OUT <= 4;  //177 / 40 = 4
    16'b10110001_00101001 : OUT <= 4;  //177 / 41 = 4
    16'b10110001_00101010 : OUT <= 4;  //177 / 42 = 4
    16'b10110001_00101011 : OUT <= 4;  //177 / 43 = 4
    16'b10110001_00101100 : OUT <= 4;  //177 / 44 = 4
    16'b10110001_00101101 : OUT <= 3;  //177 / 45 = 3
    16'b10110001_00101110 : OUT <= 3;  //177 / 46 = 3
    16'b10110001_00101111 : OUT <= 3;  //177 / 47 = 3
    16'b10110001_00110000 : OUT <= 3;  //177 / 48 = 3
    16'b10110001_00110001 : OUT <= 3;  //177 / 49 = 3
    16'b10110001_00110010 : OUT <= 3;  //177 / 50 = 3
    16'b10110001_00110011 : OUT <= 3;  //177 / 51 = 3
    16'b10110001_00110100 : OUT <= 3;  //177 / 52 = 3
    16'b10110001_00110101 : OUT <= 3;  //177 / 53 = 3
    16'b10110001_00110110 : OUT <= 3;  //177 / 54 = 3
    16'b10110001_00110111 : OUT <= 3;  //177 / 55 = 3
    16'b10110001_00111000 : OUT <= 3;  //177 / 56 = 3
    16'b10110001_00111001 : OUT <= 3;  //177 / 57 = 3
    16'b10110001_00111010 : OUT <= 3;  //177 / 58 = 3
    16'b10110001_00111011 : OUT <= 3;  //177 / 59 = 3
    16'b10110001_00111100 : OUT <= 2;  //177 / 60 = 2
    16'b10110001_00111101 : OUT <= 2;  //177 / 61 = 2
    16'b10110001_00111110 : OUT <= 2;  //177 / 62 = 2
    16'b10110001_00111111 : OUT <= 2;  //177 / 63 = 2
    16'b10110001_01000000 : OUT <= 2;  //177 / 64 = 2
    16'b10110001_01000001 : OUT <= 2;  //177 / 65 = 2
    16'b10110001_01000010 : OUT <= 2;  //177 / 66 = 2
    16'b10110001_01000011 : OUT <= 2;  //177 / 67 = 2
    16'b10110001_01000100 : OUT <= 2;  //177 / 68 = 2
    16'b10110001_01000101 : OUT <= 2;  //177 / 69 = 2
    16'b10110001_01000110 : OUT <= 2;  //177 / 70 = 2
    16'b10110001_01000111 : OUT <= 2;  //177 / 71 = 2
    16'b10110001_01001000 : OUT <= 2;  //177 / 72 = 2
    16'b10110001_01001001 : OUT <= 2;  //177 / 73 = 2
    16'b10110001_01001010 : OUT <= 2;  //177 / 74 = 2
    16'b10110001_01001011 : OUT <= 2;  //177 / 75 = 2
    16'b10110001_01001100 : OUT <= 2;  //177 / 76 = 2
    16'b10110001_01001101 : OUT <= 2;  //177 / 77 = 2
    16'b10110001_01001110 : OUT <= 2;  //177 / 78 = 2
    16'b10110001_01001111 : OUT <= 2;  //177 / 79 = 2
    16'b10110001_01010000 : OUT <= 2;  //177 / 80 = 2
    16'b10110001_01010001 : OUT <= 2;  //177 / 81 = 2
    16'b10110001_01010010 : OUT <= 2;  //177 / 82 = 2
    16'b10110001_01010011 : OUT <= 2;  //177 / 83 = 2
    16'b10110001_01010100 : OUT <= 2;  //177 / 84 = 2
    16'b10110001_01010101 : OUT <= 2;  //177 / 85 = 2
    16'b10110001_01010110 : OUT <= 2;  //177 / 86 = 2
    16'b10110001_01010111 : OUT <= 2;  //177 / 87 = 2
    16'b10110001_01011000 : OUT <= 2;  //177 / 88 = 2
    16'b10110001_01011001 : OUT <= 1;  //177 / 89 = 1
    16'b10110001_01011010 : OUT <= 1;  //177 / 90 = 1
    16'b10110001_01011011 : OUT <= 1;  //177 / 91 = 1
    16'b10110001_01011100 : OUT <= 1;  //177 / 92 = 1
    16'b10110001_01011101 : OUT <= 1;  //177 / 93 = 1
    16'b10110001_01011110 : OUT <= 1;  //177 / 94 = 1
    16'b10110001_01011111 : OUT <= 1;  //177 / 95 = 1
    16'b10110001_01100000 : OUT <= 1;  //177 / 96 = 1
    16'b10110001_01100001 : OUT <= 1;  //177 / 97 = 1
    16'b10110001_01100010 : OUT <= 1;  //177 / 98 = 1
    16'b10110001_01100011 : OUT <= 1;  //177 / 99 = 1
    16'b10110001_01100100 : OUT <= 1;  //177 / 100 = 1
    16'b10110001_01100101 : OUT <= 1;  //177 / 101 = 1
    16'b10110001_01100110 : OUT <= 1;  //177 / 102 = 1
    16'b10110001_01100111 : OUT <= 1;  //177 / 103 = 1
    16'b10110001_01101000 : OUT <= 1;  //177 / 104 = 1
    16'b10110001_01101001 : OUT <= 1;  //177 / 105 = 1
    16'b10110001_01101010 : OUT <= 1;  //177 / 106 = 1
    16'b10110001_01101011 : OUT <= 1;  //177 / 107 = 1
    16'b10110001_01101100 : OUT <= 1;  //177 / 108 = 1
    16'b10110001_01101101 : OUT <= 1;  //177 / 109 = 1
    16'b10110001_01101110 : OUT <= 1;  //177 / 110 = 1
    16'b10110001_01101111 : OUT <= 1;  //177 / 111 = 1
    16'b10110001_01110000 : OUT <= 1;  //177 / 112 = 1
    16'b10110001_01110001 : OUT <= 1;  //177 / 113 = 1
    16'b10110001_01110010 : OUT <= 1;  //177 / 114 = 1
    16'b10110001_01110011 : OUT <= 1;  //177 / 115 = 1
    16'b10110001_01110100 : OUT <= 1;  //177 / 116 = 1
    16'b10110001_01110101 : OUT <= 1;  //177 / 117 = 1
    16'b10110001_01110110 : OUT <= 1;  //177 / 118 = 1
    16'b10110001_01110111 : OUT <= 1;  //177 / 119 = 1
    16'b10110001_01111000 : OUT <= 1;  //177 / 120 = 1
    16'b10110001_01111001 : OUT <= 1;  //177 / 121 = 1
    16'b10110001_01111010 : OUT <= 1;  //177 / 122 = 1
    16'b10110001_01111011 : OUT <= 1;  //177 / 123 = 1
    16'b10110001_01111100 : OUT <= 1;  //177 / 124 = 1
    16'b10110001_01111101 : OUT <= 1;  //177 / 125 = 1
    16'b10110001_01111110 : OUT <= 1;  //177 / 126 = 1
    16'b10110001_01111111 : OUT <= 1;  //177 / 127 = 1
    16'b10110001_10000000 : OUT <= 1;  //177 / 128 = 1
    16'b10110001_10000001 : OUT <= 1;  //177 / 129 = 1
    16'b10110001_10000010 : OUT <= 1;  //177 / 130 = 1
    16'b10110001_10000011 : OUT <= 1;  //177 / 131 = 1
    16'b10110001_10000100 : OUT <= 1;  //177 / 132 = 1
    16'b10110001_10000101 : OUT <= 1;  //177 / 133 = 1
    16'b10110001_10000110 : OUT <= 1;  //177 / 134 = 1
    16'b10110001_10000111 : OUT <= 1;  //177 / 135 = 1
    16'b10110001_10001000 : OUT <= 1;  //177 / 136 = 1
    16'b10110001_10001001 : OUT <= 1;  //177 / 137 = 1
    16'b10110001_10001010 : OUT <= 1;  //177 / 138 = 1
    16'b10110001_10001011 : OUT <= 1;  //177 / 139 = 1
    16'b10110001_10001100 : OUT <= 1;  //177 / 140 = 1
    16'b10110001_10001101 : OUT <= 1;  //177 / 141 = 1
    16'b10110001_10001110 : OUT <= 1;  //177 / 142 = 1
    16'b10110001_10001111 : OUT <= 1;  //177 / 143 = 1
    16'b10110001_10010000 : OUT <= 1;  //177 / 144 = 1
    16'b10110001_10010001 : OUT <= 1;  //177 / 145 = 1
    16'b10110001_10010010 : OUT <= 1;  //177 / 146 = 1
    16'b10110001_10010011 : OUT <= 1;  //177 / 147 = 1
    16'b10110001_10010100 : OUT <= 1;  //177 / 148 = 1
    16'b10110001_10010101 : OUT <= 1;  //177 / 149 = 1
    16'b10110001_10010110 : OUT <= 1;  //177 / 150 = 1
    16'b10110001_10010111 : OUT <= 1;  //177 / 151 = 1
    16'b10110001_10011000 : OUT <= 1;  //177 / 152 = 1
    16'b10110001_10011001 : OUT <= 1;  //177 / 153 = 1
    16'b10110001_10011010 : OUT <= 1;  //177 / 154 = 1
    16'b10110001_10011011 : OUT <= 1;  //177 / 155 = 1
    16'b10110001_10011100 : OUT <= 1;  //177 / 156 = 1
    16'b10110001_10011101 : OUT <= 1;  //177 / 157 = 1
    16'b10110001_10011110 : OUT <= 1;  //177 / 158 = 1
    16'b10110001_10011111 : OUT <= 1;  //177 / 159 = 1
    16'b10110001_10100000 : OUT <= 1;  //177 / 160 = 1
    16'b10110001_10100001 : OUT <= 1;  //177 / 161 = 1
    16'b10110001_10100010 : OUT <= 1;  //177 / 162 = 1
    16'b10110001_10100011 : OUT <= 1;  //177 / 163 = 1
    16'b10110001_10100100 : OUT <= 1;  //177 / 164 = 1
    16'b10110001_10100101 : OUT <= 1;  //177 / 165 = 1
    16'b10110001_10100110 : OUT <= 1;  //177 / 166 = 1
    16'b10110001_10100111 : OUT <= 1;  //177 / 167 = 1
    16'b10110001_10101000 : OUT <= 1;  //177 / 168 = 1
    16'b10110001_10101001 : OUT <= 1;  //177 / 169 = 1
    16'b10110001_10101010 : OUT <= 1;  //177 / 170 = 1
    16'b10110001_10101011 : OUT <= 1;  //177 / 171 = 1
    16'b10110001_10101100 : OUT <= 1;  //177 / 172 = 1
    16'b10110001_10101101 : OUT <= 1;  //177 / 173 = 1
    16'b10110001_10101110 : OUT <= 1;  //177 / 174 = 1
    16'b10110001_10101111 : OUT <= 1;  //177 / 175 = 1
    16'b10110001_10110000 : OUT <= 1;  //177 / 176 = 1
    16'b10110001_10110001 : OUT <= 1;  //177 / 177 = 1
    16'b10110001_10110010 : OUT <= 0;  //177 / 178 = 0
    16'b10110001_10110011 : OUT <= 0;  //177 / 179 = 0
    16'b10110001_10110100 : OUT <= 0;  //177 / 180 = 0
    16'b10110001_10110101 : OUT <= 0;  //177 / 181 = 0
    16'b10110001_10110110 : OUT <= 0;  //177 / 182 = 0
    16'b10110001_10110111 : OUT <= 0;  //177 / 183 = 0
    16'b10110001_10111000 : OUT <= 0;  //177 / 184 = 0
    16'b10110001_10111001 : OUT <= 0;  //177 / 185 = 0
    16'b10110001_10111010 : OUT <= 0;  //177 / 186 = 0
    16'b10110001_10111011 : OUT <= 0;  //177 / 187 = 0
    16'b10110001_10111100 : OUT <= 0;  //177 / 188 = 0
    16'b10110001_10111101 : OUT <= 0;  //177 / 189 = 0
    16'b10110001_10111110 : OUT <= 0;  //177 / 190 = 0
    16'b10110001_10111111 : OUT <= 0;  //177 / 191 = 0
    16'b10110001_11000000 : OUT <= 0;  //177 / 192 = 0
    16'b10110001_11000001 : OUT <= 0;  //177 / 193 = 0
    16'b10110001_11000010 : OUT <= 0;  //177 / 194 = 0
    16'b10110001_11000011 : OUT <= 0;  //177 / 195 = 0
    16'b10110001_11000100 : OUT <= 0;  //177 / 196 = 0
    16'b10110001_11000101 : OUT <= 0;  //177 / 197 = 0
    16'b10110001_11000110 : OUT <= 0;  //177 / 198 = 0
    16'b10110001_11000111 : OUT <= 0;  //177 / 199 = 0
    16'b10110001_11001000 : OUT <= 0;  //177 / 200 = 0
    16'b10110001_11001001 : OUT <= 0;  //177 / 201 = 0
    16'b10110001_11001010 : OUT <= 0;  //177 / 202 = 0
    16'b10110001_11001011 : OUT <= 0;  //177 / 203 = 0
    16'b10110001_11001100 : OUT <= 0;  //177 / 204 = 0
    16'b10110001_11001101 : OUT <= 0;  //177 / 205 = 0
    16'b10110001_11001110 : OUT <= 0;  //177 / 206 = 0
    16'b10110001_11001111 : OUT <= 0;  //177 / 207 = 0
    16'b10110001_11010000 : OUT <= 0;  //177 / 208 = 0
    16'b10110001_11010001 : OUT <= 0;  //177 / 209 = 0
    16'b10110001_11010010 : OUT <= 0;  //177 / 210 = 0
    16'b10110001_11010011 : OUT <= 0;  //177 / 211 = 0
    16'b10110001_11010100 : OUT <= 0;  //177 / 212 = 0
    16'b10110001_11010101 : OUT <= 0;  //177 / 213 = 0
    16'b10110001_11010110 : OUT <= 0;  //177 / 214 = 0
    16'b10110001_11010111 : OUT <= 0;  //177 / 215 = 0
    16'b10110001_11011000 : OUT <= 0;  //177 / 216 = 0
    16'b10110001_11011001 : OUT <= 0;  //177 / 217 = 0
    16'b10110001_11011010 : OUT <= 0;  //177 / 218 = 0
    16'b10110001_11011011 : OUT <= 0;  //177 / 219 = 0
    16'b10110001_11011100 : OUT <= 0;  //177 / 220 = 0
    16'b10110001_11011101 : OUT <= 0;  //177 / 221 = 0
    16'b10110001_11011110 : OUT <= 0;  //177 / 222 = 0
    16'b10110001_11011111 : OUT <= 0;  //177 / 223 = 0
    16'b10110001_11100000 : OUT <= 0;  //177 / 224 = 0
    16'b10110001_11100001 : OUT <= 0;  //177 / 225 = 0
    16'b10110001_11100010 : OUT <= 0;  //177 / 226 = 0
    16'b10110001_11100011 : OUT <= 0;  //177 / 227 = 0
    16'b10110001_11100100 : OUT <= 0;  //177 / 228 = 0
    16'b10110001_11100101 : OUT <= 0;  //177 / 229 = 0
    16'b10110001_11100110 : OUT <= 0;  //177 / 230 = 0
    16'b10110001_11100111 : OUT <= 0;  //177 / 231 = 0
    16'b10110001_11101000 : OUT <= 0;  //177 / 232 = 0
    16'b10110001_11101001 : OUT <= 0;  //177 / 233 = 0
    16'b10110001_11101010 : OUT <= 0;  //177 / 234 = 0
    16'b10110001_11101011 : OUT <= 0;  //177 / 235 = 0
    16'b10110001_11101100 : OUT <= 0;  //177 / 236 = 0
    16'b10110001_11101101 : OUT <= 0;  //177 / 237 = 0
    16'b10110001_11101110 : OUT <= 0;  //177 / 238 = 0
    16'b10110001_11101111 : OUT <= 0;  //177 / 239 = 0
    16'b10110001_11110000 : OUT <= 0;  //177 / 240 = 0
    16'b10110001_11110001 : OUT <= 0;  //177 / 241 = 0
    16'b10110001_11110010 : OUT <= 0;  //177 / 242 = 0
    16'b10110001_11110011 : OUT <= 0;  //177 / 243 = 0
    16'b10110001_11110100 : OUT <= 0;  //177 / 244 = 0
    16'b10110001_11110101 : OUT <= 0;  //177 / 245 = 0
    16'b10110001_11110110 : OUT <= 0;  //177 / 246 = 0
    16'b10110001_11110111 : OUT <= 0;  //177 / 247 = 0
    16'b10110001_11111000 : OUT <= 0;  //177 / 248 = 0
    16'b10110001_11111001 : OUT <= 0;  //177 / 249 = 0
    16'b10110001_11111010 : OUT <= 0;  //177 / 250 = 0
    16'b10110001_11111011 : OUT <= 0;  //177 / 251 = 0
    16'b10110001_11111100 : OUT <= 0;  //177 / 252 = 0
    16'b10110001_11111101 : OUT <= 0;  //177 / 253 = 0
    16'b10110001_11111110 : OUT <= 0;  //177 / 254 = 0
    16'b10110001_11111111 : OUT <= 0;  //177 / 255 = 0
    16'b10110010_00000000 : OUT <= 0;  //178 / 0 = 0
    16'b10110010_00000001 : OUT <= 178;  //178 / 1 = 178
    16'b10110010_00000010 : OUT <= 89;  //178 / 2 = 89
    16'b10110010_00000011 : OUT <= 59;  //178 / 3 = 59
    16'b10110010_00000100 : OUT <= 44;  //178 / 4 = 44
    16'b10110010_00000101 : OUT <= 35;  //178 / 5 = 35
    16'b10110010_00000110 : OUT <= 29;  //178 / 6 = 29
    16'b10110010_00000111 : OUT <= 25;  //178 / 7 = 25
    16'b10110010_00001000 : OUT <= 22;  //178 / 8 = 22
    16'b10110010_00001001 : OUT <= 19;  //178 / 9 = 19
    16'b10110010_00001010 : OUT <= 17;  //178 / 10 = 17
    16'b10110010_00001011 : OUT <= 16;  //178 / 11 = 16
    16'b10110010_00001100 : OUT <= 14;  //178 / 12 = 14
    16'b10110010_00001101 : OUT <= 13;  //178 / 13 = 13
    16'b10110010_00001110 : OUT <= 12;  //178 / 14 = 12
    16'b10110010_00001111 : OUT <= 11;  //178 / 15 = 11
    16'b10110010_00010000 : OUT <= 11;  //178 / 16 = 11
    16'b10110010_00010001 : OUT <= 10;  //178 / 17 = 10
    16'b10110010_00010010 : OUT <= 9;  //178 / 18 = 9
    16'b10110010_00010011 : OUT <= 9;  //178 / 19 = 9
    16'b10110010_00010100 : OUT <= 8;  //178 / 20 = 8
    16'b10110010_00010101 : OUT <= 8;  //178 / 21 = 8
    16'b10110010_00010110 : OUT <= 8;  //178 / 22 = 8
    16'b10110010_00010111 : OUT <= 7;  //178 / 23 = 7
    16'b10110010_00011000 : OUT <= 7;  //178 / 24 = 7
    16'b10110010_00011001 : OUT <= 7;  //178 / 25 = 7
    16'b10110010_00011010 : OUT <= 6;  //178 / 26 = 6
    16'b10110010_00011011 : OUT <= 6;  //178 / 27 = 6
    16'b10110010_00011100 : OUT <= 6;  //178 / 28 = 6
    16'b10110010_00011101 : OUT <= 6;  //178 / 29 = 6
    16'b10110010_00011110 : OUT <= 5;  //178 / 30 = 5
    16'b10110010_00011111 : OUT <= 5;  //178 / 31 = 5
    16'b10110010_00100000 : OUT <= 5;  //178 / 32 = 5
    16'b10110010_00100001 : OUT <= 5;  //178 / 33 = 5
    16'b10110010_00100010 : OUT <= 5;  //178 / 34 = 5
    16'b10110010_00100011 : OUT <= 5;  //178 / 35 = 5
    16'b10110010_00100100 : OUT <= 4;  //178 / 36 = 4
    16'b10110010_00100101 : OUT <= 4;  //178 / 37 = 4
    16'b10110010_00100110 : OUT <= 4;  //178 / 38 = 4
    16'b10110010_00100111 : OUT <= 4;  //178 / 39 = 4
    16'b10110010_00101000 : OUT <= 4;  //178 / 40 = 4
    16'b10110010_00101001 : OUT <= 4;  //178 / 41 = 4
    16'b10110010_00101010 : OUT <= 4;  //178 / 42 = 4
    16'b10110010_00101011 : OUT <= 4;  //178 / 43 = 4
    16'b10110010_00101100 : OUT <= 4;  //178 / 44 = 4
    16'b10110010_00101101 : OUT <= 3;  //178 / 45 = 3
    16'b10110010_00101110 : OUT <= 3;  //178 / 46 = 3
    16'b10110010_00101111 : OUT <= 3;  //178 / 47 = 3
    16'b10110010_00110000 : OUT <= 3;  //178 / 48 = 3
    16'b10110010_00110001 : OUT <= 3;  //178 / 49 = 3
    16'b10110010_00110010 : OUT <= 3;  //178 / 50 = 3
    16'b10110010_00110011 : OUT <= 3;  //178 / 51 = 3
    16'b10110010_00110100 : OUT <= 3;  //178 / 52 = 3
    16'b10110010_00110101 : OUT <= 3;  //178 / 53 = 3
    16'b10110010_00110110 : OUT <= 3;  //178 / 54 = 3
    16'b10110010_00110111 : OUT <= 3;  //178 / 55 = 3
    16'b10110010_00111000 : OUT <= 3;  //178 / 56 = 3
    16'b10110010_00111001 : OUT <= 3;  //178 / 57 = 3
    16'b10110010_00111010 : OUT <= 3;  //178 / 58 = 3
    16'b10110010_00111011 : OUT <= 3;  //178 / 59 = 3
    16'b10110010_00111100 : OUT <= 2;  //178 / 60 = 2
    16'b10110010_00111101 : OUT <= 2;  //178 / 61 = 2
    16'b10110010_00111110 : OUT <= 2;  //178 / 62 = 2
    16'b10110010_00111111 : OUT <= 2;  //178 / 63 = 2
    16'b10110010_01000000 : OUT <= 2;  //178 / 64 = 2
    16'b10110010_01000001 : OUT <= 2;  //178 / 65 = 2
    16'b10110010_01000010 : OUT <= 2;  //178 / 66 = 2
    16'b10110010_01000011 : OUT <= 2;  //178 / 67 = 2
    16'b10110010_01000100 : OUT <= 2;  //178 / 68 = 2
    16'b10110010_01000101 : OUT <= 2;  //178 / 69 = 2
    16'b10110010_01000110 : OUT <= 2;  //178 / 70 = 2
    16'b10110010_01000111 : OUT <= 2;  //178 / 71 = 2
    16'b10110010_01001000 : OUT <= 2;  //178 / 72 = 2
    16'b10110010_01001001 : OUT <= 2;  //178 / 73 = 2
    16'b10110010_01001010 : OUT <= 2;  //178 / 74 = 2
    16'b10110010_01001011 : OUT <= 2;  //178 / 75 = 2
    16'b10110010_01001100 : OUT <= 2;  //178 / 76 = 2
    16'b10110010_01001101 : OUT <= 2;  //178 / 77 = 2
    16'b10110010_01001110 : OUT <= 2;  //178 / 78 = 2
    16'b10110010_01001111 : OUT <= 2;  //178 / 79 = 2
    16'b10110010_01010000 : OUT <= 2;  //178 / 80 = 2
    16'b10110010_01010001 : OUT <= 2;  //178 / 81 = 2
    16'b10110010_01010010 : OUT <= 2;  //178 / 82 = 2
    16'b10110010_01010011 : OUT <= 2;  //178 / 83 = 2
    16'b10110010_01010100 : OUT <= 2;  //178 / 84 = 2
    16'b10110010_01010101 : OUT <= 2;  //178 / 85 = 2
    16'b10110010_01010110 : OUT <= 2;  //178 / 86 = 2
    16'b10110010_01010111 : OUT <= 2;  //178 / 87 = 2
    16'b10110010_01011000 : OUT <= 2;  //178 / 88 = 2
    16'b10110010_01011001 : OUT <= 2;  //178 / 89 = 2
    16'b10110010_01011010 : OUT <= 1;  //178 / 90 = 1
    16'b10110010_01011011 : OUT <= 1;  //178 / 91 = 1
    16'b10110010_01011100 : OUT <= 1;  //178 / 92 = 1
    16'b10110010_01011101 : OUT <= 1;  //178 / 93 = 1
    16'b10110010_01011110 : OUT <= 1;  //178 / 94 = 1
    16'b10110010_01011111 : OUT <= 1;  //178 / 95 = 1
    16'b10110010_01100000 : OUT <= 1;  //178 / 96 = 1
    16'b10110010_01100001 : OUT <= 1;  //178 / 97 = 1
    16'b10110010_01100010 : OUT <= 1;  //178 / 98 = 1
    16'b10110010_01100011 : OUT <= 1;  //178 / 99 = 1
    16'b10110010_01100100 : OUT <= 1;  //178 / 100 = 1
    16'b10110010_01100101 : OUT <= 1;  //178 / 101 = 1
    16'b10110010_01100110 : OUT <= 1;  //178 / 102 = 1
    16'b10110010_01100111 : OUT <= 1;  //178 / 103 = 1
    16'b10110010_01101000 : OUT <= 1;  //178 / 104 = 1
    16'b10110010_01101001 : OUT <= 1;  //178 / 105 = 1
    16'b10110010_01101010 : OUT <= 1;  //178 / 106 = 1
    16'b10110010_01101011 : OUT <= 1;  //178 / 107 = 1
    16'b10110010_01101100 : OUT <= 1;  //178 / 108 = 1
    16'b10110010_01101101 : OUT <= 1;  //178 / 109 = 1
    16'b10110010_01101110 : OUT <= 1;  //178 / 110 = 1
    16'b10110010_01101111 : OUT <= 1;  //178 / 111 = 1
    16'b10110010_01110000 : OUT <= 1;  //178 / 112 = 1
    16'b10110010_01110001 : OUT <= 1;  //178 / 113 = 1
    16'b10110010_01110010 : OUT <= 1;  //178 / 114 = 1
    16'b10110010_01110011 : OUT <= 1;  //178 / 115 = 1
    16'b10110010_01110100 : OUT <= 1;  //178 / 116 = 1
    16'b10110010_01110101 : OUT <= 1;  //178 / 117 = 1
    16'b10110010_01110110 : OUT <= 1;  //178 / 118 = 1
    16'b10110010_01110111 : OUT <= 1;  //178 / 119 = 1
    16'b10110010_01111000 : OUT <= 1;  //178 / 120 = 1
    16'b10110010_01111001 : OUT <= 1;  //178 / 121 = 1
    16'b10110010_01111010 : OUT <= 1;  //178 / 122 = 1
    16'b10110010_01111011 : OUT <= 1;  //178 / 123 = 1
    16'b10110010_01111100 : OUT <= 1;  //178 / 124 = 1
    16'b10110010_01111101 : OUT <= 1;  //178 / 125 = 1
    16'b10110010_01111110 : OUT <= 1;  //178 / 126 = 1
    16'b10110010_01111111 : OUT <= 1;  //178 / 127 = 1
    16'b10110010_10000000 : OUT <= 1;  //178 / 128 = 1
    16'b10110010_10000001 : OUT <= 1;  //178 / 129 = 1
    16'b10110010_10000010 : OUT <= 1;  //178 / 130 = 1
    16'b10110010_10000011 : OUT <= 1;  //178 / 131 = 1
    16'b10110010_10000100 : OUT <= 1;  //178 / 132 = 1
    16'b10110010_10000101 : OUT <= 1;  //178 / 133 = 1
    16'b10110010_10000110 : OUT <= 1;  //178 / 134 = 1
    16'b10110010_10000111 : OUT <= 1;  //178 / 135 = 1
    16'b10110010_10001000 : OUT <= 1;  //178 / 136 = 1
    16'b10110010_10001001 : OUT <= 1;  //178 / 137 = 1
    16'b10110010_10001010 : OUT <= 1;  //178 / 138 = 1
    16'b10110010_10001011 : OUT <= 1;  //178 / 139 = 1
    16'b10110010_10001100 : OUT <= 1;  //178 / 140 = 1
    16'b10110010_10001101 : OUT <= 1;  //178 / 141 = 1
    16'b10110010_10001110 : OUT <= 1;  //178 / 142 = 1
    16'b10110010_10001111 : OUT <= 1;  //178 / 143 = 1
    16'b10110010_10010000 : OUT <= 1;  //178 / 144 = 1
    16'b10110010_10010001 : OUT <= 1;  //178 / 145 = 1
    16'b10110010_10010010 : OUT <= 1;  //178 / 146 = 1
    16'b10110010_10010011 : OUT <= 1;  //178 / 147 = 1
    16'b10110010_10010100 : OUT <= 1;  //178 / 148 = 1
    16'b10110010_10010101 : OUT <= 1;  //178 / 149 = 1
    16'b10110010_10010110 : OUT <= 1;  //178 / 150 = 1
    16'b10110010_10010111 : OUT <= 1;  //178 / 151 = 1
    16'b10110010_10011000 : OUT <= 1;  //178 / 152 = 1
    16'b10110010_10011001 : OUT <= 1;  //178 / 153 = 1
    16'b10110010_10011010 : OUT <= 1;  //178 / 154 = 1
    16'b10110010_10011011 : OUT <= 1;  //178 / 155 = 1
    16'b10110010_10011100 : OUT <= 1;  //178 / 156 = 1
    16'b10110010_10011101 : OUT <= 1;  //178 / 157 = 1
    16'b10110010_10011110 : OUT <= 1;  //178 / 158 = 1
    16'b10110010_10011111 : OUT <= 1;  //178 / 159 = 1
    16'b10110010_10100000 : OUT <= 1;  //178 / 160 = 1
    16'b10110010_10100001 : OUT <= 1;  //178 / 161 = 1
    16'b10110010_10100010 : OUT <= 1;  //178 / 162 = 1
    16'b10110010_10100011 : OUT <= 1;  //178 / 163 = 1
    16'b10110010_10100100 : OUT <= 1;  //178 / 164 = 1
    16'b10110010_10100101 : OUT <= 1;  //178 / 165 = 1
    16'b10110010_10100110 : OUT <= 1;  //178 / 166 = 1
    16'b10110010_10100111 : OUT <= 1;  //178 / 167 = 1
    16'b10110010_10101000 : OUT <= 1;  //178 / 168 = 1
    16'b10110010_10101001 : OUT <= 1;  //178 / 169 = 1
    16'b10110010_10101010 : OUT <= 1;  //178 / 170 = 1
    16'b10110010_10101011 : OUT <= 1;  //178 / 171 = 1
    16'b10110010_10101100 : OUT <= 1;  //178 / 172 = 1
    16'b10110010_10101101 : OUT <= 1;  //178 / 173 = 1
    16'b10110010_10101110 : OUT <= 1;  //178 / 174 = 1
    16'b10110010_10101111 : OUT <= 1;  //178 / 175 = 1
    16'b10110010_10110000 : OUT <= 1;  //178 / 176 = 1
    16'b10110010_10110001 : OUT <= 1;  //178 / 177 = 1
    16'b10110010_10110010 : OUT <= 1;  //178 / 178 = 1
    16'b10110010_10110011 : OUT <= 0;  //178 / 179 = 0
    16'b10110010_10110100 : OUT <= 0;  //178 / 180 = 0
    16'b10110010_10110101 : OUT <= 0;  //178 / 181 = 0
    16'b10110010_10110110 : OUT <= 0;  //178 / 182 = 0
    16'b10110010_10110111 : OUT <= 0;  //178 / 183 = 0
    16'b10110010_10111000 : OUT <= 0;  //178 / 184 = 0
    16'b10110010_10111001 : OUT <= 0;  //178 / 185 = 0
    16'b10110010_10111010 : OUT <= 0;  //178 / 186 = 0
    16'b10110010_10111011 : OUT <= 0;  //178 / 187 = 0
    16'b10110010_10111100 : OUT <= 0;  //178 / 188 = 0
    16'b10110010_10111101 : OUT <= 0;  //178 / 189 = 0
    16'b10110010_10111110 : OUT <= 0;  //178 / 190 = 0
    16'b10110010_10111111 : OUT <= 0;  //178 / 191 = 0
    16'b10110010_11000000 : OUT <= 0;  //178 / 192 = 0
    16'b10110010_11000001 : OUT <= 0;  //178 / 193 = 0
    16'b10110010_11000010 : OUT <= 0;  //178 / 194 = 0
    16'b10110010_11000011 : OUT <= 0;  //178 / 195 = 0
    16'b10110010_11000100 : OUT <= 0;  //178 / 196 = 0
    16'b10110010_11000101 : OUT <= 0;  //178 / 197 = 0
    16'b10110010_11000110 : OUT <= 0;  //178 / 198 = 0
    16'b10110010_11000111 : OUT <= 0;  //178 / 199 = 0
    16'b10110010_11001000 : OUT <= 0;  //178 / 200 = 0
    16'b10110010_11001001 : OUT <= 0;  //178 / 201 = 0
    16'b10110010_11001010 : OUT <= 0;  //178 / 202 = 0
    16'b10110010_11001011 : OUT <= 0;  //178 / 203 = 0
    16'b10110010_11001100 : OUT <= 0;  //178 / 204 = 0
    16'b10110010_11001101 : OUT <= 0;  //178 / 205 = 0
    16'b10110010_11001110 : OUT <= 0;  //178 / 206 = 0
    16'b10110010_11001111 : OUT <= 0;  //178 / 207 = 0
    16'b10110010_11010000 : OUT <= 0;  //178 / 208 = 0
    16'b10110010_11010001 : OUT <= 0;  //178 / 209 = 0
    16'b10110010_11010010 : OUT <= 0;  //178 / 210 = 0
    16'b10110010_11010011 : OUT <= 0;  //178 / 211 = 0
    16'b10110010_11010100 : OUT <= 0;  //178 / 212 = 0
    16'b10110010_11010101 : OUT <= 0;  //178 / 213 = 0
    16'b10110010_11010110 : OUT <= 0;  //178 / 214 = 0
    16'b10110010_11010111 : OUT <= 0;  //178 / 215 = 0
    16'b10110010_11011000 : OUT <= 0;  //178 / 216 = 0
    16'b10110010_11011001 : OUT <= 0;  //178 / 217 = 0
    16'b10110010_11011010 : OUT <= 0;  //178 / 218 = 0
    16'b10110010_11011011 : OUT <= 0;  //178 / 219 = 0
    16'b10110010_11011100 : OUT <= 0;  //178 / 220 = 0
    16'b10110010_11011101 : OUT <= 0;  //178 / 221 = 0
    16'b10110010_11011110 : OUT <= 0;  //178 / 222 = 0
    16'b10110010_11011111 : OUT <= 0;  //178 / 223 = 0
    16'b10110010_11100000 : OUT <= 0;  //178 / 224 = 0
    16'b10110010_11100001 : OUT <= 0;  //178 / 225 = 0
    16'b10110010_11100010 : OUT <= 0;  //178 / 226 = 0
    16'b10110010_11100011 : OUT <= 0;  //178 / 227 = 0
    16'b10110010_11100100 : OUT <= 0;  //178 / 228 = 0
    16'b10110010_11100101 : OUT <= 0;  //178 / 229 = 0
    16'b10110010_11100110 : OUT <= 0;  //178 / 230 = 0
    16'b10110010_11100111 : OUT <= 0;  //178 / 231 = 0
    16'b10110010_11101000 : OUT <= 0;  //178 / 232 = 0
    16'b10110010_11101001 : OUT <= 0;  //178 / 233 = 0
    16'b10110010_11101010 : OUT <= 0;  //178 / 234 = 0
    16'b10110010_11101011 : OUT <= 0;  //178 / 235 = 0
    16'b10110010_11101100 : OUT <= 0;  //178 / 236 = 0
    16'b10110010_11101101 : OUT <= 0;  //178 / 237 = 0
    16'b10110010_11101110 : OUT <= 0;  //178 / 238 = 0
    16'b10110010_11101111 : OUT <= 0;  //178 / 239 = 0
    16'b10110010_11110000 : OUT <= 0;  //178 / 240 = 0
    16'b10110010_11110001 : OUT <= 0;  //178 / 241 = 0
    16'b10110010_11110010 : OUT <= 0;  //178 / 242 = 0
    16'b10110010_11110011 : OUT <= 0;  //178 / 243 = 0
    16'b10110010_11110100 : OUT <= 0;  //178 / 244 = 0
    16'b10110010_11110101 : OUT <= 0;  //178 / 245 = 0
    16'b10110010_11110110 : OUT <= 0;  //178 / 246 = 0
    16'b10110010_11110111 : OUT <= 0;  //178 / 247 = 0
    16'b10110010_11111000 : OUT <= 0;  //178 / 248 = 0
    16'b10110010_11111001 : OUT <= 0;  //178 / 249 = 0
    16'b10110010_11111010 : OUT <= 0;  //178 / 250 = 0
    16'b10110010_11111011 : OUT <= 0;  //178 / 251 = 0
    16'b10110010_11111100 : OUT <= 0;  //178 / 252 = 0
    16'b10110010_11111101 : OUT <= 0;  //178 / 253 = 0
    16'b10110010_11111110 : OUT <= 0;  //178 / 254 = 0
    16'b10110010_11111111 : OUT <= 0;  //178 / 255 = 0
    16'b10110011_00000000 : OUT <= 0;  //179 / 0 = 0
    16'b10110011_00000001 : OUT <= 179;  //179 / 1 = 179
    16'b10110011_00000010 : OUT <= 89;  //179 / 2 = 89
    16'b10110011_00000011 : OUT <= 59;  //179 / 3 = 59
    16'b10110011_00000100 : OUT <= 44;  //179 / 4 = 44
    16'b10110011_00000101 : OUT <= 35;  //179 / 5 = 35
    16'b10110011_00000110 : OUT <= 29;  //179 / 6 = 29
    16'b10110011_00000111 : OUT <= 25;  //179 / 7 = 25
    16'b10110011_00001000 : OUT <= 22;  //179 / 8 = 22
    16'b10110011_00001001 : OUT <= 19;  //179 / 9 = 19
    16'b10110011_00001010 : OUT <= 17;  //179 / 10 = 17
    16'b10110011_00001011 : OUT <= 16;  //179 / 11 = 16
    16'b10110011_00001100 : OUT <= 14;  //179 / 12 = 14
    16'b10110011_00001101 : OUT <= 13;  //179 / 13 = 13
    16'b10110011_00001110 : OUT <= 12;  //179 / 14 = 12
    16'b10110011_00001111 : OUT <= 11;  //179 / 15 = 11
    16'b10110011_00010000 : OUT <= 11;  //179 / 16 = 11
    16'b10110011_00010001 : OUT <= 10;  //179 / 17 = 10
    16'b10110011_00010010 : OUT <= 9;  //179 / 18 = 9
    16'b10110011_00010011 : OUT <= 9;  //179 / 19 = 9
    16'b10110011_00010100 : OUT <= 8;  //179 / 20 = 8
    16'b10110011_00010101 : OUT <= 8;  //179 / 21 = 8
    16'b10110011_00010110 : OUT <= 8;  //179 / 22 = 8
    16'b10110011_00010111 : OUT <= 7;  //179 / 23 = 7
    16'b10110011_00011000 : OUT <= 7;  //179 / 24 = 7
    16'b10110011_00011001 : OUT <= 7;  //179 / 25 = 7
    16'b10110011_00011010 : OUT <= 6;  //179 / 26 = 6
    16'b10110011_00011011 : OUT <= 6;  //179 / 27 = 6
    16'b10110011_00011100 : OUT <= 6;  //179 / 28 = 6
    16'b10110011_00011101 : OUT <= 6;  //179 / 29 = 6
    16'b10110011_00011110 : OUT <= 5;  //179 / 30 = 5
    16'b10110011_00011111 : OUT <= 5;  //179 / 31 = 5
    16'b10110011_00100000 : OUT <= 5;  //179 / 32 = 5
    16'b10110011_00100001 : OUT <= 5;  //179 / 33 = 5
    16'b10110011_00100010 : OUT <= 5;  //179 / 34 = 5
    16'b10110011_00100011 : OUT <= 5;  //179 / 35 = 5
    16'b10110011_00100100 : OUT <= 4;  //179 / 36 = 4
    16'b10110011_00100101 : OUT <= 4;  //179 / 37 = 4
    16'b10110011_00100110 : OUT <= 4;  //179 / 38 = 4
    16'b10110011_00100111 : OUT <= 4;  //179 / 39 = 4
    16'b10110011_00101000 : OUT <= 4;  //179 / 40 = 4
    16'b10110011_00101001 : OUT <= 4;  //179 / 41 = 4
    16'b10110011_00101010 : OUT <= 4;  //179 / 42 = 4
    16'b10110011_00101011 : OUT <= 4;  //179 / 43 = 4
    16'b10110011_00101100 : OUT <= 4;  //179 / 44 = 4
    16'b10110011_00101101 : OUT <= 3;  //179 / 45 = 3
    16'b10110011_00101110 : OUT <= 3;  //179 / 46 = 3
    16'b10110011_00101111 : OUT <= 3;  //179 / 47 = 3
    16'b10110011_00110000 : OUT <= 3;  //179 / 48 = 3
    16'b10110011_00110001 : OUT <= 3;  //179 / 49 = 3
    16'b10110011_00110010 : OUT <= 3;  //179 / 50 = 3
    16'b10110011_00110011 : OUT <= 3;  //179 / 51 = 3
    16'b10110011_00110100 : OUT <= 3;  //179 / 52 = 3
    16'b10110011_00110101 : OUT <= 3;  //179 / 53 = 3
    16'b10110011_00110110 : OUT <= 3;  //179 / 54 = 3
    16'b10110011_00110111 : OUT <= 3;  //179 / 55 = 3
    16'b10110011_00111000 : OUT <= 3;  //179 / 56 = 3
    16'b10110011_00111001 : OUT <= 3;  //179 / 57 = 3
    16'b10110011_00111010 : OUT <= 3;  //179 / 58 = 3
    16'b10110011_00111011 : OUT <= 3;  //179 / 59 = 3
    16'b10110011_00111100 : OUT <= 2;  //179 / 60 = 2
    16'b10110011_00111101 : OUT <= 2;  //179 / 61 = 2
    16'b10110011_00111110 : OUT <= 2;  //179 / 62 = 2
    16'b10110011_00111111 : OUT <= 2;  //179 / 63 = 2
    16'b10110011_01000000 : OUT <= 2;  //179 / 64 = 2
    16'b10110011_01000001 : OUT <= 2;  //179 / 65 = 2
    16'b10110011_01000010 : OUT <= 2;  //179 / 66 = 2
    16'b10110011_01000011 : OUT <= 2;  //179 / 67 = 2
    16'b10110011_01000100 : OUT <= 2;  //179 / 68 = 2
    16'b10110011_01000101 : OUT <= 2;  //179 / 69 = 2
    16'b10110011_01000110 : OUT <= 2;  //179 / 70 = 2
    16'b10110011_01000111 : OUT <= 2;  //179 / 71 = 2
    16'b10110011_01001000 : OUT <= 2;  //179 / 72 = 2
    16'b10110011_01001001 : OUT <= 2;  //179 / 73 = 2
    16'b10110011_01001010 : OUT <= 2;  //179 / 74 = 2
    16'b10110011_01001011 : OUT <= 2;  //179 / 75 = 2
    16'b10110011_01001100 : OUT <= 2;  //179 / 76 = 2
    16'b10110011_01001101 : OUT <= 2;  //179 / 77 = 2
    16'b10110011_01001110 : OUT <= 2;  //179 / 78 = 2
    16'b10110011_01001111 : OUT <= 2;  //179 / 79 = 2
    16'b10110011_01010000 : OUT <= 2;  //179 / 80 = 2
    16'b10110011_01010001 : OUT <= 2;  //179 / 81 = 2
    16'b10110011_01010010 : OUT <= 2;  //179 / 82 = 2
    16'b10110011_01010011 : OUT <= 2;  //179 / 83 = 2
    16'b10110011_01010100 : OUT <= 2;  //179 / 84 = 2
    16'b10110011_01010101 : OUT <= 2;  //179 / 85 = 2
    16'b10110011_01010110 : OUT <= 2;  //179 / 86 = 2
    16'b10110011_01010111 : OUT <= 2;  //179 / 87 = 2
    16'b10110011_01011000 : OUT <= 2;  //179 / 88 = 2
    16'b10110011_01011001 : OUT <= 2;  //179 / 89 = 2
    16'b10110011_01011010 : OUT <= 1;  //179 / 90 = 1
    16'b10110011_01011011 : OUT <= 1;  //179 / 91 = 1
    16'b10110011_01011100 : OUT <= 1;  //179 / 92 = 1
    16'b10110011_01011101 : OUT <= 1;  //179 / 93 = 1
    16'b10110011_01011110 : OUT <= 1;  //179 / 94 = 1
    16'b10110011_01011111 : OUT <= 1;  //179 / 95 = 1
    16'b10110011_01100000 : OUT <= 1;  //179 / 96 = 1
    16'b10110011_01100001 : OUT <= 1;  //179 / 97 = 1
    16'b10110011_01100010 : OUT <= 1;  //179 / 98 = 1
    16'b10110011_01100011 : OUT <= 1;  //179 / 99 = 1
    16'b10110011_01100100 : OUT <= 1;  //179 / 100 = 1
    16'b10110011_01100101 : OUT <= 1;  //179 / 101 = 1
    16'b10110011_01100110 : OUT <= 1;  //179 / 102 = 1
    16'b10110011_01100111 : OUT <= 1;  //179 / 103 = 1
    16'b10110011_01101000 : OUT <= 1;  //179 / 104 = 1
    16'b10110011_01101001 : OUT <= 1;  //179 / 105 = 1
    16'b10110011_01101010 : OUT <= 1;  //179 / 106 = 1
    16'b10110011_01101011 : OUT <= 1;  //179 / 107 = 1
    16'b10110011_01101100 : OUT <= 1;  //179 / 108 = 1
    16'b10110011_01101101 : OUT <= 1;  //179 / 109 = 1
    16'b10110011_01101110 : OUT <= 1;  //179 / 110 = 1
    16'b10110011_01101111 : OUT <= 1;  //179 / 111 = 1
    16'b10110011_01110000 : OUT <= 1;  //179 / 112 = 1
    16'b10110011_01110001 : OUT <= 1;  //179 / 113 = 1
    16'b10110011_01110010 : OUT <= 1;  //179 / 114 = 1
    16'b10110011_01110011 : OUT <= 1;  //179 / 115 = 1
    16'b10110011_01110100 : OUT <= 1;  //179 / 116 = 1
    16'b10110011_01110101 : OUT <= 1;  //179 / 117 = 1
    16'b10110011_01110110 : OUT <= 1;  //179 / 118 = 1
    16'b10110011_01110111 : OUT <= 1;  //179 / 119 = 1
    16'b10110011_01111000 : OUT <= 1;  //179 / 120 = 1
    16'b10110011_01111001 : OUT <= 1;  //179 / 121 = 1
    16'b10110011_01111010 : OUT <= 1;  //179 / 122 = 1
    16'b10110011_01111011 : OUT <= 1;  //179 / 123 = 1
    16'b10110011_01111100 : OUT <= 1;  //179 / 124 = 1
    16'b10110011_01111101 : OUT <= 1;  //179 / 125 = 1
    16'b10110011_01111110 : OUT <= 1;  //179 / 126 = 1
    16'b10110011_01111111 : OUT <= 1;  //179 / 127 = 1
    16'b10110011_10000000 : OUT <= 1;  //179 / 128 = 1
    16'b10110011_10000001 : OUT <= 1;  //179 / 129 = 1
    16'b10110011_10000010 : OUT <= 1;  //179 / 130 = 1
    16'b10110011_10000011 : OUT <= 1;  //179 / 131 = 1
    16'b10110011_10000100 : OUT <= 1;  //179 / 132 = 1
    16'b10110011_10000101 : OUT <= 1;  //179 / 133 = 1
    16'b10110011_10000110 : OUT <= 1;  //179 / 134 = 1
    16'b10110011_10000111 : OUT <= 1;  //179 / 135 = 1
    16'b10110011_10001000 : OUT <= 1;  //179 / 136 = 1
    16'b10110011_10001001 : OUT <= 1;  //179 / 137 = 1
    16'b10110011_10001010 : OUT <= 1;  //179 / 138 = 1
    16'b10110011_10001011 : OUT <= 1;  //179 / 139 = 1
    16'b10110011_10001100 : OUT <= 1;  //179 / 140 = 1
    16'b10110011_10001101 : OUT <= 1;  //179 / 141 = 1
    16'b10110011_10001110 : OUT <= 1;  //179 / 142 = 1
    16'b10110011_10001111 : OUT <= 1;  //179 / 143 = 1
    16'b10110011_10010000 : OUT <= 1;  //179 / 144 = 1
    16'b10110011_10010001 : OUT <= 1;  //179 / 145 = 1
    16'b10110011_10010010 : OUT <= 1;  //179 / 146 = 1
    16'b10110011_10010011 : OUT <= 1;  //179 / 147 = 1
    16'b10110011_10010100 : OUT <= 1;  //179 / 148 = 1
    16'b10110011_10010101 : OUT <= 1;  //179 / 149 = 1
    16'b10110011_10010110 : OUT <= 1;  //179 / 150 = 1
    16'b10110011_10010111 : OUT <= 1;  //179 / 151 = 1
    16'b10110011_10011000 : OUT <= 1;  //179 / 152 = 1
    16'b10110011_10011001 : OUT <= 1;  //179 / 153 = 1
    16'b10110011_10011010 : OUT <= 1;  //179 / 154 = 1
    16'b10110011_10011011 : OUT <= 1;  //179 / 155 = 1
    16'b10110011_10011100 : OUT <= 1;  //179 / 156 = 1
    16'b10110011_10011101 : OUT <= 1;  //179 / 157 = 1
    16'b10110011_10011110 : OUT <= 1;  //179 / 158 = 1
    16'b10110011_10011111 : OUT <= 1;  //179 / 159 = 1
    16'b10110011_10100000 : OUT <= 1;  //179 / 160 = 1
    16'b10110011_10100001 : OUT <= 1;  //179 / 161 = 1
    16'b10110011_10100010 : OUT <= 1;  //179 / 162 = 1
    16'b10110011_10100011 : OUT <= 1;  //179 / 163 = 1
    16'b10110011_10100100 : OUT <= 1;  //179 / 164 = 1
    16'b10110011_10100101 : OUT <= 1;  //179 / 165 = 1
    16'b10110011_10100110 : OUT <= 1;  //179 / 166 = 1
    16'b10110011_10100111 : OUT <= 1;  //179 / 167 = 1
    16'b10110011_10101000 : OUT <= 1;  //179 / 168 = 1
    16'b10110011_10101001 : OUT <= 1;  //179 / 169 = 1
    16'b10110011_10101010 : OUT <= 1;  //179 / 170 = 1
    16'b10110011_10101011 : OUT <= 1;  //179 / 171 = 1
    16'b10110011_10101100 : OUT <= 1;  //179 / 172 = 1
    16'b10110011_10101101 : OUT <= 1;  //179 / 173 = 1
    16'b10110011_10101110 : OUT <= 1;  //179 / 174 = 1
    16'b10110011_10101111 : OUT <= 1;  //179 / 175 = 1
    16'b10110011_10110000 : OUT <= 1;  //179 / 176 = 1
    16'b10110011_10110001 : OUT <= 1;  //179 / 177 = 1
    16'b10110011_10110010 : OUT <= 1;  //179 / 178 = 1
    16'b10110011_10110011 : OUT <= 1;  //179 / 179 = 1
    16'b10110011_10110100 : OUT <= 0;  //179 / 180 = 0
    16'b10110011_10110101 : OUT <= 0;  //179 / 181 = 0
    16'b10110011_10110110 : OUT <= 0;  //179 / 182 = 0
    16'b10110011_10110111 : OUT <= 0;  //179 / 183 = 0
    16'b10110011_10111000 : OUT <= 0;  //179 / 184 = 0
    16'b10110011_10111001 : OUT <= 0;  //179 / 185 = 0
    16'b10110011_10111010 : OUT <= 0;  //179 / 186 = 0
    16'b10110011_10111011 : OUT <= 0;  //179 / 187 = 0
    16'b10110011_10111100 : OUT <= 0;  //179 / 188 = 0
    16'b10110011_10111101 : OUT <= 0;  //179 / 189 = 0
    16'b10110011_10111110 : OUT <= 0;  //179 / 190 = 0
    16'b10110011_10111111 : OUT <= 0;  //179 / 191 = 0
    16'b10110011_11000000 : OUT <= 0;  //179 / 192 = 0
    16'b10110011_11000001 : OUT <= 0;  //179 / 193 = 0
    16'b10110011_11000010 : OUT <= 0;  //179 / 194 = 0
    16'b10110011_11000011 : OUT <= 0;  //179 / 195 = 0
    16'b10110011_11000100 : OUT <= 0;  //179 / 196 = 0
    16'b10110011_11000101 : OUT <= 0;  //179 / 197 = 0
    16'b10110011_11000110 : OUT <= 0;  //179 / 198 = 0
    16'b10110011_11000111 : OUT <= 0;  //179 / 199 = 0
    16'b10110011_11001000 : OUT <= 0;  //179 / 200 = 0
    16'b10110011_11001001 : OUT <= 0;  //179 / 201 = 0
    16'b10110011_11001010 : OUT <= 0;  //179 / 202 = 0
    16'b10110011_11001011 : OUT <= 0;  //179 / 203 = 0
    16'b10110011_11001100 : OUT <= 0;  //179 / 204 = 0
    16'b10110011_11001101 : OUT <= 0;  //179 / 205 = 0
    16'b10110011_11001110 : OUT <= 0;  //179 / 206 = 0
    16'b10110011_11001111 : OUT <= 0;  //179 / 207 = 0
    16'b10110011_11010000 : OUT <= 0;  //179 / 208 = 0
    16'b10110011_11010001 : OUT <= 0;  //179 / 209 = 0
    16'b10110011_11010010 : OUT <= 0;  //179 / 210 = 0
    16'b10110011_11010011 : OUT <= 0;  //179 / 211 = 0
    16'b10110011_11010100 : OUT <= 0;  //179 / 212 = 0
    16'b10110011_11010101 : OUT <= 0;  //179 / 213 = 0
    16'b10110011_11010110 : OUT <= 0;  //179 / 214 = 0
    16'b10110011_11010111 : OUT <= 0;  //179 / 215 = 0
    16'b10110011_11011000 : OUT <= 0;  //179 / 216 = 0
    16'b10110011_11011001 : OUT <= 0;  //179 / 217 = 0
    16'b10110011_11011010 : OUT <= 0;  //179 / 218 = 0
    16'b10110011_11011011 : OUT <= 0;  //179 / 219 = 0
    16'b10110011_11011100 : OUT <= 0;  //179 / 220 = 0
    16'b10110011_11011101 : OUT <= 0;  //179 / 221 = 0
    16'b10110011_11011110 : OUT <= 0;  //179 / 222 = 0
    16'b10110011_11011111 : OUT <= 0;  //179 / 223 = 0
    16'b10110011_11100000 : OUT <= 0;  //179 / 224 = 0
    16'b10110011_11100001 : OUT <= 0;  //179 / 225 = 0
    16'b10110011_11100010 : OUT <= 0;  //179 / 226 = 0
    16'b10110011_11100011 : OUT <= 0;  //179 / 227 = 0
    16'b10110011_11100100 : OUT <= 0;  //179 / 228 = 0
    16'b10110011_11100101 : OUT <= 0;  //179 / 229 = 0
    16'b10110011_11100110 : OUT <= 0;  //179 / 230 = 0
    16'b10110011_11100111 : OUT <= 0;  //179 / 231 = 0
    16'b10110011_11101000 : OUT <= 0;  //179 / 232 = 0
    16'b10110011_11101001 : OUT <= 0;  //179 / 233 = 0
    16'b10110011_11101010 : OUT <= 0;  //179 / 234 = 0
    16'b10110011_11101011 : OUT <= 0;  //179 / 235 = 0
    16'b10110011_11101100 : OUT <= 0;  //179 / 236 = 0
    16'b10110011_11101101 : OUT <= 0;  //179 / 237 = 0
    16'b10110011_11101110 : OUT <= 0;  //179 / 238 = 0
    16'b10110011_11101111 : OUT <= 0;  //179 / 239 = 0
    16'b10110011_11110000 : OUT <= 0;  //179 / 240 = 0
    16'b10110011_11110001 : OUT <= 0;  //179 / 241 = 0
    16'b10110011_11110010 : OUT <= 0;  //179 / 242 = 0
    16'b10110011_11110011 : OUT <= 0;  //179 / 243 = 0
    16'b10110011_11110100 : OUT <= 0;  //179 / 244 = 0
    16'b10110011_11110101 : OUT <= 0;  //179 / 245 = 0
    16'b10110011_11110110 : OUT <= 0;  //179 / 246 = 0
    16'b10110011_11110111 : OUT <= 0;  //179 / 247 = 0
    16'b10110011_11111000 : OUT <= 0;  //179 / 248 = 0
    16'b10110011_11111001 : OUT <= 0;  //179 / 249 = 0
    16'b10110011_11111010 : OUT <= 0;  //179 / 250 = 0
    16'b10110011_11111011 : OUT <= 0;  //179 / 251 = 0
    16'b10110011_11111100 : OUT <= 0;  //179 / 252 = 0
    16'b10110011_11111101 : OUT <= 0;  //179 / 253 = 0
    16'b10110011_11111110 : OUT <= 0;  //179 / 254 = 0
    16'b10110011_11111111 : OUT <= 0;  //179 / 255 = 0
    16'b10110100_00000000 : OUT <= 0;  //180 / 0 = 0
    16'b10110100_00000001 : OUT <= 180;  //180 / 1 = 180
    16'b10110100_00000010 : OUT <= 90;  //180 / 2 = 90
    16'b10110100_00000011 : OUT <= 60;  //180 / 3 = 60
    16'b10110100_00000100 : OUT <= 45;  //180 / 4 = 45
    16'b10110100_00000101 : OUT <= 36;  //180 / 5 = 36
    16'b10110100_00000110 : OUT <= 30;  //180 / 6 = 30
    16'b10110100_00000111 : OUT <= 25;  //180 / 7 = 25
    16'b10110100_00001000 : OUT <= 22;  //180 / 8 = 22
    16'b10110100_00001001 : OUT <= 20;  //180 / 9 = 20
    16'b10110100_00001010 : OUT <= 18;  //180 / 10 = 18
    16'b10110100_00001011 : OUT <= 16;  //180 / 11 = 16
    16'b10110100_00001100 : OUT <= 15;  //180 / 12 = 15
    16'b10110100_00001101 : OUT <= 13;  //180 / 13 = 13
    16'b10110100_00001110 : OUT <= 12;  //180 / 14 = 12
    16'b10110100_00001111 : OUT <= 12;  //180 / 15 = 12
    16'b10110100_00010000 : OUT <= 11;  //180 / 16 = 11
    16'b10110100_00010001 : OUT <= 10;  //180 / 17 = 10
    16'b10110100_00010010 : OUT <= 10;  //180 / 18 = 10
    16'b10110100_00010011 : OUT <= 9;  //180 / 19 = 9
    16'b10110100_00010100 : OUT <= 9;  //180 / 20 = 9
    16'b10110100_00010101 : OUT <= 8;  //180 / 21 = 8
    16'b10110100_00010110 : OUT <= 8;  //180 / 22 = 8
    16'b10110100_00010111 : OUT <= 7;  //180 / 23 = 7
    16'b10110100_00011000 : OUT <= 7;  //180 / 24 = 7
    16'b10110100_00011001 : OUT <= 7;  //180 / 25 = 7
    16'b10110100_00011010 : OUT <= 6;  //180 / 26 = 6
    16'b10110100_00011011 : OUT <= 6;  //180 / 27 = 6
    16'b10110100_00011100 : OUT <= 6;  //180 / 28 = 6
    16'b10110100_00011101 : OUT <= 6;  //180 / 29 = 6
    16'b10110100_00011110 : OUT <= 6;  //180 / 30 = 6
    16'b10110100_00011111 : OUT <= 5;  //180 / 31 = 5
    16'b10110100_00100000 : OUT <= 5;  //180 / 32 = 5
    16'b10110100_00100001 : OUT <= 5;  //180 / 33 = 5
    16'b10110100_00100010 : OUT <= 5;  //180 / 34 = 5
    16'b10110100_00100011 : OUT <= 5;  //180 / 35 = 5
    16'b10110100_00100100 : OUT <= 5;  //180 / 36 = 5
    16'b10110100_00100101 : OUT <= 4;  //180 / 37 = 4
    16'b10110100_00100110 : OUT <= 4;  //180 / 38 = 4
    16'b10110100_00100111 : OUT <= 4;  //180 / 39 = 4
    16'b10110100_00101000 : OUT <= 4;  //180 / 40 = 4
    16'b10110100_00101001 : OUT <= 4;  //180 / 41 = 4
    16'b10110100_00101010 : OUT <= 4;  //180 / 42 = 4
    16'b10110100_00101011 : OUT <= 4;  //180 / 43 = 4
    16'b10110100_00101100 : OUT <= 4;  //180 / 44 = 4
    16'b10110100_00101101 : OUT <= 4;  //180 / 45 = 4
    16'b10110100_00101110 : OUT <= 3;  //180 / 46 = 3
    16'b10110100_00101111 : OUT <= 3;  //180 / 47 = 3
    16'b10110100_00110000 : OUT <= 3;  //180 / 48 = 3
    16'b10110100_00110001 : OUT <= 3;  //180 / 49 = 3
    16'b10110100_00110010 : OUT <= 3;  //180 / 50 = 3
    16'b10110100_00110011 : OUT <= 3;  //180 / 51 = 3
    16'b10110100_00110100 : OUT <= 3;  //180 / 52 = 3
    16'b10110100_00110101 : OUT <= 3;  //180 / 53 = 3
    16'b10110100_00110110 : OUT <= 3;  //180 / 54 = 3
    16'b10110100_00110111 : OUT <= 3;  //180 / 55 = 3
    16'b10110100_00111000 : OUT <= 3;  //180 / 56 = 3
    16'b10110100_00111001 : OUT <= 3;  //180 / 57 = 3
    16'b10110100_00111010 : OUT <= 3;  //180 / 58 = 3
    16'b10110100_00111011 : OUT <= 3;  //180 / 59 = 3
    16'b10110100_00111100 : OUT <= 3;  //180 / 60 = 3
    16'b10110100_00111101 : OUT <= 2;  //180 / 61 = 2
    16'b10110100_00111110 : OUT <= 2;  //180 / 62 = 2
    16'b10110100_00111111 : OUT <= 2;  //180 / 63 = 2
    16'b10110100_01000000 : OUT <= 2;  //180 / 64 = 2
    16'b10110100_01000001 : OUT <= 2;  //180 / 65 = 2
    16'b10110100_01000010 : OUT <= 2;  //180 / 66 = 2
    16'b10110100_01000011 : OUT <= 2;  //180 / 67 = 2
    16'b10110100_01000100 : OUT <= 2;  //180 / 68 = 2
    16'b10110100_01000101 : OUT <= 2;  //180 / 69 = 2
    16'b10110100_01000110 : OUT <= 2;  //180 / 70 = 2
    16'b10110100_01000111 : OUT <= 2;  //180 / 71 = 2
    16'b10110100_01001000 : OUT <= 2;  //180 / 72 = 2
    16'b10110100_01001001 : OUT <= 2;  //180 / 73 = 2
    16'b10110100_01001010 : OUT <= 2;  //180 / 74 = 2
    16'b10110100_01001011 : OUT <= 2;  //180 / 75 = 2
    16'b10110100_01001100 : OUT <= 2;  //180 / 76 = 2
    16'b10110100_01001101 : OUT <= 2;  //180 / 77 = 2
    16'b10110100_01001110 : OUT <= 2;  //180 / 78 = 2
    16'b10110100_01001111 : OUT <= 2;  //180 / 79 = 2
    16'b10110100_01010000 : OUT <= 2;  //180 / 80 = 2
    16'b10110100_01010001 : OUT <= 2;  //180 / 81 = 2
    16'b10110100_01010010 : OUT <= 2;  //180 / 82 = 2
    16'b10110100_01010011 : OUT <= 2;  //180 / 83 = 2
    16'b10110100_01010100 : OUT <= 2;  //180 / 84 = 2
    16'b10110100_01010101 : OUT <= 2;  //180 / 85 = 2
    16'b10110100_01010110 : OUT <= 2;  //180 / 86 = 2
    16'b10110100_01010111 : OUT <= 2;  //180 / 87 = 2
    16'b10110100_01011000 : OUT <= 2;  //180 / 88 = 2
    16'b10110100_01011001 : OUT <= 2;  //180 / 89 = 2
    16'b10110100_01011010 : OUT <= 2;  //180 / 90 = 2
    16'b10110100_01011011 : OUT <= 1;  //180 / 91 = 1
    16'b10110100_01011100 : OUT <= 1;  //180 / 92 = 1
    16'b10110100_01011101 : OUT <= 1;  //180 / 93 = 1
    16'b10110100_01011110 : OUT <= 1;  //180 / 94 = 1
    16'b10110100_01011111 : OUT <= 1;  //180 / 95 = 1
    16'b10110100_01100000 : OUT <= 1;  //180 / 96 = 1
    16'b10110100_01100001 : OUT <= 1;  //180 / 97 = 1
    16'b10110100_01100010 : OUT <= 1;  //180 / 98 = 1
    16'b10110100_01100011 : OUT <= 1;  //180 / 99 = 1
    16'b10110100_01100100 : OUT <= 1;  //180 / 100 = 1
    16'b10110100_01100101 : OUT <= 1;  //180 / 101 = 1
    16'b10110100_01100110 : OUT <= 1;  //180 / 102 = 1
    16'b10110100_01100111 : OUT <= 1;  //180 / 103 = 1
    16'b10110100_01101000 : OUT <= 1;  //180 / 104 = 1
    16'b10110100_01101001 : OUT <= 1;  //180 / 105 = 1
    16'b10110100_01101010 : OUT <= 1;  //180 / 106 = 1
    16'b10110100_01101011 : OUT <= 1;  //180 / 107 = 1
    16'b10110100_01101100 : OUT <= 1;  //180 / 108 = 1
    16'b10110100_01101101 : OUT <= 1;  //180 / 109 = 1
    16'b10110100_01101110 : OUT <= 1;  //180 / 110 = 1
    16'b10110100_01101111 : OUT <= 1;  //180 / 111 = 1
    16'b10110100_01110000 : OUT <= 1;  //180 / 112 = 1
    16'b10110100_01110001 : OUT <= 1;  //180 / 113 = 1
    16'b10110100_01110010 : OUT <= 1;  //180 / 114 = 1
    16'b10110100_01110011 : OUT <= 1;  //180 / 115 = 1
    16'b10110100_01110100 : OUT <= 1;  //180 / 116 = 1
    16'b10110100_01110101 : OUT <= 1;  //180 / 117 = 1
    16'b10110100_01110110 : OUT <= 1;  //180 / 118 = 1
    16'b10110100_01110111 : OUT <= 1;  //180 / 119 = 1
    16'b10110100_01111000 : OUT <= 1;  //180 / 120 = 1
    16'b10110100_01111001 : OUT <= 1;  //180 / 121 = 1
    16'b10110100_01111010 : OUT <= 1;  //180 / 122 = 1
    16'b10110100_01111011 : OUT <= 1;  //180 / 123 = 1
    16'b10110100_01111100 : OUT <= 1;  //180 / 124 = 1
    16'b10110100_01111101 : OUT <= 1;  //180 / 125 = 1
    16'b10110100_01111110 : OUT <= 1;  //180 / 126 = 1
    16'b10110100_01111111 : OUT <= 1;  //180 / 127 = 1
    16'b10110100_10000000 : OUT <= 1;  //180 / 128 = 1
    16'b10110100_10000001 : OUT <= 1;  //180 / 129 = 1
    16'b10110100_10000010 : OUT <= 1;  //180 / 130 = 1
    16'b10110100_10000011 : OUT <= 1;  //180 / 131 = 1
    16'b10110100_10000100 : OUT <= 1;  //180 / 132 = 1
    16'b10110100_10000101 : OUT <= 1;  //180 / 133 = 1
    16'b10110100_10000110 : OUT <= 1;  //180 / 134 = 1
    16'b10110100_10000111 : OUT <= 1;  //180 / 135 = 1
    16'b10110100_10001000 : OUT <= 1;  //180 / 136 = 1
    16'b10110100_10001001 : OUT <= 1;  //180 / 137 = 1
    16'b10110100_10001010 : OUT <= 1;  //180 / 138 = 1
    16'b10110100_10001011 : OUT <= 1;  //180 / 139 = 1
    16'b10110100_10001100 : OUT <= 1;  //180 / 140 = 1
    16'b10110100_10001101 : OUT <= 1;  //180 / 141 = 1
    16'b10110100_10001110 : OUT <= 1;  //180 / 142 = 1
    16'b10110100_10001111 : OUT <= 1;  //180 / 143 = 1
    16'b10110100_10010000 : OUT <= 1;  //180 / 144 = 1
    16'b10110100_10010001 : OUT <= 1;  //180 / 145 = 1
    16'b10110100_10010010 : OUT <= 1;  //180 / 146 = 1
    16'b10110100_10010011 : OUT <= 1;  //180 / 147 = 1
    16'b10110100_10010100 : OUT <= 1;  //180 / 148 = 1
    16'b10110100_10010101 : OUT <= 1;  //180 / 149 = 1
    16'b10110100_10010110 : OUT <= 1;  //180 / 150 = 1
    16'b10110100_10010111 : OUT <= 1;  //180 / 151 = 1
    16'b10110100_10011000 : OUT <= 1;  //180 / 152 = 1
    16'b10110100_10011001 : OUT <= 1;  //180 / 153 = 1
    16'b10110100_10011010 : OUT <= 1;  //180 / 154 = 1
    16'b10110100_10011011 : OUT <= 1;  //180 / 155 = 1
    16'b10110100_10011100 : OUT <= 1;  //180 / 156 = 1
    16'b10110100_10011101 : OUT <= 1;  //180 / 157 = 1
    16'b10110100_10011110 : OUT <= 1;  //180 / 158 = 1
    16'b10110100_10011111 : OUT <= 1;  //180 / 159 = 1
    16'b10110100_10100000 : OUT <= 1;  //180 / 160 = 1
    16'b10110100_10100001 : OUT <= 1;  //180 / 161 = 1
    16'b10110100_10100010 : OUT <= 1;  //180 / 162 = 1
    16'b10110100_10100011 : OUT <= 1;  //180 / 163 = 1
    16'b10110100_10100100 : OUT <= 1;  //180 / 164 = 1
    16'b10110100_10100101 : OUT <= 1;  //180 / 165 = 1
    16'b10110100_10100110 : OUT <= 1;  //180 / 166 = 1
    16'b10110100_10100111 : OUT <= 1;  //180 / 167 = 1
    16'b10110100_10101000 : OUT <= 1;  //180 / 168 = 1
    16'b10110100_10101001 : OUT <= 1;  //180 / 169 = 1
    16'b10110100_10101010 : OUT <= 1;  //180 / 170 = 1
    16'b10110100_10101011 : OUT <= 1;  //180 / 171 = 1
    16'b10110100_10101100 : OUT <= 1;  //180 / 172 = 1
    16'b10110100_10101101 : OUT <= 1;  //180 / 173 = 1
    16'b10110100_10101110 : OUT <= 1;  //180 / 174 = 1
    16'b10110100_10101111 : OUT <= 1;  //180 / 175 = 1
    16'b10110100_10110000 : OUT <= 1;  //180 / 176 = 1
    16'b10110100_10110001 : OUT <= 1;  //180 / 177 = 1
    16'b10110100_10110010 : OUT <= 1;  //180 / 178 = 1
    16'b10110100_10110011 : OUT <= 1;  //180 / 179 = 1
    16'b10110100_10110100 : OUT <= 1;  //180 / 180 = 1
    16'b10110100_10110101 : OUT <= 0;  //180 / 181 = 0
    16'b10110100_10110110 : OUT <= 0;  //180 / 182 = 0
    16'b10110100_10110111 : OUT <= 0;  //180 / 183 = 0
    16'b10110100_10111000 : OUT <= 0;  //180 / 184 = 0
    16'b10110100_10111001 : OUT <= 0;  //180 / 185 = 0
    16'b10110100_10111010 : OUT <= 0;  //180 / 186 = 0
    16'b10110100_10111011 : OUT <= 0;  //180 / 187 = 0
    16'b10110100_10111100 : OUT <= 0;  //180 / 188 = 0
    16'b10110100_10111101 : OUT <= 0;  //180 / 189 = 0
    16'b10110100_10111110 : OUT <= 0;  //180 / 190 = 0
    16'b10110100_10111111 : OUT <= 0;  //180 / 191 = 0
    16'b10110100_11000000 : OUT <= 0;  //180 / 192 = 0
    16'b10110100_11000001 : OUT <= 0;  //180 / 193 = 0
    16'b10110100_11000010 : OUT <= 0;  //180 / 194 = 0
    16'b10110100_11000011 : OUT <= 0;  //180 / 195 = 0
    16'b10110100_11000100 : OUT <= 0;  //180 / 196 = 0
    16'b10110100_11000101 : OUT <= 0;  //180 / 197 = 0
    16'b10110100_11000110 : OUT <= 0;  //180 / 198 = 0
    16'b10110100_11000111 : OUT <= 0;  //180 / 199 = 0
    16'b10110100_11001000 : OUT <= 0;  //180 / 200 = 0
    16'b10110100_11001001 : OUT <= 0;  //180 / 201 = 0
    16'b10110100_11001010 : OUT <= 0;  //180 / 202 = 0
    16'b10110100_11001011 : OUT <= 0;  //180 / 203 = 0
    16'b10110100_11001100 : OUT <= 0;  //180 / 204 = 0
    16'b10110100_11001101 : OUT <= 0;  //180 / 205 = 0
    16'b10110100_11001110 : OUT <= 0;  //180 / 206 = 0
    16'b10110100_11001111 : OUT <= 0;  //180 / 207 = 0
    16'b10110100_11010000 : OUT <= 0;  //180 / 208 = 0
    16'b10110100_11010001 : OUT <= 0;  //180 / 209 = 0
    16'b10110100_11010010 : OUT <= 0;  //180 / 210 = 0
    16'b10110100_11010011 : OUT <= 0;  //180 / 211 = 0
    16'b10110100_11010100 : OUT <= 0;  //180 / 212 = 0
    16'b10110100_11010101 : OUT <= 0;  //180 / 213 = 0
    16'b10110100_11010110 : OUT <= 0;  //180 / 214 = 0
    16'b10110100_11010111 : OUT <= 0;  //180 / 215 = 0
    16'b10110100_11011000 : OUT <= 0;  //180 / 216 = 0
    16'b10110100_11011001 : OUT <= 0;  //180 / 217 = 0
    16'b10110100_11011010 : OUT <= 0;  //180 / 218 = 0
    16'b10110100_11011011 : OUT <= 0;  //180 / 219 = 0
    16'b10110100_11011100 : OUT <= 0;  //180 / 220 = 0
    16'b10110100_11011101 : OUT <= 0;  //180 / 221 = 0
    16'b10110100_11011110 : OUT <= 0;  //180 / 222 = 0
    16'b10110100_11011111 : OUT <= 0;  //180 / 223 = 0
    16'b10110100_11100000 : OUT <= 0;  //180 / 224 = 0
    16'b10110100_11100001 : OUT <= 0;  //180 / 225 = 0
    16'b10110100_11100010 : OUT <= 0;  //180 / 226 = 0
    16'b10110100_11100011 : OUT <= 0;  //180 / 227 = 0
    16'b10110100_11100100 : OUT <= 0;  //180 / 228 = 0
    16'b10110100_11100101 : OUT <= 0;  //180 / 229 = 0
    16'b10110100_11100110 : OUT <= 0;  //180 / 230 = 0
    16'b10110100_11100111 : OUT <= 0;  //180 / 231 = 0
    16'b10110100_11101000 : OUT <= 0;  //180 / 232 = 0
    16'b10110100_11101001 : OUT <= 0;  //180 / 233 = 0
    16'b10110100_11101010 : OUT <= 0;  //180 / 234 = 0
    16'b10110100_11101011 : OUT <= 0;  //180 / 235 = 0
    16'b10110100_11101100 : OUT <= 0;  //180 / 236 = 0
    16'b10110100_11101101 : OUT <= 0;  //180 / 237 = 0
    16'b10110100_11101110 : OUT <= 0;  //180 / 238 = 0
    16'b10110100_11101111 : OUT <= 0;  //180 / 239 = 0
    16'b10110100_11110000 : OUT <= 0;  //180 / 240 = 0
    16'b10110100_11110001 : OUT <= 0;  //180 / 241 = 0
    16'b10110100_11110010 : OUT <= 0;  //180 / 242 = 0
    16'b10110100_11110011 : OUT <= 0;  //180 / 243 = 0
    16'b10110100_11110100 : OUT <= 0;  //180 / 244 = 0
    16'b10110100_11110101 : OUT <= 0;  //180 / 245 = 0
    16'b10110100_11110110 : OUT <= 0;  //180 / 246 = 0
    16'b10110100_11110111 : OUT <= 0;  //180 / 247 = 0
    16'b10110100_11111000 : OUT <= 0;  //180 / 248 = 0
    16'b10110100_11111001 : OUT <= 0;  //180 / 249 = 0
    16'b10110100_11111010 : OUT <= 0;  //180 / 250 = 0
    16'b10110100_11111011 : OUT <= 0;  //180 / 251 = 0
    16'b10110100_11111100 : OUT <= 0;  //180 / 252 = 0
    16'b10110100_11111101 : OUT <= 0;  //180 / 253 = 0
    16'b10110100_11111110 : OUT <= 0;  //180 / 254 = 0
    16'b10110100_11111111 : OUT <= 0;  //180 / 255 = 0
    16'b10110101_00000000 : OUT <= 0;  //181 / 0 = 0
    16'b10110101_00000001 : OUT <= 181;  //181 / 1 = 181
    16'b10110101_00000010 : OUT <= 90;  //181 / 2 = 90
    16'b10110101_00000011 : OUT <= 60;  //181 / 3 = 60
    16'b10110101_00000100 : OUT <= 45;  //181 / 4 = 45
    16'b10110101_00000101 : OUT <= 36;  //181 / 5 = 36
    16'b10110101_00000110 : OUT <= 30;  //181 / 6 = 30
    16'b10110101_00000111 : OUT <= 25;  //181 / 7 = 25
    16'b10110101_00001000 : OUT <= 22;  //181 / 8 = 22
    16'b10110101_00001001 : OUT <= 20;  //181 / 9 = 20
    16'b10110101_00001010 : OUT <= 18;  //181 / 10 = 18
    16'b10110101_00001011 : OUT <= 16;  //181 / 11 = 16
    16'b10110101_00001100 : OUT <= 15;  //181 / 12 = 15
    16'b10110101_00001101 : OUT <= 13;  //181 / 13 = 13
    16'b10110101_00001110 : OUT <= 12;  //181 / 14 = 12
    16'b10110101_00001111 : OUT <= 12;  //181 / 15 = 12
    16'b10110101_00010000 : OUT <= 11;  //181 / 16 = 11
    16'b10110101_00010001 : OUT <= 10;  //181 / 17 = 10
    16'b10110101_00010010 : OUT <= 10;  //181 / 18 = 10
    16'b10110101_00010011 : OUT <= 9;  //181 / 19 = 9
    16'b10110101_00010100 : OUT <= 9;  //181 / 20 = 9
    16'b10110101_00010101 : OUT <= 8;  //181 / 21 = 8
    16'b10110101_00010110 : OUT <= 8;  //181 / 22 = 8
    16'b10110101_00010111 : OUT <= 7;  //181 / 23 = 7
    16'b10110101_00011000 : OUT <= 7;  //181 / 24 = 7
    16'b10110101_00011001 : OUT <= 7;  //181 / 25 = 7
    16'b10110101_00011010 : OUT <= 6;  //181 / 26 = 6
    16'b10110101_00011011 : OUT <= 6;  //181 / 27 = 6
    16'b10110101_00011100 : OUT <= 6;  //181 / 28 = 6
    16'b10110101_00011101 : OUT <= 6;  //181 / 29 = 6
    16'b10110101_00011110 : OUT <= 6;  //181 / 30 = 6
    16'b10110101_00011111 : OUT <= 5;  //181 / 31 = 5
    16'b10110101_00100000 : OUT <= 5;  //181 / 32 = 5
    16'b10110101_00100001 : OUT <= 5;  //181 / 33 = 5
    16'b10110101_00100010 : OUT <= 5;  //181 / 34 = 5
    16'b10110101_00100011 : OUT <= 5;  //181 / 35 = 5
    16'b10110101_00100100 : OUT <= 5;  //181 / 36 = 5
    16'b10110101_00100101 : OUT <= 4;  //181 / 37 = 4
    16'b10110101_00100110 : OUT <= 4;  //181 / 38 = 4
    16'b10110101_00100111 : OUT <= 4;  //181 / 39 = 4
    16'b10110101_00101000 : OUT <= 4;  //181 / 40 = 4
    16'b10110101_00101001 : OUT <= 4;  //181 / 41 = 4
    16'b10110101_00101010 : OUT <= 4;  //181 / 42 = 4
    16'b10110101_00101011 : OUT <= 4;  //181 / 43 = 4
    16'b10110101_00101100 : OUT <= 4;  //181 / 44 = 4
    16'b10110101_00101101 : OUT <= 4;  //181 / 45 = 4
    16'b10110101_00101110 : OUT <= 3;  //181 / 46 = 3
    16'b10110101_00101111 : OUT <= 3;  //181 / 47 = 3
    16'b10110101_00110000 : OUT <= 3;  //181 / 48 = 3
    16'b10110101_00110001 : OUT <= 3;  //181 / 49 = 3
    16'b10110101_00110010 : OUT <= 3;  //181 / 50 = 3
    16'b10110101_00110011 : OUT <= 3;  //181 / 51 = 3
    16'b10110101_00110100 : OUT <= 3;  //181 / 52 = 3
    16'b10110101_00110101 : OUT <= 3;  //181 / 53 = 3
    16'b10110101_00110110 : OUT <= 3;  //181 / 54 = 3
    16'b10110101_00110111 : OUT <= 3;  //181 / 55 = 3
    16'b10110101_00111000 : OUT <= 3;  //181 / 56 = 3
    16'b10110101_00111001 : OUT <= 3;  //181 / 57 = 3
    16'b10110101_00111010 : OUT <= 3;  //181 / 58 = 3
    16'b10110101_00111011 : OUT <= 3;  //181 / 59 = 3
    16'b10110101_00111100 : OUT <= 3;  //181 / 60 = 3
    16'b10110101_00111101 : OUT <= 2;  //181 / 61 = 2
    16'b10110101_00111110 : OUT <= 2;  //181 / 62 = 2
    16'b10110101_00111111 : OUT <= 2;  //181 / 63 = 2
    16'b10110101_01000000 : OUT <= 2;  //181 / 64 = 2
    16'b10110101_01000001 : OUT <= 2;  //181 / 65 = 2
    16'b10110101_01000010 : OUT <= 2;  //181 / 66 = 2
    16'b10110101_01000011 : OUT <= 2;  //181 / 67 = 2
    16'b10110101_01000100 : OUT <= 2;  //181 / 68 = 2
    16'b10110101_01000101 : OUT <= 2;  //181 / 69 = 2
    16'b10110101_01000110 : OUT <= 2;  //181 / 70 = 2
    16'b10110101_01000111 : OUT <= 2;  //181 / 71 = 2
    16'b10110101_01001000 : OUT <= 2;  //181 / 72 = 2
    16'b10110101_01001001 : OUT <= 2;  //181 / 73 = 2
    16'b10110101_01001010 : OUT <= 2;  //181 / 74 = 2
    16'b10110101_01001011 : OUT <= 2;  //181 / 75 = 2
    16'b10110101_01001100 : OUT <= 2;  //181 / 76 = 2
    16'b10110101_01001101 : OUT <= 2;  //181 / 77 = 2
    16'b10110101_01001110 : OUT <= 2;  //181 / 78 = 2
    16'b10110101_01001111 : OUT <= 2;  //181 / 79 = 2
    16'b10110101_01010000 : OUT <= 2;  //181 / 80 = 2
    16'b10110101_01010001 : OUT <= 2;  //181 / 81 = 2
    16'b10110101_01010010 : OUT <= 2;  //181 / 82 = 2
    16'b10110101_01010011 : OUT <= 2;  //181 / 83 = 2
    16'b10110101_01010100 : OUT <= 2;  //181 / 84 = 2
    16'b10110101_01010101 : OUT <= 2;  //181 / 85 = 2
    16'b10110101_01010110 : OUT <= 2;  //181 / 86 = 2
    16'b10110101_01010111 : OUT <= 2;  //181 / 87 = 2
    16'b10110101_01011000 : OUT <= 2;  //181 / 88 = 2
    16'b10110101_01011001 : OUT <= 2;  //181 / 89 = 2
    16'b10110101_01011010 : OUT <= 2;  //181 / 90 = 2
    16'b10110101_01011011 : OUT <= 1;  //181 / 91 = 1
    16'b10110101_01011100 : OUT <= 1;  //181 / 92 = 1
    16'b10110101_01011101 : OUT <= 1;  //181 / 93 = 1
    16'b10110101_01011110 : OUT <= 1;  //181 / 94 = 1
    16'b10110101_01011111 : OUT <= 1;  //181 / 95 = 1
    16'b10110101_01100000 : OUT <= 1;  //181 / 96 = 1
    16'b10110101_01100001 : OUT <= 1;  //181 / 97 = 1
    16'b10110101_01100010 : OUT <= 1;  //181 / 98 = 1
    16'b10110101_01100011 : OUT <= 1;  //181 / 99 = 1
    16'b10110101_01100100 : OUT <= 1;  //181 / 100 = 1
    16'b10110101_01100101 : OUT <= 1;  //181 / 101 = 1
    16'b10110101_01100110 : OUT <= 1;  //181 / 102 = 1
    16'b10110101_01100111 : OUT <= 1;  //181 / 103 = 1
    16'b10110101_01101000 : OUT <= 1;  //181 / 104 = 1
    16'b10110101_01101001 : OUT <= 1;  //181 / 105 = 1
    16'b10110101_01101010 : OUT <= 1;  //181 / 106 = 1
    16'b10110101_01101011 : OUT <= 1;  //181 / 107 = 1
    16'b10110101_01101100 : OUT <= 1;  //181 / 108 = 1
    16'b10110101_01101101 : OUT <= 1;  //181 / 109 = 1
    16'b10110101_01101110 : OUT <= 1;  //181 / 110 = 1
    16'b10110101_01101111 : OUT <= 1;  //181 / 111 = 1
    16'b10110101_01110000 : OUT <= 1;  //181 / 112 = 1
    16'b10110101_01110001 : OUT <= 1;  //181 / 113 = 1
    16'b10110101_01110010 : OUT <= 1;  //181 / 114 = 1
    16'b10110101_01110011 : OUT <= 1;  //181 / 115 = 1
    16'b10110101_01110100 : OUT <= 1;  //181 / 116 = 1
    16'b10110101_01110101 : OUT <= 1;  //181 / 117 = 1
    16'b10110101_01110110 : OUT <= 1;  //181 / 118 = 1
    16'b10110101_01110111 : OUT <= 1;  //181 / 119 = 1
    16'b10110101_01111000 : OUT <= 1;  //181 / 120 = 1
    16'b10110101_01111001 : OUT <= 1;  //181 / 121 = 1
    16'b10110101_01111010 : OUT <= 1;  //181 / 122 = 1
    16'b10110101_01111011 : OUT <= 1;  //181 / 123 = 1
    16'b10110101_01111100 : OUT <= 1;  //181 / 124 = 1
    16'b10110101_01111101 : OUT <= 1;  //181 / 125 = 1
    16'b10110101_01111110 : OUT <= 1;  //181 / 126 = 1
    16'b10110101_01111111 : OUT <= 1;  //181 / 127 = 1
    16'b10110101_10000000 : OUT <= 1;  //181 / 128 = 1
    16'b10110101_10000001 : OUT <= 1;  //181 / 129 = 1
    16'b10110101_10000010 : OUT <= 1;  //181 / 130 = 1
    16'b10110101_10000011 : OUT <= 1;  //181 / 131 = 1
    16'b10110101_10000100 : OUT <= 1;  //181 / 132 = 1
    16'b10110101_10000101 : OUT <= 1;  //181 / 133 = 1
    16'b10110101_10000110 : OUT <= 1;  //181 / 134 = 1
    16'b10110101_10000111 : OUT <= 1;  //181 / 135 = 1
    16'b10110101_10001000 : OUT <= 1;  //181 / 136 = 1
    16'b10110101_10001001 : OUT <= 1;  //181 / 137 = 1
    16'b10110101_10001010 : OUT <= 1;  //181 / 138 = 1
    16'b10110101_10001011 : OUT <= 1;  //181 / 139 = 1
    16'b10110101_10001100 : OUT <= 1;  //181 / 140 = 1
    16'b10110101_10001101 : OUT <= 1;  //181 / 141 = 1
    16'b10110101_10001110 : OUT <= 1;  //181 / 142 = 1
    16'b10110101_10001111 : OUT <= 1;  //181 / 143 = 1
    16'b10110101_10010000 : OUT <= 1;  //181 / 144 = 1
    16'b10110101_10010001 : OUT <= 1;  //181 / 145 = 1
    16'b10110101_10010010 : OUT <= 1;  //181 / 146 = 1
    16'b10110101_10010011 : OUT <= 1;  //181 / 147 = 1
    16'b10110101_10010100 : OUT <= 1;  //181 / 148 = 1
    16'b10110101_10010101 : OUT <= 1;  //181 / 149 = 1
    16'b10110101_10010110 : OUT <= 1;  //181 / 150 = 1
    16'b10110101_10010111 : OUT <= 1;  //181 / 151 = 1
    16'b10110101_10011000 : OUT <= 1;  //181 / 152 = 1
    16'b10110101_10011001 : OUT <= 1;  //181 / 153 = 1
    16'b10110101_10011010 : OUT <= 1;  //181 / 154 = 1
    16'b10110101_10011011 : OUT <= 1;  //181 / 155 = 1
    16'b10110101_10011100 : OUT <= 1;  //181 / 156 = 1
    16'b10110101_10011101 : OUT <= 1;  //181 / 157 = 1
    16'b10110101_10011110 : OUT <= 1;  //181 / 158 = 1
    16'b10110101_10011111 : OUT <= 1;  //181 / 159 = 1
    16'b10110101_10100000 : OUT <= 1;  //181 / 160 = 1
    16'b10110101_10100001 : OUT <= 1;  //181 / 161 = 1
    16'b10110101_10100010 : OUT <= 1;  //181 / 162 = 1
    16'b10110101_10100011 : OUT <= 1;  //181 / 163 = 1
    16'b10110101_10100100 : OUT <= 1;  //181 / 164 = 1
    16'b10110101_10100101 : OUT <= 1;  //181 / 165 = 1
    16'b10110101_10100110 : OUT <= 1;  //181 / 166 = 1
    16'b10110101_10100111 : OUT <= 1;  //181 / 167 = 1
    16'b10110101_10101000 : OUT <= 1;  //181 / 168 = 1
    16'b10110101_10101001 : OUT <= 1;  //181 / 169 = 1
    16'b10110101_10101010 : OUT <= 1;  //181 / 170 = 1
    16'b10110101_10101011 : OUT <= 1;  //181 / 171 = 1
    16'b10110101_10101100 : OUT <= 1;  //181 / 172 = 1
    16'b10110101_10101101 : OUT <= 1;  //181 / 173 = 1
    16'b10110101_10101110 : OUT <= 1;  //181 / 174 = 1
    16'b10110101_10101111 : OUT <= 1;  //181 / 175 = 1
    16'b10110101_10110000 : OUT <= 1;  //181 / 176 = 1
    16'b10110101_10110001 : OUT <= 1;  //181 / 177 = 1
    16'b10110101_10110010 : OUT <= 1;  //181 / 178 = 1
    16'b10110101_10110011 : OUT <= 1;  //181 / 179 = 1
    16'b10110101_10110100 : OUT <= 1;  //181 / 180 = 1
    16'b10110101_10110101 : OUT <= 1;  //181 / 181 = 1
    16'b10110101_10110110 : OUT <= 0;  //181 / 182 = 0
    16'b10110101_10110111 : OUT <= 0;  //181 / 183 = 0
    16'b10110101_10111000 : OUT <= 0;  //181 / 184 = 0
    16'b10110101_10111001 : OUT <= 0;  //181 / 185 = 0
    16'b10110101_10111010 : OUT <= 0;  //181 / 186 = 0
    16'b10110101_10111011 : OUT <= 0;  //181 / 187 = 0
    16'b10110101_10111100 : OUT <= 0;  //181 / 188 = 0
    16'b10110101_10111101 : OUT <= 0;  //181 / 189 = 0
    16'b10110101_10111110 : OUT <= 0;  //181 / 190 = 0
    16'b10110101_10111111 : OUT <= 0;  //181 / 191 = 0
    16'b10110101_11000000 : OUT <= 0;  //181 / 192 = 0
    16'b10110101_11000001 : OUT <= 0;  //181 / 193 = 0
    16'b10110101_11000010 : OUT <= 0;  //181 / 194 = 0
    16'b10110101_11000011 : OUT <= 0;  //181 / 195 = 0
    16'b10110101_11000100 : OUT <= 0;  //181 / 196 = 0
    16'b10110101_11000101 : OUT <= 0;  //181 / 197 = 0
    16'b10110101_11000110 : OUT <= 0;  //181 / 198 = 0
    16'b10110101_11000111 : OUT <= 0;  //181 / 199 = 0
    16'b10110101_11001000 : OUT <= 0;  //181 / 200 = 0
    16'b10110101_11001001 : OUT <= 0;  //181 / 201 = 0
    16'b10110101_11001010 : OUT <= 0;  //181 / 202 = 0
    16'b10110101_11001011 : OUT <= 0;  //181 / 203 = 0
    16'b10110101_11001100 : OUT <= 0;  //181 / 204 = 0
    16'b10110101_11001101 : OUT <= 0;  //181 / 205 = 0
    16'b10110101_11001110 : OUT <= 0;  //181 / 206 = 0
    16'b10110101_11001111 : OUT <= 0;  //181 / 207 = 0
    16'b10110101_11010000 : OUT <= 0;  //181 / 208 = 0
    16'b10110101_11010001 : OUT <= 0;  //181 / 209 = 0
    16'b10110101_11010010 : OUT <= 0;  //181 / 210 = 0
    16'b10110101_11010011 : OUT <= 0;  //181 / 211 = 0
    16'b10110101_11010100 : OUT <= 0;  //181 / 212 = 0
    16'b10110101_11010101 : OUT <= 0;  //181 / 213 = 0
    16'b10110101_11010110 : OUT <= 0;  //181 / 214 = 0
    16'b10110101_11010111 : OUT <= 0;  //181 / 215 = 0
    16'b10110101_11011000 : OUT <= 0;  //181 / 216 = 0
    16'b10110101_11011001 : OUT <= 0;  //181 / 217 = 0
    16'b10110101_11011010 : OUT <= 0;  //181 / 218 = 0
    16'b10110101_11011011 : OUT <= 0;  //181 / 219 = 0
    16'b10110101_11011100 : OUT <= 0;  //181 / 220 = 0
    16'b10110101_11011101 : OUT <= 0;  //181 / 221 = 0
    16'b10110101_11011110 : OUT <= 0;  //181 / 222 = 0
    16'b10110101_11011111 : OUT <= 0;  //181 / 223 = 0
    16'b10110101_11100000 : OUT <= 0;  //181 / 224 = 0
    16'b10110101_11100001 : OUT <= 0;  //181 / 225 = 0
    16'b10110101_11100010 : OUT <= 0;  //181 / 226 = 0
    16'b10110101_11100011 : OUT <= 0;  //181 / 227 = 0
    16'b10110101_11100100 : OUT <= 0;  //181 / 228 = 0
    16'b10110101_11100101 : OUT <= 0;  //181 / 229 = 0
    16'b10110101_11100110 : OUT <= 0;  //181 / 230 = 0
    16'b10110101_11100111 : OUT <= 0;  //181 / 231 = 0
    16'b10110101_11101000 : OUT <= 0;  //181 / 232 = 0
    16'b10110101_11101001 : OUT <= 0;  //181 / 233 = 0
    16'b10110101_11101010 : OUT <= 0;  //181 / 234 = 0
    16'b10110101_11101011 : OUT <= 0;  //181 / 235 = 0
    16'b10110101_11101100 : OUT <= 0;  //181 / 236 = 0
    16'b10110101_11101101 : OUT <= 0;  //181 / 237 = 0
    16'b10110101_11101110 : OUT <= 0;  //181 / 238 = 0
    16'b10110101_11101111 : OUT <= 0;  //181 / 239 = 0
    16'b10110101_11110000 : OUT <= 0;  //181 / 240 = 0
    16'b10110101_11110001 : OUT <= 0;  //181 / 241 = 0
    16'b10110101_11110010 : OUT <= 0;  //181 / 242 = 0
    16'b10110101_11110011 : OUT <= 0;  //181 / 243 = 0
    16'b10110101_11110100 : OUT <= 0;  //181 / 244 = 0
    16'b10110101_11110101 : OUT <= 0;  //181 / 245 = 0
    16'b10110101_11110110 : OUT <= 0;  //181 / 246 = 0
    16'b10110101_11110111 : OUT <= 0;  //181 / 247 = 0
    16'b10110101_11111000 : OUT <= 0;  //181 / 248 = 0
    16'b10110101_11111001 : OUT <= 0;  //181 / 249 = 0
    16'b10110101_11111010 : OUT <= 0;  //181 / 250 = 0
    16'b10110101_11111011 : OUT <= 0;  //181 / 251 = 0
    16'b10110101_11111100 : OUT <= 0;  //181 / 252 = 0
    16'b10110101_11111101 : OUT <= 0;  //181 / 253 = 0
    16'b10110101_11111110 : OUT <= 0;  //181 / 254 = 0
    16'b10110101_11111111 : OUT <= 0;  //181 / 255 = 0
    16'b10110110_00000000 : OUT <= 0;  //182 / 0 = 0
    16'b10110110_00000001 : OUT <= 182;  //182 / 1 = 182
    16'b10110110_00000010 : OUT <= 91;  //182 / 2 = 91
    16'b10110110_00000011 : OUT <= 60;  //182 / 3 = 60
    16'b10110110_00000100 : OUT <= 45;  //182 / 4 = 45
    16'b10110110_00000101 : OUT <= 36;  //182 / 5 = 36
    16'b10110110_00000110 : OUT <= 30;  //182 / 6 = 30
    16'b10110110_00000111 : OUT <= 26;  //182 / 7 = 26
    16'b10110110_00001000 : OUT <= 22;  //182 / 8 = 22
    16'b10110110_00001001 : OUT <= 20;  //182 / 9 = 20
    16'b10110110_00001010 : OUT <= 18;  //182 / 10 = 18
    16'b10110110_00001011 : OUT <= 16;  //182 / 11 = 16
    16'b10110110_00001100 : OUT <= 15;  //182 / 12 = 15
    16'b10110110_00001101 : OUT <= 14;  //182 / 13 = 14
    16'b10110110_00001110 : OUT <= 13;  //182 / 14 = 13
    16'b10110110_00001111 : OUT <= 12;  //182 / 15 = 12
    16'b10110110_00010000 : OUT <= 11;  //182 / 16 = 11
    16'b10110110_00010001 : OUT <= 10;  //182 / 17 = 10
    16'b10110110_00010010 : OUT <= 10;  //182 / 18 = 10
    16'b10110110_00010011 : OUT <= 9;  //182 / 19 = 9
    16'b10110110_00010100 : OUT <= 9;  //182 / 20 = 9
    16'b10110110_00010101 : OUT <= 8;  //182 / 21 = 8
    16'b10110110_00010110 : OUT <= 8;  //182 / 22 = 8
    16'b10110110_00010111 : OUT <= 7;  //182 / 23 = 7
    16'b10110110_00011000 : OUT <= 7;  //182 / 24 = 7
    16'b10110110_00011001 : OUT <= 7;  //182 / 25 = 7
    16'b10110110_00011010 : OUT <= 7;  //182 / 26 = 7
    16'b10110110_00011011 : OUT <= 6;  //182 / 27 = 6
    16'b10110110_00011100 : OUT <= 6;  //182 / 28 = 6
    16'b10110110_00011101 : OUT <= 6;  //182 / 29 = 6
    16'b10110110_00011110 : OUT <= 6;  //182 / 30 = 6
    16'b10110110_00011111 : OUT <= 5;  //182 / 31 = 5
    16'b10110110_00100000 : OUT <= 5;  //182 / 32 = 5
    16'b10110110_00100001 : OUT <= 5;  //182 / 33 = 5
    16'b10110110_00100010 : OUT <= 5;  //182 / 34 = 5
    16'b10110110_00100011 : OUT <= 5;  //182 / 35 = 5
    16'b10110110_00100100 : OUT <= 5;  //182 / 36 = 5
    16'b10110110_00100101 : OUT <= 4;  //182 / 37 = 4
    16'b10110110_00100110 : OUT <= 4;  //182 / 38 = 4
    16'b10110110_00100111 : OUT <= 4;  //182 / 39 = 4
    16'b10110110_00101000 : OUT <= 4;  //182 / 40 = 4
    16'b10110110_00101001 : OUT <= 4;  //182 / 41 = 4
    16'b10110110_00101010 : OUT <= 4;  //182 / 42 = 4
    16'b10110110_00101011 : OUT <= 4;  //182 / 43 = 4
    16'b10110110_00101100 : OUT <= 4;  //182 / 44 = 4
    16'b10110110_00101101 : OUT <= 4;  //182 / 45 = 4
    16'b10110110_00101110 : OUT <= 3;  //182 / 46 = 3
    16'b10110110_00101111 : OUT <= 3;  //182 / 47 = 3
    16'b10110110_00110000 : OUT <= 3;  //182 / 48 = 3
    16'b10110110_00110001 : OUT <= 3;  //182 / 49 = 3
    16'b10110110_00110010 : OUT <= 3;  //182 / 50 = 3
    16'b10110110_00110011 : OUT <= 3;  //182 / 51 = 3
    16'b10110110_00110100 : OUT <= 3;  //182 / 52 = 3
    16'b10110110_00110101 : OUT <= 3;  //182 / 53 = 3
    16'b10110110_00110110 : OUT <= 3;  //182 / 54 = 3
    16'b10110110_00110111 : OUT <= 3;  //182 / 55 = 3
    16'b10110110_00111000 : OUT <= 3;  //182 / 56 = 3
    16'b10110110_00111001 : OUT <= 3;  //182 / 57 = 3
    16'b10110110_00111010 : OUT <= 3;  //182 / 58 = 3
    16'b10110110_00111011 : OUT <= 3;  //182 / 59 = 3
    16'b10110110_00111100 : OUT <= 3;  //182 / 60 = 3
    16'b10110110_00111101 : OUT <= 2;  //182 / 61 = 2
    16'b10110110_00111110 : OUT <= 2;  //182 / 62 = 2
    16'b10110110_00111111 : OUT <= 2;  //182 / 63 = 2
    16'b10110110_01000000 : OUT <= 2;  //182 / 64 = 2
    16'b10110110_01000001 : OUT <= 2;  //182 / 65 = 2
    16'b10110110_01000010 : OUT <= 2;  //182 / 66 = 2
    16'b10110110_01000011 : OUT <= 2;  //182 / 67 = 2
    16'b10110110_01000100 : OUT <= 2;  //182 / 68 = 2
    16'b10110110_01000101 : OUT <= 2;  //182 / 69 = 2
    16'b10110110_01000110 : OUT <= 2;  //182 / 70 = 2
    16'b10110110_01000111 : OUT <= 2;  //182 / 71 = 2
    16'b10110110_01001000 : OUT <= 2;  //182 / 72 = 2
    16'b10110110_01001001 : OUT <= 2;  //182 / 73 = 2
    16'b10110110_01001010 : OUT <= 2;  //182 / 74 = 2
    16'b10110110_01001011 : OUT <= 2;  //182 / 75 = 2
    16'b10110110_01001100 : OUT <= 2;  //182 / 76 = 2
    16'b10110110_01001101 : OUT <= 2;  //182 / 77 = 2
    16'b10110110_01001110 : OUT <= 2;  //182 / 78 = 2
    16'b10110110_01001111 : OUT <= 2;  //182 / 79 = 2
    16'b10110110_01010000 : OUT <= 2;  //182 / 80 = 2
    16'b10110110_01010001 : OUT <= 2;  //182 / 81 = 2
    16'b10110110_01010010 : OUT <= 2;  //182 / 82 = 2
    16'b10110110_01010011 : OUT <= 2;  //182 / 83 = 2
    16'b10110110_01010100 : OUT <= 2;  //182 / 84 = 2
    16'b10110110_01010101 : OUT <= 2;  //182 / 85 = 2
    16'b10110110_01010110 : OUT <= 2;  //182 / 86 = 2
    16'b10110110_01010111 : OUT <= 2;  //182 / 87 = 2
    16'b10110110_01011000 : OUT <= 2;  //182 / 88 = 2
    16'b10110110_01011001 : OUT <= 2;  //182 / 89 = 2
    16'b10110110_01011010 : OUT <= 2;  //182 / 90 = 2
    16'b10110110_01011011 : OUT <= 2;  //182 / 91 = 2
    16'b10110110_01011100 : OUT <= 1;  //182 / 92 = 1
    16'b10110110_01011101 : OUT <= 1;  //182 / 93 = 1
    16'b10110110_01011110 : OUT <= 1;  //182 / 94 = 1
    16'b10110110_01011111 : OUT <= 1;  //182 / 95 = 1
    16'b10110110_01100000 : OUT <= 1;  //182 / 96 = 1
    16'b10110110_01100001 : OUT <= 1;  //182 / 97 = 1
    16'b10110110_01100010 : OUT <= 1;  //182 / 98 = 1
    16'b10110110_01100011 : OUT <= 1;  //182 / 99 = 1
    16'b10110110_01100100 : OUT <= 1;  //182 / 100 = 1
    16'b10110110_01100101 : OUT <= 1;  //182 / 101 = 1
    16'b10110110_01100110 : OUT <= 1;  //182 / 102 = 1
    16'b10110110_01100111 : OUT <= 1;  //182 / 103 = 1
    16'b10110110_01101000 : OUT <= 1;  //182 / 104 = 1
    16'b10110110_01101001 : OUT <= 1;  //182 / 105 = 1
    16'b10110110_01101010 : OUT <= 1;  //182 / 106 = 1
    16'b10110110_01101011 : OUT <= 1;  //182 / 107 = 1
    16'b10110110_01101100 : OUT <= 1;  //182 / 108 = 1
    16'b10110110_01101101 : OUT <= 1;  //182 / 109 = 1
    16'b10110110_01101110 : OUT <= 1;  //182 / 110 = 1
    16'b10110110_01101111 : OUT <= 1;  //182 / 111 = 1
    16'b10110110_01110000 : OUT <= 1;  //182 / 112 = 1
    16'b10110110_01110001 : OUT <= 1;  //182 / 113 = 1
    16'b10110110_01110010 : OUT <= 1;  //182 / 114 = 1
    16'b10110110_01110011 : OUT <= 1;  //182 / 115 = 1
    16'b10110110_01110100 : OUT <= 1;  //182 / 116 = 1
    16'b10110110_01110101 : OUT <= 1;  //182 / 117 = 1
    16'b10110110_01110110 : OUT <= 1;  //182 / 118 = 1
    16'b10110110_01110111 : OUT <= 1;  //182 / 119 = 1
    16'b10110110_01111000 : OUT <= 1;  //182 / 120 = 1
    16'b10110110_01111001 : OUT <= 1;  //182 / 121 = 1
    16'b10110110_01111010 : OUT <= 1;  //182 / 122 = 1
    16'b10110110_01111011 : OUT <= 1;  //182 / 123 = 1
    16'b10110110_01111100 : OUT <= 1;  //182 / 124 = 1
    16'b10110110_01111101 : OUT <= 1;  //182 / 125 = 1
    16'b10110110_01111110 : OUT <= 1;  //182 / 126 = 1
    16'b10110110_01111111 : OUT <= 1;  //182 / 127 = 1
    16'b10110110_10000000 : OUT <= 1;  //182 / 128 = 1
    16'b10110110_10000001 : OUT <= 1;  //182 / 129 = 1
    16'b10110110_10000010 : OUT <= 1;  //182 / 130 = 1
    16'b10110110_10000011 : OUT <= 1;  //182 / 131 = 1
    16'b10110110_10000100 : OUT <= 1;  //182 / 132 = 1
    16'b10110110_10000101 : OUT <= 1;  //182 / 133 = 1
    16'b10110110_10000110 : OUT <= 1;  //182 / 134 = 1
    16'b10110110_10000111 : OUT <= 1;  //182 / 135 = 1
    16'b10110110_10001000 : OUT <= 1;  //182 / 136 = 1
    16'b10110110_10001001 : OUT <= 1;  //182 / 137 = 1
    16'b10110110_10001010 : OUT <= 1;  //182 / 138 = 1
    16'b10110110_10001011 : OUT <= 1;  //182 / 139 = 1
    16'b10110110_10001100 : OUT <= 1;  //182 / 140 = 1
    16'b10110110_10001101 : OUT <= 1;  //182 / 141 = 1
    16'b10110110_10001110 : OUT <= 1;  //182 / 142 = 1
    16'b10110110_10001111 : OUT <= 1;  //182 / 143 = 1
    16'b10110110_10010000 : OUT <= 1;  //182 / 144 = 1
    16'b10110110_10010001 : OUT <= 1;  //182 / 145 = 1
    16'b10110110_10010010 : OUT <= 1;  //182 / 146 = 1
    16'b10110110_10010011 : OUT <= 1;  //182 / 147 = 1
    16'b10110110_10010100 : OUT <= 1;  //182 / 148 = 1
    16'b10110110_10010101 : OUT <= 1;  //182 / 149 = 1
    16'b10110110_10010110 : OUT <= 1;  //182 / 150 = 1
    16'b10110110_10010111 : OUT <= 1;  //182 / 151 = 1
    16'b10110110_10011000 : OUT <= 1;  //182 / 152 = 1
    16'b10110110_10011001 : OUT <= 1;  //182 / 153 = 1
    16'b10110110_10011010 : OUT <= 1;  //182 / 154 = 1
    16'b10110110_10011011 : OUT <= 1;  //182 / 155 = 1
    16'b10110110_10011100 : OUT <= 1;  //182 / 156 = 1
    16'b10110110_10011101 : OUT <= 1;  //182 / 157 = 1
    16'b10110110_10011110 : OUT <= 1;  //182 / 158 = 1
    16'b10110110_10011111 : OUT <= 1;  //182 / 159 = 1
    16'b10110110_10100000 : OUT <= 1;  //182 / 160 = 1
    16'b10110110_10100001 : OUT <= 1;  //182 / 161 = 1
    16'b10110110_10100010 : OUT <= 1;  //182 / 162 = 1
    16'b10110110_10100011 : OUT <= 1;  //182 / 163 = 1
    16'b10110110_10100100 : OUT <= 1;  //182 / 164 = 1
    16'b10110110_10100101 : OUT <= 1;  //182 / 165 = 1
    16'b10110110_10100110 : OUT <= 1;  //182 / 166 = 1
    16'b10110110_10100111 : OUT <= 1;  //182 / 167 = 1
    16'b10110110_10101000 : OUT <= 1;  //182 / 168 = 1
    16'b10110110_10101001 : OUT <= 1;  //182 / 169 = 1
    16'b10110110_10101010 : OUT <= 1;  //182 / 170 = 1
    16'b10110110_10101011 : OUT <= 1;  //182 / 171 = 1
    16'b10110110_10101100 : OUT <= 1;  //182 / 172 = 1
    16'b10110110_10101101 : OUT <= 1;  //182 / 173 = 1
    16'b10110110_10101110 : OUT <= 1;  //182 / 174 = 1
    16'b10110110_10101111 : OUT <= 1;  //182 / 175 = 1
    16'b10110110_10110000 : OUT <= 1;  //182 / 176 = 1
    16'b10110110_10110001 : OUT <= 1;  //182 / 177 = 1
    16'b10110110_10110010 : OUT <= 1;  //182 / 178 = 1
    16'b10110110_10110011 : OUT <= 1;  //182 / 179 = 1
    16'b10110110_10110100 : OUT <= 1;  //182 / 180 = 1
    16'b10110110_10110101 : OUT <= 1;  //182 / 181 = 1
    16'b10110110_10110110 : OUT <= 1;  //182 / 182 = 1
    16'b10110110_10110111 : OUT <= 0;  //182 / 183 = 0
    16'b10110110_10111000 : OUT <= 0;  //182 / 184 = 0
    16'b10110110_10111001 : OUT <= 0;  //182 / 185 = 0
    16'b10110110_10111010 : OUT <= 0;  //182 / 186 = 0
    16'b10110110_10111011 : OUT <= 0;  //182 / 187 = 0
    16'b10110110_10111100 : OUT <= 0;  //182 / 188 = 0
    16'b10110110_10111101 : OUT <= 0;  //182 / 189 = 0
    16'b10110110_10111110 : OUT <= 0;  //182 / 190 = 0
    16'b10110110_10111111 : OUT <= 0;  //182 / 191 = 0
    16'b10110110_11000000 : OUT <= 0;  //182 / 192 = 0
    16'b10110110_11000001 : OUT <= 0;  //182 / 193 = 0
    16'b10110110_11000010 : OUT <= 0;  //182 / 194 = 0
    16'b10110110_11000011 : OUT <= 0;  //182 / 195 = 0
    16'b10110110_11000100 : OUT <= 0;  //182 / 196 = 0
    16'b10110110_11000101 : OUT <= 0;  //182 / 197 = 0
    16'b10110110_11000110 : OUT <= 0;  //182 / 198 = 0
    16'b10110110_11000111 : OUT <= 0;  //182 / 199 = 0
    16'b10110110_11001000 : OUT <= 0;  //182 / 200 = 0
    16'b10110110_11001001 : OUT <= 0;  //182 / 201 = 0
    16'b10110110_11001010 : OUT <= 0;  //182 / 202 = 0
    16'b10110110_11001011 : OUT <= 0;  //182 / 203 = 0
    16'b10110110_11001100 : OUT <= 0;  //182 / 204 = 0
    16'b10110110_11001101 : OUT <= 0;  //182 / 205 = 0
    16'b10110110_11001110 : OUT <= 0;  //182 / 206 = 0
    16'b10110110_11001111 : OUT <= 0;  //182 / 207 = 0
    16'b10110110_11010000 : OUT <= 0;  //182 / 208 = 0
    16'b10110110_11010001 : OUT <= 0;  //182 / 209 = 0
    16'b10110110_11010010 : OUT <= 0;  //182 / 210 = 0
    16'b10110110_11010011 : OUT <= 0;  //182 / 211 = 0
    16'b10110110_11010100 : OUT <= 0;  //182 / 212 = 0
    16'b10110110_11010101 : OUT <= 0;  //182 / 213 = 0
    16'b10110110_11010110 : OUT <= 0;  //182 / 214 = 0
    16'b10110110_11010111 : OUT <= 0;  //182 / 215 = 0
    16'b10110110_11011000 : OUT <= 0;  //182 / 216 = 0
    16'b10110110_11011001 : OUT <= 0;  //182 / 217 = 0
    16'b10110110_11011010 : OUT <= 0;  //182 / 218 = 0
    16'b10110110_11011011 : OUT <= 0;  //182 / 219 = 0
    16'b10110110_11011100 : OUT <= 0;  //182 / 220 = 0
    16'b10110110_11011101 : OUT <= 0;  //182 / 221 = 0
    16'b10110110_11011110 : OUT <= 0;  //182 / 222 = 0
    16'b10110110_11011111 : OUT <= 0;  //182 / 223 = 0
    16'b10110110_11100000 : OUT <= 0;  //182 / 224 = 0
    16'b10110110_11100001 : OUT <= 0;  //182 / 225 = 0
    16'b10110110_11100010 : OUT <= 0;  //182 / 226 = 0
    16'b10110110_11100011 : OUT <= 0;  //182 / 227 = 0
    16'b10110110_11100100 : OUT <= 0;  //182 / 228 = 0
    16'b10110110_11100101 : OUT <= 0;  //182 / 229 = 0
    16'b10110110_11100110 : OUT <= 0;  //182 / 230 = 0
    16'b10110110_11100111 : OUT <= 0;  //182 / 231 = 0
    16'b10110110_11101000 : OUT <= 0;  //182 / 232 = 0
    16'b10110110_11101001 : OUT <= 0;  //182 / 233 = 0
    16'b10110110_11101010 : OUT <= 0;  //182 / 234 = 0
    16'b10110110_11101011 : OUT <= 0;  //182 / 235 = 0
    16'b10110110_11101100 : OUT <= 0;  //182 / 236 = 0
    16'b10110110_11101101 : OUT <= 0;  //182 / 237 = 0
    16'b10110110_11101110 : OUT <= 0;  //182 / 238 = 0
    16'b10110110_11101111 : OUT <= 0;  //182 / 239 = 0
    16'b10110110_11110000 : OUT <= 0;  //182 / 240 = 0
    16'b10110110_11110001 : OUT <= 0;  //182 / 241 = 0
    16'b10110110_11110010 : OUT <= 0;  //182 / 242 = 0
    16'b10110110_11110011 : OUT <= 0;  //182 / 243 = 0
    16'b10110110_11110100 : OUT <= 0;  //182 / 244 = 0
    16'b10110110_11110101 : OUT <= 0;  //182 / 245 = 0
    16'b10110110_11110110 : OUT <= 0;  //182 / 246 = 0
    16'b10110110_11110111 : OUT <= 0;  //182 / 247 = 0
    16'b10110110_11111000 : OUT <= 0;  //182 / 248 = 0
    16'b10110110_11111001 : OUT <= 0;  //182 / 249 = 0
    16'b10110110_11111010 : OUT <= 0;  //182 / 250 = 0
    16'b10110110_11111011 : OUT <= 0;  //182 / 251 = 0
    16'b10110110_11111100 : OUT <= 0;  //182 / 252 = 0
    16'b10110110_11111101 : OUT <= 0;  //182 / 253 = 0
    16'b10110110_11111110 : OUT <= 0;  //182 / 254 = 0
    16'b10110110_11111111 : OUT <= 0;  //182 / 255 = 0
    16'b10110111_00000000 : OUT <= 0;  //183 / 0 = 0
    16'b10110111_00000001 : OUT <= 183;  //183 / 1 = 183
    16'b10110111_00000010 : OUT <= 91;  //183 / 2 = 91
    16'b10110111_00000011 : OUT <= 61;  //183 / 3 = 61
    16'b10110111_00000100 : OUT <= 45;  //183 / 4 = 45
    16'b10110111_00000101 : OUT <= 36;  //183 / 5 = 36
    16'b10110111_00000110 : OUT <= 30;  //183 / 6 = 30
    16'b10110111_00000111 : OUT <= 26;  //183 / 7 = 26
    16'b10110111_00001000 : OUT <= 22;  //183 / 8 = 22
    16'b10110111_00001001 : OUT <= 20;  //183 / 9 = 20
    16'b10110111_00001010 : OUT <= 18;  //183 / 10 = 18
    16'b10110111_00001011 : OUT <= 16;  //183 / 11 = 16
    16'b10110111_00001100 : OUT <= 15;  //183 / 12 = 15
    16'b10110111_00001101 : OUT <= 14;  //183 / 13 = 14
    16'b10110111_00001110 : OUT <= 13;  //183 / 14 = 13
    16'b10110111_00001111 : OUT <= 12;  //183 / 15 = 12
    16'b10110111_00010000 : OUT <= 11;  //183 / 16 = 11
    16'b10110111_00010001 : OUT <= 10;  //183 / 17 = 10
    16'b10110111_00010010 : OUT <= 10;  //183 / 18 = 10
    16'b10110111_00010011 : OUT <= 9;  //183 / 19 = 9
    16'b10110111_00010100 : OUT <= 9;  //183 / 20 = 9
    16'b10110111_00010101 : OUT <= 8;  //183 / 21 = 8
    16'b10110111_00010110 : OUT <= 8;  //183 / 22 = 8
    16'b10110111_00010111 : OUT <= 7;  //183 / 23 = 7
    16'b10110111_00011000 : OUT <= 7;  //183 / 24 = 7
    16'b10110111_00011001 : OUT <= 7;  //183 / 25 = 7
    16'b10110111_00011010 : OUT <= 7;  //183 / 26 = 7
    16'b10110111_00011011 : OUT <= 6;  //183 / 27 = 6
    16'b10110111_00011100 : OUT <= 6;  //183 / 28 = 6
    16'b10110111_00011101 : OUT <= 6;  //183 / 29 = 6
    16'b10110111_00011110 : OUT <= 6;  //183 / 30 = 6
    16'b10110111_00011111 : OUT <= 5;  //183 / 31 = 5
    16'b10110111_00100000 : OUT <= 5;  //183 / 32 = 5
    16'b10110111_00100001 : OUT <= 5;  //183 / 33 = 5
    16'b10110111_00100010 : OUT <= 5;  //183 / 34 = 5
    16'b10110111_00100011 : OUT <= 5;  //183 / 35 = 5
    16'b10110111_00100100 : OUT <= 5;  //183 / 36 = 5
    16'b10110111_00100101 : OUT <= 4;  //183 / 37 = 4
    16'b10110111_00100110 : OUT <= 4;  //183 / 38 = 4
    16'b10110111_00100111 : OUT <= 4;  //183 / 39 = 4
    16'b10110111_00101000 : OUT <= 4;  //183 / 40 = 4
    16'b10110111_00101001 : OUT <= 4;  //183 / 41 = 4
    16'b10110111_00101010 : OUT <= 4;  //183 / 42 = 4
    16'b10110111_00101011 : OUT <= 4;  //183 / 43 = 4
    16'b10110111_00101100 : OUT <= 4;  //183 / 44 = 4
    16'b10110111_00101101 : OUT <= 4;  //183 / 45 = 4
    16'b10110111_00101110 : OUT <= 3;  //183 / 46 = 3
    16'b10110111_00101111 : OUT <= 3;  //183 / 47 = 3
    16'b10110111_00110000 : OUT <= 3;  //183 / 48 = 3
    16'b10110111_00110001 : OUT <= 3;  //183 / 49 = 3
    16'b10110111_00110010 : OUT <= 3;  //183 / 50 = 3
    16'b10110111_00110011 : OUT <= 3;  //183 / 51 = 3
    16'b10110111_00110100 : OUT <= 3;  //183 / 52 = 3
    16'b10110111_00110101 : OUT <= 3;  //183 / 53 = 3
    16'b10110111_00110110 : OUT <= 3;  //183 / 54 = 3
    16'b10110111_00110111 : OUT <= 3;  //183 / 55 = 3
    16'b10110111_00111000 : OUT <= 3;  //183 / 56 = 3
    16'b10110111_00111001 : OUT <= 3;  //183 / 57 = 3
    16'b10110111_00111010 : OUT <= 3;  //183 / 58 = 3
    16'b10110111_00111011 : OUT <= 3;  //183 / 59 = 3
    16'b10110111_00111100 : OUT <= 3;  //183 / 60 = 3
    16'b10110111_00111101 : OUT <= 3;  //183 / 61 = 3
    16'b10110111_00111110 : OUT <= 2;  //183 / 62 = 2
    16'b10110111_00111111 : OUT <= 2;  //183 / 63 = 2
    16'b10110111_01000000 : OUT <= 2;  //183 / 64 = 2
    16'b10110111_01000001 : OUT <= 2;  //183 / 65 = 2
    16'b10110111_01000010 : OUT <= 2;  //183 / 66 = 2
    16'b10110111_01000011 : OUT <= 2;  //183 / 67 = 2
    16'b10110111_01000100 : OUT <= 2;  //183 / 68 = 2
    16'b10110111_01000101 : OUT <= 2;  //183 / 69 = 2
    16'b10110111_01000110 : OUT <= 2;  //183 / 70 = 2
    16'b10110111_01000111 : OUT <= 2;  //183 / 71 = 2
    16'b10110111_01001000 : OUT <= 2;  //183 / 72 = 2
    16'b10110111_01001001 : OUT <= 2;  //183 / 73 = 2
    16'b10110111_01001010 : OUT <= 2;  //183 / 74 = 2
    16'b10110111_01001011 : OUT <= 2;  //183 / 75 = 2
    16'b10110111_01001100 : OUT <= 2;  //183 / 76 = 2
    16'b10110111_01001101 : OUT <= 2;  //183 / 77 = 2
    16'b10110111_01001110 : OUT <= 2;  //183 / 78 = 2
    16'b10110111_01001111 : OUT <= 2;  //183 / 79 = 2
    16'b10110111_01010000 : OUT <= 2;  //183 / 80 = 2
    16'b10110111_01010001 : OUT <= 2;  //183 / 81 = 2
    16'b10110111_01010010 : OUT <= 2;  //183 / 82 = 2
    16'b10110111_01010011 : OUT <= 2;  //183 / 83 = 2
    16'b10110111_01010100 : OUT <= 2;  //183 / 84 = 2
    16'b10110111_01010101 : OUT <= 2;  //183 / 85 = 2
    16'b10110111_01010110 : OUT <= 2;  //183 / 86 = 2
    16'b10110111_01010111 : OUT <= 2;  //183 / 87 = 2
    16'b10110111_01011000 : OUT <= 2;  //183 / 88 = 2
    16'b10110111_01011001 : OUT <= 2;  //183 / 89 = 2
    16'b10110111_01011010 : OUT <= 2;  //183 / 90 = 2
    16'b10110111_01011011 : OUT <= 2;  //183 / 91 = 2
    16'b10110111_01011100 : OUT <= 1;  //183 / 92 = 1
    16'b10110111_01011101 : OUT <= 1;  //183 / 93 = 1
    16'b10110111_01011110 : OUT <= 1;  //183 / 94 = 1
    16'b10110111_01011111 : OUT <= 1;  //183 / 95 = 1
    16'b10110111_01100000 : OUT <= 1;  //183 / 96 = 1
    16'b10110111_01100001 : OUT <= 1;  //183 / 97 = 1
    16'b10110111_01100010 : OUT <= 1;  //183 / 98 = 1
    16'b10110111_01100011 : OUT <= 1;  //183 / 99 = 1
    16'b10110111_01100100 : OUT <= 1;  //183 / 100 = 1
    16'b10110111_01100101 : OUT <= 1;  //183 / 101 = 1
    16'b10110111_01100110 : OUT <= 1;  //183 / 102 = 1
    16'b10110111_01100111 : OUT <= 1;  //183 / 103 = 1
    16'b10110111_01101000 : OUT <= 1;  //183 / 104 = 1
    16'b10110111_01101001 : OUT <= 1;  //183 / 105 = 1
    16'b10110111_01101010 : OUT <= 1;  //183 / 106 = 1
    16'b10110111_01101011 : OUT <= 1;  //183 / 107 = 1
    16'b10110111_01101100 : OUT <= 1;  //183 / 108 = 1
    16'b10110111_01101101 : OUT <= 1;  //183 / 109 = 1
    16'b10110111_01101110 : OUT <= 1;  //183 / 110 = 1
    16'b10110111_01101111 : OUT <= 1;  //183 / 111 = 1
    16'b10110111_01110000 : OUT <= 1;  //183 / 112 = 1
    16'b10110111_01110001 : OUT <= 1;  //183 / 113 = 1
    16'b10110111_01110010 : OUT <= 1;  //183 / 114 = 1
    16'b10110111_01110011 : OUT <= 1;  //183 / 115 = 1
    16'b10110111_01110100 : OUT <= 1;  //183 / 116 = 1
    16'b10110111_01110101 : OUT <= 1;  //183 / 117 = 1
    16'b10110111_01110110 : OUT <= 1;  //183 / 118 = 1
    16'b10110111_01110111 : OUT <= 1;  //183 / 119 = 1
    16'b10110111_01111000 : OUT <= 1;  //183 / 120 = 1
    16'b10110111_01111001 : OUT <= 1;  //183 / 121 = 1
    16'b10110111_01111010 : OUT <= 1;  //183 / 122 = 1
    16'b10110111_01111011 : OUT <= 1;  //183 / 123 = 1
    16'b10110111_01111100 : OUT <= 1;  //183 / 124 = 1
    16'b10110111_01111101 : OUT <= 1;  //183 / 125 = 1
    16'b10110111_01111110 : OUT <= 1;  //183 / 126 = 1
    16'b10110111_01111111 : OUT <= 1;  //183 / 127 = 1
    16'b10110111_10000000 : OUT <= 1;  //183 / 128 = 1
    16'b10110111_10000001 : OUT <= 1;  //183 / 129 = 1
    16'b10110111_10000010 : OUT <= 1;  //183 / 130 = 1
    16'b10110111_10000011 : OUT <= 1;  //183 / 131 = 1
    16'b10110111_10000100 : OUT <= 1;  //183 / 132 = 1
    16'b10110111_10000101 : OUT <= 1;  //183 / 133 = 1
    16'b10110111_10000110 : OUT <= 1;  //183 / 134 = 1
    16'b10110111_10000111 : OUT <= 1;  //183 / 135 = 1
    16'b10110111_10001000 : OUT <= 1;  //183 / 136 = 1
    16'b10110111_10001001 : OUT <= 1;  //183 / 137 = 1
    16'b10110111_10001010 : OUT <= 1;  //183 / 138 = 1
    16'b10110111_10001011 : OUT <= 1;  //183 / 139 = 1
    16'b10110111_10001100 : OUT <= 1;  //183 / 140 = 1
    16'b10110111_10001101 : OUT <= 1;  //183 / 141 = 1
    16'b10110111_10001110 : OUT <= 1;  //183 / 142 = 1
    16'b10110111_10001111 : OUT <= 1;  //183 / 143 = 1
    16'b10110111_10010000 : OUT <= 1;  //183 / 144 = 1
    16'b10110111_10010001 : OUT <= 1;  //183 / 145 = 1
    16'b10110111_10010010 : OUT <= 1;  //183 / 146 = 1
    16'b10110111_10010011 : OUT <= 1;  //183 / 147 = 1
    16'b10110111_10010100 : OUT <= 1;  //183 / 148 = 1
    16'b10110111_10010101 : OUT <= 1;  //183 / 149 = 1
    16'b10110111_10010110 : OUT <= 1;  //183 / 150 = 1
    16'b10110111_10010111 : OUT <= 1;  //183 / 151 = 1
    16'b10110111_10011000 : OUT <= 1;  //183 / 152 = 1
    16'b10110111_10011001 : OUT <= 1;  //183 / 153 = 1
    16'b10110111_10011010 : OUT <= 1;  //183 / 154 = 1
    16'b10110111_10011011 : OUT <= 1;  //183 / 155 = 1
    16'b10110111_10011100 : OUT <= 1;  //183 / 156 = 1
    16'b10110111_10011101 : OUT <= 1;  //183 / 157 = 1
    16'b10110111_10011110 : OUT <= 1;  //183 / 158 = 1
    16'b10110111_10011111 : OUT <= 1;  //183 / 159 = 1
    16'b10110111_10100000 : OUT <= 1;  //183 / 160 = 1
    16'b10110111_10100001 : OUT <= 1;  //183 / 161 = 1
    16'b10110111_10100010 : OUT <= 1;  //183 / 162 = 1
    16'b10110111_10100011 : OUT <= 1;  //183 / 163 = 1
    16'b10110111_10100100 : OUT <= 1;  //183 / 164 = 1
    16'b10110111_10100101 : OUT <= 1;  //183 / 165 = 1
    16'b10110111_10100110 : OUT <= 1;  //183 / 166 = 1
    16'b10110111_10100111 : OUT <= 1;  //183 / 167 = 1
    16'b10110111_10101000 : OUT <= 1;  //183 / 168 = 1
    16'b10110111_10101001 : OUT <= 1;  //183 / 169 = 1
    16'b10110111_10101010 : OUT <= 1;  //183 / 170 = 1
    16'b10110111_10101011 : OUT <= 1;  //183 / 171 = 1
    16'b10110111_10101100 : OUT <= 1;  //183 / 172 = 1
    16'b10110111_10101101 : OUT <= 1;  //183 / 173 = 1
    16'b10110111_10101110 : OUT <= 1;  //183 / 174 = 1
    16'b10110111_10101111 : OUT <= 1;  //183 / 175 = 1
    16'b10110111_10110000 : OUT <= 1;  //183 / 176 = 1
    16'b10110111_10110001 : OUT <= 1;  //183 / 177 = 1
    16'b10110111_10110010 : OUT <= 1;  //183 / 178 = 1
    16'b10110111_10110011 : OUT <= 1;  //183 / 179 = 1
    16'b10110111_10110100 : OUT <= 1;  //183 / 180 = 1
    16'b10110111_10110101 : OUT <= 1;  //183 / 181 = 1
    16'b10110111_10110110 : OUT <= 1;  //183 / 182 = 1
    16'b10110111_10110111 : OUT <= 1;  //183 / 183 = 1
    16'b10110111_10111000 : OUT <= 0;  //183 / 184 = 0
    16'b10110111_10111001 : OUT <= 0;  //183 / 185 = 0
    16'b10110111_10111010 : OUT <= 0;  //183 / 186 = 0
    16'b10110111_10111011 : OUT <= 0;  //183 / 187 = 0
    16'b10110111_10111100 : OUT <= 0;  //183 / 188 = 0
    16'b10110111_10111101 : OUT <= 0;  //183 / 189 = 0
    16'b10110111_10111110 : OUT <= 0;  //183 / 190 = 0
    16'b10110111_10111111 : OUT <= 0;  //183 / 191 = 0
    16'b10110111_11000000 : OUT <= 0;  //183 / 192 = 0
    16'b10110111_11000001 : OUT <= 0;  //183 / 193 = 0
    16'b10110111_11000010 : OUT <= 0;  //183 / 194 = 0
    16'b10110111_11000011 : OUT <= 0;  //183 / 195 = 0
    16'b10110111_11000100 : OUT <= 0;  //183 / 196 = 0
    16'b10110111_11000101 : OUT <= 0;  //183 / 197 = 0
    16'b10110111_11000110 : OUT <= 0;  //183 / 198 = 0
    16'b10110111_11000111 : OUT <= 0;  //183 / 199 = 0
    16'b10110111_11001000 : OUT <= 0;  //183 / 200 = 0
    16'b10110111_11001001 : OUT <= 0;  //183 / 201 = 0
    16'b10110111_11001010 : OUT <= 0;  //183 / 202 = 0
    16'b10110111_11001011 : OUT <= 0;  //183 / 203 = 0
    16'b10110111_11001100 : OUT <= 0;  //183 / 204 = 0
    16'b10110111_11001101 : OUT <= 0;  //183 / 205 = 0
    16'b10110111_11001110 : OUT <= 0;  //183 / 206 = 0
    16'b10110111_11001111 : OUT <= 0;  //183 / 207 = 0
    16'b10110111_11010000 : OUT <= 0;  //183 / 208 = 0
    16'b10110111_11010001 : OUT <= 0;  //183 / 209 = 0
    16'b10110111_11010010 : OUT <= 0;  //183 / 210 = 0
    16'b10110111_11010011 : OUT <= 0;  //183 / 211 = 0
    16'b10110111_11010100 : OUT <= 0;  //183 / 212 = 0
    16'b10110111_11010101 : OUT <= 0;  //183 / 213 = 0
    16'b10110111_11010110 : OUT <= 0;  //183 / 214 = 0
    16'b10110111_11010111 : OUT <= 0;  //183 / 215 = 0
    16'b10110111_11011000 : OUT <= 0;  //183 / 216 = 0
    16'b10110111_11011001 : OUT <= 0;  //183 / 217 = 0
    16'b10110111_11011010 : OUT <= 0;  //183 / 218 = 0
    16'b10110111_11011011 : OUT <= 0;  //183 / 219 = 0
    16'b10110111_11011100 : OUT <= 0;  //183 / 220 = 0
    16'b10110111_11011101 : OUT <= 0;  //183 / 221 = 0
    16'b10110111_11011110 : OUT <= 0;  //183 / 222 = 0
    16'b10110111_11011111 : OUT <= 0;  //183 / 223 = 0
    16'b10110111_11100000 : OUT <= 0;  //183 / 224 = 0
    16'b10110111_11100001 : OUT <= 0;  //183 / 225 = 0
    16'b10110111_11100010 : OUT <= 0;  //183 / 226 = 0
    16'b10110111_11100011 : OUT <= 0;  //183 / 227 = 0
    16'b10110111_11100100 : OUT <= 0;  //183 / 228 = 0
    16'b10110111_11100101 : OUT <= 0;  //183 / 229 = 0
    16'b10110111_11100110 : OUT <= 0;  //183 / 230 = 0
    16'b10110111_11100111 : OUT <= 0;  //183 / 231 = 0
    16'b10110111_11101000 : OUT <= 0;  //183 / 232 = 0
    16'b10110111_11101001 : OUT <= 0;  //183 / 233 = 0
    16'b10110111_11101010 : OUT <= 0;  //183 / 234 = 0
    16'b10110111_11101011 : OUT <= 0;  //183 / 235 = 0
    16'b10110111_11101100 : OUT <= 0;  //183 / 236 = 0
    16'b10110111_11101101 : OUT <= 0;  //183 / 237 = 0
    16'b10110111_11101110 : OUT <= 0;  //183 / 238 = 0
    16'b10110111_11101111 : OUT <= 0;  //183 / 239 = 0
    16'b10110111_11110000 : OUT <= 0;  //183 / 240 = 0
    16'b10110111_11110001 : OUT <= 0;  //183 / 241 = 0
    16'b10110111_11110010 : OUT <= 0;  //183 / 242 = 0
    16'b10110111_11110011 : OUT <= 0;  //183 / 243 = 0
    16'b10110111_11110100 : OUT <= 0;  //183 / 244 = 0
    16'b10110111_11110101 : OUT <= 0;  //183 / 245 = 0
    16'b10110111_11110110 : OUT <= 0;  //183 / 246 = 0
    16'b10110111_11110111 : OUT <= 0;  //183 / 247 = 0
    16'b10110111_11111000 : OUT <= 0;  //183 / 248 = 0
    16'b10110111_11111001 : OUT <= 0;  //183 / 249 = 0
    16'b10110111_11111010 : OUT <= 0;  //183 / 250 = 0
    16'b10110111_11111011 : OUT <= 0;  //183 / 251 = 0
    16'b10110111_11111100 : OUT <= 0;  //183 / 252 = 0
    16'b10110111_11111101 : OUT <= 0;  //183 / 253 = 0
    16'b10110111_11111110 : OUT <= 0;  //183 / 254 = 0
    16'b10110111_11111111 : OUT <= 0;  //183 / 255 = 0
    16'b10111000_00000000 : OUT <= 0;  //184 / 0 = 0
    16'b10111000_00000001 : OUT <= 184;  //184 / 1 = 184
    16'b10111000_00000010 : OUT <= 92;  //184 / 2 = 92
    16'b10111000_00000011 : OUT <= 61;  //184 / 3 = 61
    16'b10111000_00000100 : OUT <= 46;  //184 / 4 = 46
    16'b10111000_00000101 : OUT <= 36;  //184 / 5 = 36
    16'b10111000_00000110 : OUT <= 30;  //184 / 6 = 30
    16'b10111000_00000111 : OUT <= 26;  //184 / 7 = 26
    16'b10111000_00001000 : OUT <= 23;  //184 / 8 = 23
    16'b10111000_00001001 : OUT <= 20;  //184 / 9 = 20
    16'b10111000_00001010 : OUT <= 18;  //184 / 10 = 18
    16'b10111000_00001011 : OUT <= 16;  //184 / 11 = 16
    16'b10111000_00001100 : OUT <= 15;  //184 / 12 = 15
    16'b10111000_00001101 : OUT <= 14;  //184 / 13 = 14
    16'b10111000_00001110 : OUT <= 13;  //184 / 14 = 13
    16'b10111000_00001111 : OUT <= 12;  //184 / 15 = 12
    16'b10111000_00010000 : OUT <= 11;  //184 / 16 = 11
    16'b10111000_00010001 : OUT <= 10;  //184 / 17 = 10
    16'b10111000_00010010 : OUT <= 10;  //184 / 18 = 10
    16'b10111000_00010011 : OUT <= 9;  //184 / 19 = 9
    16'b10111000_00010100 : OUT <= 9;  //184 / 20 = 9
    16'b10111000_00010101 : OUT <= 8;  //184 / 21 = 8
    16'b10111000_00010110 : OUT <= 8;  //184 / 22 = 8
    16'b10111000_00010111 : OUT <= 8;  //184 / 23 = 8
    16'b10111000_00011000 : OUT <= 7;  //184 / 24 = 7
    16'b10111000_00011001 : OUT <= 7;  //184 / 25 = 7
    16'b10111000_00011010 : OUT <= 7;  //184 / 26 = 7
    16'b10111000_00011011 : OUT <= 6;  //184 / 27 = 6
    16'b10111000_00011100 : OUT <= 6;  //184 / 28 = 6
    16'b10111000_00011101 : OUT <= 6;  //184 / 29 = 6
    16'b10111000_00011110 : OUT <= 6;  //184 / 30 = 6
    16'b10111000_00011111 : OUT <= 5;  //184 / 31 = 5
    16'b10111000_00100000 : OUT <= 5;  //184 / 32 = 5
    16'b10111000_00100001 : OUT <= 5;  //184 / 33 = 5
    16'b10111000_00100010 : OUT <= 5;  //184 / 34 = 5
    16'b10111000_00100011 : OUT <= 5;  //184 / 35 = 5
    16'b10111000_00100100 : OUT <= 5;  //184 / 36 = 5
    16'b10111000_00100101 : OUT <= 4;  //184 / 37 = 4
    16'b10111000_00100110 : OUT <= 4;  //184 / 38 = 4
    16'b10111000_00100111 : OUT <= 4;  //184 / 39 = 4
    16'b10111000_00101000 : OUT <= 4;  //184 / 40 = 4
    16'b10111000_00101001 : OUT <= 4;  //184 / 41 = 4
    16'b10111000_00101010 : OUT <= 4;  //184 / 42 = 4
    16'b10111000_00101011 : OUT <= 4;  //184 / 43 = 4
    16'b10111000_00101100 : OUT <= 4;  //184 / 44 = 4
    16'b10111000_00101101 : OUT <= 4;  //184 / 45 = 4
    16'b10111000_00101110 : OUT <= 4;  //184 / 46 = 4
    16'b10111000_00101111 : OUT <= 3;  //184 / 47 = 3
    16'b10111000_00110000 : OUT <= 3;  //184 / 48 = 3
    16'b10111000_00110001 : OUT <= 3;  //184 / 49 = 3
    16'b10111000_00110010 : OUT <= 3;  //184 / 50 = 3
    16'b10111000_00110011 : OUT <= 3;  //184 / 51 = 3
    16'b10111000_00110100 : OUT <= 3;  //184 / 52 = 3
    16'b10111000_00110101 : OUT <= 3;  //184 / 53 = 3
    16'b10111000_00110110 : OUT <= 3;  //184 / 54 = 3
    16'b10111000_00110111 : OUT <= 3;  //184 / 55 = 3
    16'b10111000_00111000 : OUT <= 3;  //184 / 56 = 3
    16'b10111000_00111001 : OUT <= 3;  //184 / 57 = 3
    16'b10111000_00111010 : OUT <= 3;  //184 / 58 = 3
    16'b10111000_00111011 : OUT <= 3;  //184 / 59 = 3
    16'b10111000_00111100 : OUT <= 3;  //184 / 60 = 3
    16'b10111000_00111101 : OUT <= 3;  //184 / 61 = 3
    16'b10111000_00111110 : OUT <= 2;  //184 / 62 = 2
    16'b10111000_00111111 : OUT <= 2;  //184 / 63 = 2
    16'b10111000_01000000 : OUT <= 2;  //184 / 64 = 2
    16'b10111000_01000001 : OUT <= 2;  //184 / 65 = 2
    16'b10111000_01000010 : OUT <= 2;  //184 / 66 = 2
    16'b10111000_01000011 : OUT <= 2;  //184 / 67 = 2
    16'b10111000_01000100 : OUT <= 2;  //184 / 68 = 2
    16'b10111000_01000101 : OUT <= 2;  //184 / 69 = 2
    16'b10111000_01000110 : OUT <= 2;  //184 / 70 = 2
    16'b10111000_01000111 : OUT <= 2;  //184 / 71 = 2
    16'b10111000_01001000 : OUT <= 2;  //184 / 72 = 2
    16'b10111000_01001001 : OUT <= 2;  //184 / 73 = 2
    16'b10111000_01001010 : OUT <= 2;  //184 / 74 = 2
    16'b10111000_01001011 : OUT <= 2;  //184 / 75 = 2
    16'b10111000_01001100 : OUT <= 2;  //184 / 76 = 2
    16'b10111000_01001101 : OUT <= 2;  //184 / 77 = 2
    16'b10111000_01001110 : OUT <= 2;  //184 / 78 = 2
    16'b10111000_01001111 : OUT <= 2;  //184 / 79 = 2
    16'b10111000_01010000 : OUT <= 2;  //184 / 80 = 2
    16'b10111000_01010001 : OUT <= 2;  //184 / 81 = 2
    16'b10111000_01010010 : OUT <= 2;  //184 / 82 = 2
    16'b10111000_01010011 : OUT <= 2;  //184 / 83 = 2
    16'b10111000_01010100 : OUT <= 2;  //184 / 84 = 2
    16'b10111000_01010101 : OUT <= 2;  //184 / 85 = 2
    16'b10111000_01010110 : OUT <= 2;  //184 / 86 = 2
    16'b10111000_01010111 : OUT <= 2;  //184 / 87 = 2
    16'b10111000_01011000 : OUT <= 2;  //184 / 88 = 2
    16'b10111000_01011001 : OUT <= 2;  //184 / 89 = 2
    16'b10111000_01011010 : OUT <= 2;  //184 / 90 = 2
    16'b10111000_01011011 : OUT <= 2;  //184 / 91 = 2
    16'b10111000_01011100 : OUT <= 2;  //184 / 92 = 2
    16'b10111000_01011101 : OUT <= 1;  //184 / 93 = 1
    16'b10111000_01011110 : OUT <= 1;  //184 / 94 = 1
    16'b10111000_01011111 : OUT <= 1;  //184 / 95 = 1
    16'b10111000_01100000 : OUT <= 1;  //184 / 96 = 1
    16'b10111000_01100001 : OUT <= 1;  //184 / 97 = 1
    16'b10111000_01100010 : OUT <= 1;  //184 / 98 = 1
    16'b10111000_01100011 : OUT <= 1;  //184 / 99 = 1
    16'b10111000_01100100 : OUT <= 1;  //184 / 100 = 1
    16'b10111000_01100101 : OUT <= 1;  //184 / 101 = 1
    16'b10111000_01100110 : OUT <= 1;  //184 / 102 = 1
    16'b10111000_01100111 : OUT <= 1;  //184 / 103 = 1
    16'b10111000_01101000 : OUT <= 1;  //184 / 104 = 1
    16'b10111000_01101001 : OUT <= 1;  //184 / 105 = 1
    16'b10111000_01101010 : OUT <= 1;  //184 / 106 = 1
    16'b10111000_01101011 : OUT <= 1;  //184 / 107 = 1
    16'b10111000_01101100 : OUT <= 1;  //184 / 108 = 1
    16'b10111000_01101101 : OUT <= 1;  //184 / 109 = 1
    16'b10111000_01101110 : OUT <= 1;  //184 / 110 = 1
    16'b10111000_01101111 : OUT <= 1;  //184 / 111 = 1
    16'b10111000_01110000 : OUT <= 1;  //184 / 112 = 1
    16'b10111000_01110001 : OUT <= 1;  //184 / 113 = 1
    16'b10111000_01110010 : OUT <= 1;  //184 / 114 = 1
    16'b10111000_01110011 : OUT <= 1;  //184 / 115 = 1
    16'b10111000_01110100 : OUT <= 1;  //184 / 116 = 1
    16'b10111000_01110101 : OUT <= 1;  //184 / 117 = 1
    16'b10111000_01110110 : OUT <= 1;  //184 / 118 = 1
    16'b10111000_01110111 : OUT <= 1;  //184 / 119 = 1
    16'b10111000_01111000 : OUT <= 1;  //184 / 120 = 1
    16'b10111000_01111001 : OUT <= 1;  //184 / 121 = 1
    16'b10111000_01111010 : OUT <= 1;  //184 / 122 = 1
    16'b10111000_01111011 : OUT <= 1;  //184 / 123 = 1
    16'b10111000_01111100 : OUT <= 1;  //184 / 124 = 1
    16'b10111000_01111101 : OUT <= 1;  //184 / 125 = 1
    16'b10111000_01111110 : OUT <= 1;  //184 / 126 = 1
    16'b10111000_01111111 : OUT <= 1;  //184 / 127 = 1
    16'b10111000_10000000 : OUT <= 1;  //184 / 128 = 1
    16'b10111000_10000001 : OUT <= 1;  //184 / 129 = 1
    16'b10111000_10000010 : OUT <= 1;  //184 / 130 = 1
    16'b10111000_10000011 : OUT <= 1;  //184 / 131 = 1
    16'b10111000_10000100 : OUT <= 1;  //184 / 132 = 1
    16'b10111000_10000101 : OUT <= 1;  //184 / 133 = 1
    16'b10111000_10000110 : OUT <= 1;  //184 / 134 = 1
    16'b10111000_10000111 : OUT <= 1;  //184 / 135 = 1
    16'b10111000_10001000 : OUT <= 1;  //184 / 136 = 1
    16'b10111000_10001001 : OUT <= 1;  //184 / 137 = 1
    16'b10111000_10001010 : OUT <= 1;  //184 / 138 = 1
    16'b10111000_10001011 : OUT <= 1;  //184 / 139 = 1
    16'b10111000_10001100 : OUT <= 1;  //184 / 140 = 1
    16'b10111000_10001101 : OUT <= 1;  //184 / 141 = 1
    16'b10111000_10001110 : OUT <= 1;  //184 / 142 = 1
    16'b10111000_10001111 : OUT <= 1;  //184 / 143 = 1
    16'b10111000_10010000 : OUT <= 1;  //184 / 144 = 1
    16'b10111000_10010001 : OUT <= 1;  //184 / 145 = 1
    16'b10111000_10010010 : OUT <= 1;  //184 / 146 = 1
    16'b10111000_10010011 : OUT <= 1;  //184 / 147 = 1
    16'b10111000_10010100 : OUT <= 1;  //184 / 148 = 1
    16'b10111000_10010101 : OUT <= 1;  //184 / 149 = 1
    16'b10111000_10010110 : OUT <= 1;  //184 / 150 = 1
    16'b10111000_10010111 : OUT <= 1;  //184 / 151 = 1
    16'b10111000_10011000 : OUT <= 1;  //184 / 152 = 1
    16'b10111000_10011001 : OUT <= 1;  //184 / 153 = 1
    16'b10111000_10011010 : OUT <= 1;  //184 / 154 = 1
    16'b10111000_10011011 : OUT <= 1;  //184 / 155 = 1
    16'b10111000_10011100 : OUT <= 1;  //184 / 156 = 1
    16'b10111000_10011101 : OUT <= 1;  //184 / 157 = 1
    16'b10111000_10011110 : OUT <= 1;  //184 / 158 = 1
    16'b10111000_10011111 : OUT <= 1;  //184 / 159 = 1
    16'b10111000_10100000 : OUT <= 1;  //184 / 160 = 1
    16'b10111000_10100001 : OUT <= 1;  //184 / 161 = 1
    16'b10111000_10100010 : OUT <= 1;  //184 / 162 = 1
    16'b10111000_10100011 : OUT <= 1;  //184 / 163 = 1
    16'b10111000_10100100 : OUT <= 1;  //184 / 164 = 1
    16'b10111000_10100101 : OUT <= 1;  //184 / 165 = 1
    16'b10111000_10100110 : OUT <= 1;  //184 / 166 = 1
    16'b10111000_10100111 : OUT <= 1;  //184 / 167 = 1
    16'b10111000_10101000 : OUT <= 1;  //184 / 168 = 1
    16'b10111000_10101001 : OUT <= 1;  //184 / 169 = 1
    16'b10111000_10101010 : OUT <= 1;  //184 / 170 = 1
    16'b10111000_10101011 : OUT <= 1;  //184 / 171 = 1
    16'b10111000_10101100 : OUT <= 1;  //184 / 172 = 1
    16'b10111000_10101101 : OUT <= 1;  //184 / 173 = 1
    16'b10111000_10101110 : OUT <= 1;  //184 / 174 = 1
    16'b10111000_10101111 : OUT <= 1;  //184 / 175 = 1
    16'b10111000_10110000 : OUT <= 1;  //184 / 176 = 1
    16'b10111000_10110001 : OUT <= 1;  //184 / 177 = 1
    16'b10111000_10110010 : OUT <= 1;  //184 / 178 = 1
    16'b10111000_10110011 : OUT <= 1;  //184 / 179 = 1
    16'b10111000_10110100 : OUT <= 1;  //184 / 180 = 1
    16'b10111000_10110101 : OUT <= 1;  //184 / 181 = 1
    16'b10111000_10110110 : OUT <= 1;  //184 / 182 = 1
    16'b10111000_10110111 : OUT <= 1;  //184 / 183 = 1
    16'b10111000_10111000 : OUT <= 1;  //184 / 184 = 1
    16'b10111000_10111001 : OUT <= 0;  //184 / 185 = 0
    16'b10111000_10111010 : OUT <= 0;  //184 / 186 = 0
    16'b10111000_10111011 : OUT <= 0;  //184 / 187 = 0
    16'b10111000_10111100 : OUT <= 0;  //184 / 188 = 0
    16'b10111000_10111101 : OUT <= 0;  //184 / 189 = 0
    16'b10111000_10111110 : OUT <= 0;  //184 / 190 = 0
    16'b10111000_10111111 : OUT <= 0;  //184 / 191 = 0
    16'b10111000_11000000 : OUT <= 0;  //184 / 192 = 0
    16'b10111000_11000001 : OUT <= 0;  //184 / 193 = 0
    16'b10111000_11000010 : OUT <= 0;  //184 / 194 = 0
    16'b10111000_11000011 : OUT <= 0;  //184 / 195 = 0
    16'b10111000_11000100 : OUT <= 0;  //184 / 196 = 0
    16'b10111000_11000101 : OUT <= 0;  //184 / 197 = 0
    16'b10111000_11000110 : OUT <= 0;  //184 / 198 = 0
    16'b10111000_11000111 : OUT <= 0;  //184 / 199 = 0
    16'b10111000_11001000 : OUT <= 0;  //184 / 200 = 0
    16'b10111000_11001001 : OUT <= 0;  //184 / 201 = 0
    16'b10111000_11001010 : OUT <= 0;  //184 / 202 = 0
    16'b10111000_11001011 : OUT <= 0;  //184 / 203 = 0
    16'b10111000_11001100 : OUT <= 0;  //184 / 204 = 0
    16'b10111000_11001101 : OUT <= 0;  //184 / 205 = 0
    16'b10111000_11001110 : OUT <= 0;  //184 / 206 = 0
    16'b10111000_11001111 : OUT <= 0;  //184 / 207 = 0
    16'b10111000_11010000 : OUT <= 0;  //184 / 208 = 0
    16'b10111000_11010001 : OUT <= 0;  //184 / 209 = 0
    16'b10111000_11010010 : OUT <= 0;  //184 / 210 = 0
    16'b10111000_11010011 : OUT <= 0;  //184 / 211 = 0
    16'b10111000_11010100 : OUT <= 0;  //184 / 212 = 0
    16'b10111000_11010101 : OUT <= 0;  //184 / 213 = 0
    16'b10111000_11010110 : OUT <= 0;  //184 / 214 = 0
    16'b10111000_11010111 : OUT <= 0;  //184 / 215 = 0
    16'b10111000_11011000 : OUT <= 0;  //184 / 216 = 0
    16'b10111000_11011001 : OUT <= 0;  //184 / 217 = 0
    16'b10111000_11011010 : OUT <= 0;  //184 / 218 = 0
    16'b10111000_11011011 : OUT <= 0;  //184 / 219 = 0
    16'b10111000_11011100 : OUT <= 0;  //184 / 220 = 0
    16'b10111000_11011101 : OUT <= 0;  //184 / 221 = 0
    16'b10111000_11011110 : OUT <= 0;  //184 / 222 = 0
    16'b10111000_11011111 : OUT <= 0;  //184 / 223 = 0
    16'b10111000_11100000 : OUT <= 0;  //184 / 224 = 0
    16'b10111000_11100001 : OUT <= 0;  //184 / 225 = 0
    16'b10111000_11100010 : OUT <= 0;  //184 / 226 = 0
    16'b10111000_11100011 : OUT <= 0;  //184 / 227 = 0
    16'b10111000_11100100 : OUT <= 0;  //184 / 228 = 0
    16'b10111000_11100101 : OUT <= 0;  //184 / 229 = 0
    16'b10111000_11100110 : OUT <= 0;  //184 / 230 = 0
    16'b10111000_11100111 : OUT <= 0;  //184 / 231 = 0
    16'b10111000_11101000 : OUT <= 0;  //184 / 232 = 0
    16'b10111000_11101001 : OUT <= 0;  //184 / 233 = 0
    16'b10111000_11101010 : OUT <= 0;  //184 / 234 = 0
    16'b10111000_11101011 : OUT <= 0;  //184 / 235 = 0
    16'b10111000_11101100 : OUT <= 0;  //184 / 236 = 0
    16'b10111000_11101101 : OUT <= 0;  //184 / 237 = 0
    16'b10111000_11101110 : OUT <= 0;  //184 / 238 = 0
    16'b10111000_11101111 : OUT <= 0;  //184 / 239 = 0
    16'b10111000_11110000 : OUT <= 0;  //184 / 240 = 0
    16'b10111000_11110001 : OUT <= 0;  //184 / 241 = 0
    16'b10111000_11110010 : OUT <= 0;  //184 / 242 = 0
    16'b10111000_11110011 : OUT <= 0;  //184 / 243 = 0
    16'b10111000_11110100 : OUT <= 0;  //184 / 244 = 0
    16'b10111000_11110101 : OUT <= 0;  //184 / 245 = 0
    16'b10111000_11110110 : OUT <= 0;  //184 / 246 = 0
    16'b10111000_11110111 : OUT <= 0;  //184 / 247 = 0
    16'b10111000_11111000 : OUT <= 0;  //184 / 248 = 0
    16'b10111000_11111001 : OUT <= 0;  //184 / 249 = 0
    16'b10111000_11111010 : OUT <= 0;  //184 / 250 = 0
    16'b10111000_11111011 : OUT <= 0;  //184 / 251 = 0
    16'b10111000_11111100 : OUT <= 0;  //184 / 252 = 0
    16'b10111000_11111101 : OUT <= 0;  //184 / 253 = 0
    16'b10111000_11111110 : OUT <= 0;  //184 / 254 = 0
    16'b10111000_11111111 : OUT <= 0;  //184 / 255 = 0
    16'b10111001_00000000 : OUT <= 0;  //185 / 0 = 0
    16'b10111001_00000001 : OUT <= 185;  //185 / 1 = 185
    16'b10111001_00000010 : OUT <= 92;  //185 / 2 = 92
    16'b10111001_00000011 : OUT <= 61;  //185 / 3 = 61
    16'b10111001_00000100 : OUT <= 46;  //185 / 4 = 46
    16'b10111001_00000101 : OUT <= 37;  //185 / 5 = 37
    16'b10111001_00000110 : OUT <= 30;  //185 / 6 = 30
    16'b10111001_00000111 : OUT <= 26;  //185 / 7 = 26
    16'b10111001_00001000 : OUT <= 23;  //185 / 8 = 23
    16'b10111001_00001001 : OUT <= 20;  //185 / 9 = 20
    16'b10111001_00001010 : OUT <= 18;  //185 / 10 = 18
    16'b10111001_00001011 : OUT <= 16;  //185 / 11 = 16
    16'b10111001_00001100 : OUT <= 15;  //185 / 12 = 15
    16'b10111001_00001101 : OUT <= 14;  //185 / 13 = 14
    16'b10111001_00001110 : OUT <= 13;  //185 / 14 = 13
    16'b10111001_00001111 : OUT <= 12;  //185 / 15 = 12
    16'b10111001_00010000 : OUT <= 11;  //185 / 16 = 11
    16'b10111001_00010001 : OUT <= 10;  //185 / 17 = 10
    16'b10111001_00010010 : OUT <= 10;  //185 / 18 = 10
    16'b10111001_00010011 : OUT <= 9;  //185 / 19 = 9
    16'b10111001_00010100 : OUT <= 9;  //185 / 20 = 9
    16'b10111001_00010101 : OUT <= 8;  //185 / 21 = 8
    16'b10111001_00010110 : OUT <= 8;  //185 / 22 = 8
    16'b10111001_00010111 : OUT <= 8;  //185 / 23 = 8
    16'b10111001_00011000 : OUT <= 7;  //185 / 24 = 7
    16'b10111001_00011001 : OUT <= 7;  //185 / 25 = 7
    16'b10111001_00011010 : OUT <= 7;  //185 / 26 = 7
    16'b10111001_00011011 : OUT <= 6;  //185 / 27 = 6
    16'b10111001_00011100 : OUT <= 6;  //185 / 28 = 6
    16'b10111001_00011101 : OUT <= 6;  //185 / 29 = 6
    16'b10111001_00011110 : OUT <= 6;  //185 / 30 = 6
    16'b10111001_00011111 : OUT <= 5;  //185 / 31 = 5
    16'b10111001_00100000 : OUT <= 5;  //185 / 32 = 5
    16'b10111001_00100001 : OUT <= 5;  //185 / 33 = 5
    16'b10111001_00100010 : OUT <= 5;  //185 / 34 = 5
    16'b10111001_00100011 : OUT <= 5;  //185 / 35 = 5
    16'b10111001_00100100 : OUT <= 5;  //185 / 36 = 5
    16'b10111001_00100101 : OUT <= 5;  //185 / 37 = 5
    16'b10111001_00100110 : OUT <= 4;  //185 / 38 = 4
    16'b10111001_00100111 : OUT <= 4;  //185 / 39 = 4
    16'b10111001_00101000 : OUT <= 4;  //185 / 40 = 4
    16'b10111001_00101001 : OUT <= 4;  //185 / 41 = 4
    16'b10111001_00101010 : OUT <= 4;  //185 / 42 = 4
    16'b10111001_00101011 : OUT <= 4;  //185 / 43 = 4
    16'b10111001_00101100 : OUT <= 4;  //185 / 44 = 4
    16'b10111001_00101101 : OUT <= 4;  //185 / 45 = 4
    16'b10111001_00101110 : OUT <= 4;  //185 / 46 = 4
    16'b10111001_00101111 : OUT <= 3;  //185 / 47 = 3
    16'b10111001_00110000 : OUT <= 3;  //185 / 48 = 3
    16'b10111001_00110001 : OUT <= 3;  //185 / 49 = 3
    16'b10111001_00110010 : OUT <= 3;  //185 / 50 = 3
    16'b10111001_00110011 : OUT <= 3;  //185 / 51 = 3
    16'b10111001_00110100 : OUT <= 3;  //185 / 52 = 3
    16'b10111001_00110101 : OUT <= 3;  //185 / 53 = 3
    16'b10111001_00110110 : OUT <= 3;  //185 / 54 = 3
    16'b10111001_00110111 : OUT <= 3;  //185 / 55 = 3
    16'b10111001_00111000 : OUT <= 3;  //185 / 56 = 3
    16'b10111001_00111001 : OUT <= 3;  //185 / 57 = 3
    16'b10111001_00111010 : OUT <= 3;  //185 / 58 = 3
    16'b10111001_00111011 : OUT <= 3;  //185 / 59 = 3
    16'b10111001_00111100 : OUT <= 3;  //185 / 60 = 3
    16'b10111001_00111101 : OUT <= 3;  //185 / 61 = 3
    16'b10111001_00111110 : OUT <= 2;  //185 / 62 = 2
    16'b10111001_00111111 : OUT <= 2;  //185 / 63 = 2
    16'b10111001_01000000 : OUT <= 2;  //185 / 64 = 2
    16'b10111001_01000001 : OUT <= 2;  //185 / 65 = 2
    16'b10111001_01000010 : OUT <= 2;  //185 / 66 = 2
    16'b10111001_01000011 : OUT <= 2;  //185 / 67 = 2
    16'b10111001_01000100 : OUT <= 2;  //185 / 68 = 2
    16'b10111001_01000101 : OUT <= 2;  //185 / 69 = 2
    16'b10111001_01000110 : OUT <= 2;  //185 / 70 = 2
    16'b10111001_01000111 : OUT <= 2;  //185 / 71 = 2
    16'b10111001_01001000 : OUT <= 2;  //185 / 72 = 2
    16'b10111001_01001001 : OUT <= 2;  //185 / 73 = 2
    16'b10111001_01001010 : OUT <= 2;  //185 / 74 = 2
    16'b10111001_01001011 : OUT <= 2;  //185 / 75 = 2
    16'b10111001_01001100 : OUT <= 2;  //185 / 76 = 2
    16'b10111001_01001101 : OUT <= 2;  //185 / 77 = 2
    16'b10111001_01001110 : OUT <= 2;  //185 / 78 = 2
    16'b10111001_01001111 : OUT <= 2;  //185 / 79 = 2
    16'b10111001_01010000 : OUT <= 2;  //185 / 80 = 2
    16'b10111001_01010001 : OUT <= 2;  //185 / 81 = 2
    16'b10111001_01010010 : OUT <= 2;  //185 / 82 = 2
    16'b10111001_01010011 : OUT <= 2;  //185 / 83 = 2
    16'b10111001_01010100 : OUT <= 2;  //185 / 84 = 2
    16'b10111001_01010101 : OUT <= 2;  //185 / 85 = 2
    16'b10111001_01010110 : OUT <= 2;  //185 / 86 = 2
    16'b10111001_01010111 : OUT <= 2;  //185 / 87 = 2
    16'b10111001_01011000 : OUT <= 2;  //185 / 88 = 2
    16'b10111001_01011001 : OUT <= 2;  //185 / 89 = 2
    16'b10111001_01011010 : OUT <= 2;  //185 / 90 = 2
    16'b10111001_01011011 : OUT <= 2;  //185 / 91 = 2
    16'b10111001_01011100 : OUT <= 2;  //185 / 92 = 2
    16'b10111001_01011101 : OUT <= 1;  //185 / 93 = 1
    16'b10111001_01011110 : OUT <= 1;  //185 / 94 = 1
    16'b10111001_01011111 : OUT <= 1;  //185 / 95 = 1
    16'b10111001_01100000 : OUT <= 1;  //185 / 96 = 1
    16'b10111001_01100001 : OUT <= 1;  //185 / 97 = 1
    16'b10111001_01100010 : OUT <= 1;  //185 / 98 = 1
    16'b10111001_01100011 : OUT <= 1;  //185 / 99 = 1
    16'b10111001_01100100 : OUT <= 1;  //185 / 100 = 1
    16'b10111001_01100101 : OUT <= 1;  //185 / 101 = 1
    16'b10111001_01100110 : OUT <= 1;  //185 / 102 = 1
    16'b10111001_01100111 : OUT <= 1;  //185 / 103 = 1
    16'b10111001_01101000 : OUT <= 1;  //185 / 104 = 1
    16'b10111001_01101001 : OUT <= 1;  //185 / 105 = 1
    16'b10111001_01101010 : OUT <= 1;  //185 / 106 = 1
    16'b10111001_01101011 : OUT <= 1;  //185 / 107 = 1
    16'b10111001_01101100 : OUT <= 1;  //185 / 108 = 1
    16'b10111001_01101101 : OUT <= 1;  //185 / 109 = 1
    16'b10111001_01101110 : OUT <= 1;  //185 / 110 = 1
    16'b10111001_01101111 : OUT <= 1;  //185 / 111 = 1
    16'b10111001_01110000 : OUT <= 1;  //185 / 112 = 1
    16'b10111001_01110001 : OUT <= 1;  //185 / 113 = 1
    16'b10111001_01110010 : OUT <= 1;  //185 / 114 = 1
    16'b10111001_01110011 : OUT <= 1;  //185 / 115 = 1
    16'b10111001_01110100 : OUT <= 1;  //185 / 116 = 1
    16'b10111001_01110101 : OUT <= 1;  //185 / 117 = 1
    16'b10111001_01110110 : OUT <= 1;  //185 / 118 = 1
    16'b10111001_01110111 : OUT <= 1;  //185 / 119 = 1
    16'b10111001_01111000 : OUT <= 1;  //185 / 120 = 1
    16'b10111001_01111001 : OUT <= 1;  //185 / 121 = 1
    16'b10111001_01111010 : OUT <= 1;  //185 / 122 = 1
    16'b10111001_01111011 : OUT <= 1;  //185 / 123 = 1
    16'b10111001_01111100 : OUT <= 1;  //185 / 124 = 1
    16'b10111001_01111101 : OUT <= 1;  //185 / 125 = 1
    16'b10111001_01111110 : OUT <= 1;  //185 / 126 = 1
    16'b10111001_01111111 : OUT <= 1;  //185 / 127 = 1
    16'b10111001_10000000 : OUT <= 1;  //185 / 128 = 1
    16'b10111001_10000001 : OUT <= 1;  //185 / 129 = 1
    16'b10111001_10000010 : OUT <= 1;  //185 / 130 = 1
    16'b10111001_10000011 : OUT <= 1;  //185 / 131 = 1
    16'b10111001_10000100 : OUT <= 1;  //185 / 132 = 1
    16'b10111001_10000101 : OUT <= 1;  //185 / 133 = 1
    16'b10111001_10000110 : OUT <= 1;  //185 / 134 = 1
    16'b10111001_10000111 : OUT <= 1;  //185 / 135 = 1
    16'b10111001_10001000 : OUT <= 1;  //185 / 136 = 1
    16'b10111001_10001001 : OUT <= 1;  //185 / 137 = 1
    16'b10111001_10001010 : OUT <= 1;  //185 / 138 = 1
    16'b10111001_10001011 : OUT <= 1;  //185 / 139 = 1
    16'b10111001_10001100 : OUT <= 1;  //185 / 140 = 1
    16'b10111001_10001101 : OUT <= 1;  //185 / 141 = 1
    16'b10111001_10001110 : OUT <= 1;  //185 / 142 = 1
    16'b10111001_10001111 : OUT <= 1;  //185 / 143 = 1
    16'b10111001_10010000 : OUT <= 1;  //185 / 144 = 1
    16'b10111001_10010001 : OUT <= 1;  //185 / 145 = 1
    16'b10111001_10010010 : OUT <= 1;  //185 / 146 = 1
    16'b10111001_10010011 : OUT <= 1;  //185 / 147 = 1
    16'b10111001_10010100 : OUT <= 1;  //185 / 148 = 1
    16'b10111001_10010101 : OUT <= 1;  //185 / 149 = 1
    16'b10111001_10010110 : OUT <= 1;  //185 / 150 = 1
    16'b10111001_10010111 : OUT <= 1;  //185 / 151 = 1
    16'b10111001_10011000 : OUT <= 1;  //185 / 152 = 1
    16'b10111001_10011001 : OUT <= 1;  //185 / 153 = 1
    16'b10111001_10011010 : OUT <= 1;  //185 / 154 = 1
    16'b10111001_10011011 : OUT <= 1;  //185 / 155 = 1
    16'b10111001_10011100 : OUT <= 1;  //185 / 156 = 1
    16'b10111001_10011101 : OUT <= 1;  //185 / 157 = 1
    16'b10111001_10011110 : OUT <= 1;  //185 / 158 = 1
    16'b10111001_10011111 : OUT <= 1;  //185 / 159 = 1
    16'b10111001_10100000 : OUT <= 1;  //185 / 160 = 1
    16'b10111001_10100001 : OUT <= 1;  //185 / 161 = 1
    16'b10111001_10100010 : OUT <= 1;  //185 / 162 = 1
    16'b10111001_10100011 : OUT <= 1;  //185 / 163 = 1
    16'b10111001_10100100 : OUT <= 1;  //185 / 164 = 1
    16'b10111001_10100101 : OUT <= 1;  //185 / 165 = 1
    16'b10111001_10100110 : OUT <= 1;  //185 / 166 = 1
    16'b10111001_10100111 : OUT <= 1;  //185 / 167 = 1
    16'b10111001_10101000 : OUT <= 1;  //185 / 168 = 1
    16'b10111001_10101001 : OUT <= 1;  //185 / 169 = 1
    16'b10111001_10101010 : OUT <= 1;  //185 / 170 = 1
    16'b10111001_10101011 : OUT <= 1;  //185 / 171 = 1
    16'b10111001_10101100 : OUT <= 1;  //185 / 172 = 1
    16'b10111001_10101101 : OUT <= 1;  //185 / 173 = 1
    16'b10111001_10101110 : OUT <= 1;  //185 / 174 = 1
    16'b10111001_10101111 : OUT <= 1;  //185 / 175 = 1
    16'b10111001_10110000 : OUT <= 1;  //185 / 176 = 1
    16'b10111001_10110001 : OUT <= 1;  //185 / 177 = 1
    16'b10111001_10110010 : OUT <= 1;  //185 / 178 = 1
    16'b10111001_10110011 : OUT <= 1;  //185 / 179 = 1
    16'b10111001_10110100 : OUT <= 1;  //185 / 180 = 1
    16'b10111001_10110101 : OUT <= 1;  //185 / 181 = 1
    16'b10111001_10110110 : OUT <= 1;  //185 / 182 = 1
    16'b10111001_10110111 : OUT <= 1;  //185 / 183 = 1
    16'b10111001_10111000 : OUT <= 1;  //185 / 184 = 1
    16'b10111001_10111001 : OUT <= 1;  //185 / 185 = 1
    16'b10111001_10111010 : OUT <= 0;  //185 / 186 = 0
    16'b10111001_10111011 : OUT <= 0;  //185 / 187 = 0
    16'b10111001_10111100 : OUT <= 0;  //185 / 188 = 0
    16'b10111001_10111101 : OUT <= 0;  //185 / 189 = 0
    16'b10111001_10111110 : OUT <= 0;  //185 / 190 = 0
    16'b10111001_10111111 : OUT <= 0;  //185 / 191 = 0
    16'b10111001_11000000 : OUT <= 0;  //185 / 192 = 0
    16'b10111001_11000001 : OUT <= 0;  //185 / 193 = 0
    16'b10111001_11000010 : OUT <= 0;  //185 / 194 = 0
    16'b10111001_11000011 : OUT <= 0;  //185 / 195 = 0
    16'b10111001_11000100 : OUT <= 0;  //185 / 196 = 0
    16'b10111001_11000101 : OUT <= 0;  //185 / 197 = 0
    16'b10111001_11000110 : OUT <= 0;  //185 / 198 = 0
    16'b10111001_11000111 : OUT <= 0;  //185 / 199 = 0
    16'b10111001_11001000 : OUT <= 0;  //185 / 200 = 0
    16'b10111001_11001001 : OUT <= 0;  //185 / 201 = 0
    16'b10111001_11001010 : OUT <= 0;  //185 / 202 = 0
    16'b10111001_11001011 : OUT <= 0;  //185 / 203 = 0
    16'b10111001_11001100 : OUT <= 0;  //185 / 204 = 0
    16'b10111001_11001101 : OUT <= 0;  //185 / 205 = 0
    16'b10111001_11001110 : OUT <= 0;  //185 / 206 = 0
    16'b10111001_11001111 : OUT <= 0;  //185 / 207 = 0
    16'b10111001_11010000 : OUT <= 0;  //185 / 208 = 0
    16'b10111001_11010001 : OUT <= 0;  //185 / 209 = 0
    16'b10111001_11010010 : OUT <= 0;  //185 / 210 = 0
    16'b10111001_11010011 : OUT <= 0;  //185 / 211 = 0
    16'b10111001_11010100 : OUT <= 0;  //185 / 212 = 0
    16'b10111001_11010101 : OUT <= 0;  //185 / 213 = 0
    16'b10111001_11010110 : OUT <= 0;  //185 / 214 = 0
    16'b10111001_11010111 : OUT <= 0;  //185 / 215 = 0
    16'b10111001_11011000 : OUT <= 0;  //185 / 216 = 0
    16'b10111001_11011001 : OUT <= 0;  //185 / 217 = 0
    16'b10111001_11011010 : OUT <= 0;  //185 / 218 = 0
    16'b10111001_11011011 : OUT <= 0;  //185 / 219 = 0
    16'b10111001_11011100 : OUT <= 0;  //185 / 220 = 0
    16'b10111001_11011101 : OUT <= 0;  //185 / 221 = 0
    16'b10111001_11011110 : OUT <= 0;  //185 / 222 = 0
    16'b10111001_11011111 : OUT <= 0;  //185 / 223 = 0
    16'b10111001_11100000 : OUT <= 0;  //185 / 224 = 0
    16'b10111001_11100001 : OUT <= 0;  //185 / 225 = 0
    16'b10111001_11100010 : OUT <= 0;  //185 / 226 = 0
    16'b10111001_11100011 : OUT <= 0;  //185 / 227 = 0
    16'b10111001_11100100 : OUT <= 0;  //185 / 228 = 0
    16'b10111001_11100101 : OUT <= 0;  //185 / 229 = 0
    16'b10111001_11100110 : OUT <= 0;  //185 / 230 = 0
    16'b10111001_11100111 : OUT <= 0;  //185 / 231 = 0
    16'b10111001_11101000 : OUT <= 0;  //185 / 232 = 0
    16'b10111001_11101001 : OUT <= 0;  //185 / 233 = 0
    16'b10111001_11101010 : OUT <= 0;  //185 / 234 = 0
    16'b10111001_11101011 : OUT <= 0;  //185 / 235 = 0
    16'b10111001_11101100 : OUT <= 0;  //185 / 236 = 0
    16'b10111001_11101101 : OUT <= 0;  //185 / 237 = 0
    16'b10111001_11101110 : OUT <= 0;  //185 / 238 = 0
    16'b10111001_11101111 : OUT <= 0;  //185 / 239 = 0
    16'b10111001_11110000 : OUT <= 0;  //185 / 240 = 0
    16'b10111001_11110001 : OUT <= 0;  //185 / 241 = 0
    16'b10111001_11110010 : OUT <= 0;  //185 / 242 = 0
    16'b10111001_11110011 : OUT <= 0;  //185 / 243 = 0
    16'b10111001_11110100 : OUT <= 0;  //185 / 244 = 0
    16'b10111001_11110101 : OUT <= 0;  //185 / 245 = 0
    16'b10111001_11110110 : OUT <= 0;  //185 / 246 = 0
    16'b10111001_11110111 : OUT <= 0;  //185 / 247 = 0
    16'b10111001_11111000 : OUT <= 0;  //185 / 248 = 0
    16'b10111001_11111001 : OUT <= 0;  //185 / 249 = 0
    16'b10111001_11111010 : OUT <= 0;  //185 / 250 = 0
    16'b10111001_11111011 : OUT <= 0;  //185 / 251 = 0
    16'b10111001_11111100 : OUT <= 0;  //185 / 252 = 0
    16'b10111001_11111101 : OUT <= 0;  //185 / 253 = 0
    16'b10111001_11111110 : OUT <= 0;  //185 / 254 = 0
    16'b10111001_11111111 : OUT <= 0;  //185 / 255 = 0
    16'b10111010_00000000 : OUT <= 0;  //186 / 0 = 0
    16'b10111010_00000001 : OUT <= 186;  //186 / 1 = 186
    16'b10111010_00000010 : OUT <= 93;  //186 / 2 = 93
    16'b10111010_00000011 : OUT <= 62;  //186 / 3 = 62
    16'b10111010_00000100 : OUT <= 46;  //186 / 4 = 46
    16'b10111010_00000101 : OUT <= 37;  //186 / 5 = 37
    16'b10111010_00000110 : OUT <= 31;  //186 / 6 = 31
    16'b10111010_00000111 : OUT <= 26;  //186 / 7 = 26
    16'b10111010_00001000 : OUT <= 23;  //186 / 8 = 23
    16'b10111010_00001001 : OUT <= 20;  //186 / 9 = 20
    16'b10111010_00001010 : OUT <= 18;  //186 / 10 = 18
    16'b10111010_00001011 : OUT <= 16;  //186 / 11 = 16
    16'b10111010_00001100 : OUT <= 15;  //186 / 12 = 15
    16'b10111010_00001101 : OUT <= 14;  //186 / 13 = 14
    16'b10111010_00001110 : OUT <= 13;  //186 / 14 = 13
    16'b10111010_00001111 : OUT <= 12;  //186 / 15 = 12
    16'b10111010_00010000 : OUT <= 11;  //186 / 16 = 11
    16'b10111010_00010001 : OUT <= 10;  //186 / 17 = 10
    16'b10111010_00010010 : OUT <= 10;  //186 / 18 = 10
    16'b10111010_00010011 : OUT <= 9;  //186 / 19 = 9
    16'b10111010_00010100 : OUT <= 9;  //186 / 20 = 9
    16'b10111010_00010101 : OUT <= 8;  //186 / 21 = 8
    16'b10111010_00010110 : OUT <= 8;  //186 / 22 = 8
    16'b10111010_00010111 : OUT <= 8;  //186 / 23 = 8
    16'b10111010_00011000 : OUT <= 7;  //186 / 24 = 7
    16'b10111010_00011001 : OUT <= 7;  //186 / 25 = 7
    16'b10111010_00011010 : OUT <= 7;  //186 / 26 = 7
    16'b10111010_00011011 : OUT <= 6;  //186 / 27 = 6
    16'b10111010_00011100 : OUT <= 6;  //186 / 28 = 6
    16'b10111010_00011101 : OUT <= 6;  //186 / 29 = 6
    16'b10111010_00011110 : OUT <= 6;  //186 / 30 = 6
    16'b10111010_00011111 : OUT <= 6;  //186 / 31 = 6
    16'b10111010_00100000 : OUT <= 5;  //186 / 32 = 5
    16'b10111010_00100001 : OUT <= 5;  //186 / 33 = 5
    16'b10111010_00100010 : OUT <= 5;  //186 / 34 = 5
    16'b10111010_00100011 : OUT <= 5;  //186 / 35 = 5
    16'b10111010_00100100 : OUT <= 5;  //186 / 36 = 5
    16'b10111010_00100101 : OUT <= 5;  //186 / 37 = 5
    16'b10111010_00100110 : OUT <= 4;  //186 / 38 = 4
    16'b10111010_00100111 : OUT <= 4;  //186 / 39 = 4
    16'b10111010_00101000 : OUT <= 4;  //186 / 40 = 4
    16'b10111010_00101001 : OUT <= 4;  //186 / 41 = 4
    16'b10111010_00101010 : OUT <= 4;  //186 / 42 = 4
    16'b10111010_00101011 : OUT <= 4;  //186 / 43 = 4
    16'b10111010_00101100 : OUT <= 4;  //186 / 44 = 4
    16'b10111010_00101101 : OUT <= 4;  //186 / 45 = 4
    16'b10111010_00101110 : OUT <= 4;  //186 / 46 = 4
    16'b10111010_00101111 : OUT <= 3;  //186 / 47 = 3
    16'b10111010_00110000 : OUT <= 3;  //186 / 48 = 3
    16'b10111010_00110001 : OUT <= 3;  //186 / 49 = 3
    16'b10111010_00110010 : OUT <= 3;  //186 / 50 = 3
    16'b10111010_00110011 : OUT <= 3;  //186 / 51 = 3
    16'b10111010_00110100 : OUT <= 3;  //186 / 52 = 3
    16'b10111010_00110101 : OUT <= 3;  //186 / 53 = 3
    16'b10111010_00110110 : OUT <= 3;  //186 / 54 = 3
    16'b10111010_00110111 : OUT <= 3;  //186 / 55 = 3
    16'b10111010_00111000 : OUT <= 3;  //186 / 56 = 3
    16'b10111010_00111001 : OUT <= 3;  //186 / 57 = 3
    16'b10111010_00111010 : OUT <= 3;  //186 / 58 = 3
    16'b10111010_00111011 : OUT <= 3;  //186 / 59 = 3
    16'b10111010_00111100 : OUT <= 3;  //186 / 60 = 3
    16'b10111010_00111101 : OUT <= 3;  //186 / 61 = 3
    16'b10111010_00111110 : OUT <= 3;  //186 / 62 = 3
    16'b10111010_00111111 : OUT <= 2;  //186 / 63 = 2
    16'b10111010_01000000 : OUT <= 2;  //186 / 64 = 2
    16'b10111010_01000001 : OUT <= 2;  //186 / 65 = 2
    16'b10111010_01000010 : OUT <= 2;  //186 / 66 = 2
    16'b10111010_01000011 : OUT <= 2;  //186 / 67 = 2
    16'b10111010_01000100 : OUT <= 2;  //186 / 68 = 2
    16'b10111010_01000101 : OUT <= 2;  //186 / 69 = 2
    16'b10111010_01000110 : OUT <= 2;  //186 / 70 = 2
    16'b10111010_01000111 : OUT <= 2;  //186 / 71 = 2
    16'b10111010_01001000 : OUT <= 2;  //186 / 72 = 2
    16'b10111010_01001001 : OUT <= 2;  //186 / 73 = 2
    16'b10111010_01001010 : OUT <= 2;  //186 / 74 = 2
    16'b10111010_01001011 : OUT <= 2;  //186 / 75 = 2
    16'b10111010_01001100 : OUT <= 2;  //186 / 76 = 2
    16'b10111010_01001101 : OUT <= 2;  //186 / 77 = 2
    16'b10111010_01001110 : OUT <= 2;  //186 / 78 = 2
    16'b10111010_01001111 : OUT <= 2;  //186 / 79 = 2
    16'b10111010_01010000 : OUT <= 2;  //186 / 80 = 2
    16'b10111010_01010001 : OUT <= 2;  //186 / 81 = 2
    16'b10111010_01010010 : OUT <= 2;  //186 / 82 = 2
    16'b10111010_01010011 : OUT <= 2;  //186 / 83 = 2
    16'b10111010_01010100 : OUT <= 2;  //186 / 84 = 2
    16'b10111010_01010101 : OUT <= 2;  //186 / 85 = 2
    16'b10111010_01010110 : OUT <= 2;  //186 / 86 = 2
    16'b10111010_01010111 : OUT <= 2;  //186 / 87 = 2
    16'b10111010_01011000 : OUT <= 2;  //186 / 88 = 2
    16'b10111010_01011001 : OUT <= 2;  //186 / 89 = 2
    16'b10111010_01011010 : OUT <= 2;  //186 / 90 = 2
    16'b10111010_01011011 : OUT <= 2;  //186 / 91 = 2
    16'b10111010_01011100 : OUT <= 2;  //186 / 92 = 2
    16'b10111010_01011101 : OUT <= 2;  //186 / 93 = 2
    16'b10111010_01011110 : OUT <= 1;  //186 / 94 = 1
    16'b10111010_01011111 : OUT <= 1;  //186 / 95 = 1
    16'b10111010_01100000 : OUT <= 1;  //186 / 96 = 1
    16'b10111010_01100001 : OUT <= 1;  //186 / 97 = 1
    16'b10111010_01100010 : OUT <= 1;  //186 / 98 = 1
    16'b10111010_01100011 : OUT <= 1;  //186 / 99 = 1
    16'b10111010_01100100 : OUT <= 1;  //186 / 100 = 1
    16'b10111010_01100101 : OUT <= 1;  //186 / 101 = 1
    16'b10111010_01100110 : OUT <= 1;  //186 / 102 = 1
    16'b10111010_01100111 : OUT <= 1;  //186 / 103 = 1
    16'b10111010_01101000 : OUT <= 1;  //186 / 104 = 1
    16'b10111010_01101001 : OUT <= 1;  //186 / 105 = 1
    16'b10111010_01101010 : OUT <= 1;  //186 / 106 = 1
    16'b10111010_01101011 : OUT <= 1;  //186 / 107 = 1
    16'b10111010_01101100 : OUT <= 1;  //186 / 108 = 1
    16'b10111010_01101101 : OUT <= 1;  //186 / 109 = 1
    16'b10111010_01101110 : OUT <= 1;  //186 / 110 = 1
    16'b10111010_01101111 : OUT <= 1;  //186 / 111 = 1
    16'b10111010_01110000 : OUT <= 1;  //186 / 112 = 1
    16'b10111010_01110001 : OUT <= 1;  //186 / 113 = 1
    16'b10111010_01110010 : OUT <= 1;  //186 / 114 = 1
    16'b10111010_01110011 : OUT <= 1;  //186 / 115 = 1
    16'b10111010_01110100 : OUT <= 1;  //186 / 116 = 1
    16'b10111010_01110101 : OUT <= 1;  //186 / 117 = 1
    16'b10111010_01110110 : OUT <= 1;  //186 / 118 = 1
    16'b10111010_01110111 : OUT <= 1;  //186 / 119 = 1
    16'b10111010_01111000 : OUT <= 1;  //186 / 120 = 1
    16'b10111010_01111001 : OUT <= 1;  //186 / 121 = 1
    16'b10111010_01111010 : OUT <= 1;  //186 / 122 = 1
    16'b10111010_01111011 : OUT <= 1;  //186 / 123 = 1
    16'b10111010_01111100 : OUT <= 1;  //186 / 124 = 1
    16'b10111010_01111101 : OUT <= 1;  //186 / 125 = 1
    16'b10111010_01111110 : OUT <= 1;  //186 / 126 = 1
    16'b10111010_01111111 : OUT <= 1;  //186 / 127 = 1
    16'b10111010_10000000 : OUT <= 1;  //186 / 128 = 1
    16'b10111010_10000001 : OUT <= 1;  //186 / 129 = 1
    16'b10111010_10000010 : OUT <= 1;  //186 / 130 = 1
    16'b10111010_10000011 : OUT <= 1;  //186 / 131 = 1
    16'b10111010_10000100 : OUT <= 1;  //186 / 132 = 1
    16'b10111010_10000101 : OUT <= 1;  //186 / 133 = 1
    16'b10111010_10000110 : OUT <= 1;  //186 / 134 = 1
    16'b10111010_10000111 : OUT <= 1;  //186 / 135 = 1
    16'b10111010_10001000 : OUT <= 1;  //186 / 136 = 1
    16'b10111010_10001001 : OUT <= 1;  //186 / 137 = 1
    16'b10111010_10001010 : OUT <= 1;  //186 / 138 = 1
    16'b10111010_10001011 : OUT <= 1;  //186 / 139 = 1
    16'b10111010_10001100 : OUT <= 1;  //186 / 140 = 1
    16'b10111010_10001101 : OUT <= 1;  //186 / 141 = 1
    16'b10111010_10001110 : OUT <= 1;  //186 / 142 = 1
    16'b10111010_10001111 : OUT <= 1;  //186 / 143 = 1
    16'b10111010_10010000 : OUT <= 1;  //186 / 144 = 1
    16'b10111010_10010001 : OUT <= 1;  //186 / 145 = 1
    16'b10111010_10010010 : OUT <= 1;  //186 / 146 = 1
    16'b10111010_10010011 : OUT <= 1;  //186 / 147 = 1
    16'b10111010_10010100 : OUT <= 1;  //186 / 148 = 1
    16'b10111010_10010101 : OUT <= 1;  //186 / 149 = 1
    16'b10111010_10010110 : OUT <= 1;  //186 / 150 = 1
    16'b10111010_10010111 : OUT <= 1;  //186 / 151 = 1
    16'b10111010_10011000 : OUT <= 1;  //186 / 152 = 1
    16'b10111010_10011001 : OUT <= 1;  //186 / 153 = 1
    16'b10111010_10011010 : OUT <= 1;  //186 / 154 = 1
    16'b10111010_10011011 : OUT <= 1;  //186 / 155 = 1
    16'b10111010_10011100 : OUT <= 1;  //186 / 156 = 1
    16'b10111010_10011101 : OUT <= 1;  //186 / 157 = 1
    16'b10111010_10011110 : OUT <= 1;  //186 / 158 = 1
    16'b10111010_10011111 : OUT <= 1;  //186 / 159 = 1
    16'b10111010_10100000 : OUT <= 1;  //186 / 160 = 1
    16'b10111010_10100001 : OUT <= 1;  //186 / 161 = 1
    16'b10111010_10100010 : OUT <= 1;  //186 / 162 = 1
    16'b10111010_10100011 : OUT <= 1;  //186 / 163 = 1
    16'b10111010_10100100 : OUT <= 1;  //186 / 164 = 1
    16'b10111010_10100101 : OUT <= 1;  //186 / 165 = 1
    16'b10111010_10100110 : OUT <= 1;  //186 / 166 = 1
    16'b10111010_10100111 : OUT <= 1;  //186 / 167 = 1
    16'b10111010_10101000 : OUT <= 1;  //186 / 168 = 1
    16'b10111010_10101001 : OUT <= 1;  //186 / 169 = 1
    16'b10111010_10101010 : OUT <= 1;  //186 / 170 = 1
    16'b10111010_10101011 : OUT <= 1;  //186 / 171 = 1
    16'b10111010_10101100 : OUT <= 1;  //186 / 172 = 1
    16'b10111010_10101101 : OUT <= 1;  //186 / 173 = 1
    16'b10111010_10101110 : OUT <= 1;  //186 / 174 = 1
    16'b10111010_10101111 : OUT <= 1;  //186 / 175 = 1
    16'b10111010_10110000 : OUT <= 1;  //186 / 176 = 1
    16'b10111010_10110001 : OUT <= 1;  //186 / 177 = 1
    16'b10111010_10110010 : OUT <= 1;  //186 / 178 = 1
    16'b10111010_10110011 : OUT <= 1;  //186 / 179 = 1
    16'b10111010_10110100 : OUT <= 1;  //186 / 180 = 1
    16'b10111010_10110101 : OUT <= 1;  //186 / 181 = 1
    16'b10111010_10110110 : OUT <= 1;  //186 / 182 = 1
    16'b10111010_10110111 : OUT <= 1;  //186 / 183 = 1
    16'b10111010_10111000 : OUT <= 1;  //186 / 184 = 1
    16'b10111010_10111001 : OUT <= 1;  //186 / 185 = 1
    16'b10111010_10111010 : OUT <= 1;  //186 / 186 = 1
    16'b10111010_10111011 : OUT <= 0;  //186 / 187 = 0
    16'b10111010_10111100 : OUT <= 0;  //186 / 188 = 0
    16'b10111010_10111101 : OUT <= 0;  //186 / 189 = 0
    16'b10111010_10111110 : OUT <= 0;  //186 / 190 = 0
    16'b10111010_10111111 : OUT <= 0;  //186 / 191 = 0
    16'b10111010_11000000 : OUT <= 0;  //186 / 192 = 0
    16'b10111010_11000001 : OUT <= 0;  //186 / 193 = 0
    16'b10111010_11000010 : OUT <= 0;  //186 / 194 = 0
    16'b10111010_11000011 : OUT <= 0;  //186 / 195 = 0
    16'b10111010_11000100 : OUT <= 0;  //186 / 196 = 0
    16'b10111010_11000101 : OUT <= 0;  //186 / 197 = 0
    16'b10111010_11000110 : OUT <= 0;  //186 / 198 = 0
    16'b10111010_11000111 : OUT <= 0;  //186 / 199 = 0
    16'b10111010_11001000 : OUT <= 0;  //186 / 200 = 0
    16'b10111010_11001001 : OUT <= 0;  //186 / 201 = 0
    16'b10111010_11001010 : OUT <= 0;  //186 / 202 = 0
    16'b10111010_11001011 : OUT <= 0;  //186 / 203 = 0
    16'b10111010_11001100 : OUT <= 0;  //186 / 204 = 0
    16'b10111010_11001101 : OUT <= 0;  //186 / 205 = 0
    16'b10111010_11001110 : OUT <= 0;  //186 / 206 = 0
    16'b10111010_11001111 : OUT <= 0;  //186 / 207 = 0
    16'b10111010_11010000 : OUT <= 0;  //186 / 208 = 0
    16'b10111010_11010001 : OUT <= 0;  //186 / 209 = 0
    16'b10111010_11010010 : OUT <= 0;  //186 / 210 = 0
    16'b10111010_11010011 : OUT <= 0;  //186 / 211 = 0
    16'b10111010_11010100 : OUT <= 0;  //186 / 212 = 0
    16'b10111010_11010101 : OUT <= 0;  //186 / 213 = 0
    16'b10111010_11010110 : OUT <= 0;  //186 / 214 = 0
    16'b10111010_11010111 : OUT <= 0;  //186 / 215 = 0
    16'b10111010_11011000 : OUT <= 0;  //186 / 216 = 0
    16'b10111010_11011001 : OUT <= 0;  //186 / 217 = 0
    16'b10111010_11011010 : OUT <= 0;  //186 / 218 = 0
    16'b10111010_11011011 : OUT <= 0;  //186 / 219 = 0
    16'b10111010_11011100 : OUT <= 0;  //186 / 220 = 0
    16'b10111010_11011101 : OUT <= 0;  //186 / 221 = 0
    16'b10111010_11011110 : OUT <= 0;  //186 / 222 = 0
    16'b10111010_11011111 : OUT <= 0;  //186 / 223 = 0
    16'b10111010_11100000 : OUT <= 0;  //186 / 224 = 0
    16'b10111010_11100001 : OUT <= 0;  //186 / 225 = 0
    16'b10111010_11100010 : OUT <= 0;  //186 / 226 = 0
    16'b10111010_11100011 : OUT <= 0;  //186 / 227 = 0
    16'b10111010_11100100 : OUT <= 0;  //186 / 228 = 0
    16'b10111010_11100101 : OUT <= 0;  //186 / 229 = 0
    16'b10111010_11100110 : OUT <= 0;  //186 / 230 = 0
    16'b10111010_11100111 : OUT <= 0;  //186 / 231 = 0
    16'b10111010_11101000 : OUT <= 0;  //186 / 232 = 0
    16'b10111010_11101001 : OUT <= 0;  //186 / 233 = 0
    16'b10111010_11101010 : OUT <= 0;  //186 / 234 = 0
    16'b10111010_11101011 : OUT <= 0;  //186 / 235 = 0
    16'b10111010_11101100 : OUT <= 0;  //186 / 236 = 0
    16'b10111010_11101101 : OUT <= 0;  //186 / 237 = 0
    16'b10111010_11101110 : OUT <= 0;  //186 / 238 = 0
    16'b10111010_11101111 : OUT <= 0;  //186 / 239 = 0
    16'b10111010_11110000 : OUT <= 0;  //186 / 240 = 0
    16'b10111010_11110001 : OUT <= 0;  //186 / 241 = 0
    16'b10111010_11110010 : OUT <= 0;  //186 / 242 = 0
    16'b10111010_11110011 : OUT <= 0;  //186 / 243 = 0
    16'b10111010_11110100 : OUT <= 0;  //186 / 244 = 0
    16'b10111010_11110101 : OUT <= 0;  //186 / 245 = 0
    16'b10111010_11110110 : OUT <= 0;  //186 / 246 = 0
    16'b10111010_11110111 : OUT <= 0;  //186 / 247 = 0
    16'b10111010_11111000 : OUT <= 0;  //186 / 248 = 0
    16'b10111010_11111001 : OUT <= 0;  //186 / 249 = 0
    16'b10111010_11111010 : OUT <= 0;  //186 / 250 = 0
    16'b10111010_11111011 : OUT <= 0;  //186 / 251 = 0
    16'b10111010_11111100 : OUT <= 0;  //186 / 252 = 0
    16'b10111010_11111101 : OUT <= 0;  //186 / 253 = 0
    16'b10111010_11111110 : OUT <= 0;  //186 / 254 = 0
    16'b10111010_11111111 : OUT <= 0;  //186 / 255 = 0
    16'b10111011_00000000 : OUT <= 0;  //187 / 0 = 0
    16'b10111011_00000001 : OUT <= 187;  //187 / 1 = 187
    16'b10111011_00000010 : OUT <= 93;  //187 / 2 = 93
    16'b10111011_00000011 : OUT <= 62;  //187 / 3 = 62
    16'b10111011_00000100 : OUT <= 46;  //187 / 4 = 46
    16'b10111011_00000101 : OUT <= 37;  //187 / 5 = 37
    16'b10111011_00000110 : OUT <= 31;  //187 / 6 = 31
    16'b10111011_00000111 : OUT <= 26;  //187 / 7 = 26
    16'b10111011_00001000 : OUT <= 23;  //187 / 8 = 23
    16'b10111011_00001001 : OUT <= 20;  //187 / 9 = 20
    16'b10111011_00001010 : OUT <= 18;  //187 / 10 = 18
    16'b10111011_00001011 : OUT <= 17;  //187 / 11 = 17
    16'b10111011_00001100 : OUT <= 15;  //187 / 12 = 15
    16'b10111011_00001101 : OUT <= 14;  //187 / 13 = 14
    16'b10111011_00001110 : OUT <= 13;  //187 / 14 = 13
    16'b10111011_00001111 : OUT <= 12;  //187 / 15 = 12
    16'b10111011_00010000 : OUT <= 11;  //187 / 16 = 11
    16'b10111011_00010001 : OUT <= 11;  //187 / 17 = 11
    16'b10111011_00010010 : OUT <= 10;  //187 / 18 = 10
    16'b10111011_00010011 : OUT <= 9;  //187 / 19 = 9
    16'b10111011_00010100 : OUT <= 9;  //187 / 20 = 9
    16'b10111011_00010101 : OUT <= 8;  //187 / 21 = 8
    16'b10111011_00010110 : OUT <= 8;  //187 / 22 = 8
    16'b10111011_00010111 : OUT <= 8;  //187 / 23 = 8
    16'b10111011_00011000 : OUT <= 7;  //187 / 24 = 7
    16'b10111011_00011001 : OUT <= 7;  //187 / 25 = 7
    16'b10111011_00011010 : OUT <= 7;  //187 / 26 = 7
    16'b10111011_00011011 : OUT <= 6;  //187 / 27 = 6
    16'b10111011_00011100 : OUT <= 6;  //187 / 28 = 6
    16'b10111011_00011101 : OUT <= 6;  //187 / 29 = 6
    16'b10111011_00011110 : OUT <= 6;  //187 / 30 = 6
    16'b10111011_00011111 : OUT <= 6;  //187 / 31 = 6
    16'b10111011_00100000 : OUT <= 5;  //187 / 32 = 5
    16'b10111011_00100001 : OUT <= 5;  //187 / 33 = 5
    16'b10111011_00100010 : OUT <= 5;  //187 / 34 = 5
    16'b10111011_00100011 : OUT <= 5;  //187 / 35 = 5
    16'b10111011_00100100 : OUT <= 5;  //187 / 36 = 5
    16'b10111011_00100101 : OUT <= 5;  //187 / 37 = 5
    16'b10111011_00100110 : OUT <= 4;  //187 / 38 = 4
    16'b10111011_00100111 : OUT <= 4;  //187 / 39 = 4
    16'b10111011_00101000 : OUT <= 4;  //187 / 40 = 4
    16'b10111011_00101001 : OUT <= 4;  //187 / 41 = 4
    16'b10111011_00101010 : OUT <= 4;  //187 / 42 = 4
    16'b10111011_00101011 : OUT <= 4;  //187 / 43 = 4
    16'b10111011_00101100 : OUT <= 4;  //187 / 44 = 4
    16'b10111011_00101101 : OUT <= 4;  //187 / 45 = 4
    16'b10111011_00101110 : OUT <= 4;  //187 / 46 = 4
    16'b10111011_00101111 : OUT <= 3;  //187 / 47 = 3
    16'b10111011_00110000 : OUT <= 3;  //187 / 48 = 3
    16'b10111011_00110001 : OUT <= 3;  //187 / 49 = 3
    16'b10111011_00110010 : OUT <= 3;  //187 / 50 = 3
    16'b10111011_00110011 : OUT <= 3;  //187 / 51 = 3
    16'b10111011_00110100 : OUT <= 3;  //187 / 52 = 3
    16'b10111011_00110101 : OUT <= 3;  //187 / 53 = 3
    16'b10111011_00110110 : OUT <= 3;  //187 / 54 = 3
    16'b10111011_00110111 : OUT <= 3;  //187 / 55 = 3
    16'b10111011_00111000 : OUT <= 3;  //187 / 56 = 3
    16'b10111011_00111001 : OUT <= 3;  //187 / 57 = 3
    16'b10111011_00111010 : OUT <= 3;  //187 / 58 = 3
    16'b10111011_00111011 : OUT <= 3;  //187 / 59 = 3
    16'b10111011_00111100 : OUT <= 3;  //187 / 60 = 3
    16'b10111011_00111101 : OUT <= 3;  //187 / 61 = 3
    16'b10111011_00111110 : OUT <= 3;  //187 / 62 = 3
    16'b10111011_00111111 : OUT <= 2;  //187 / 63 = 2
    16'b10111011_01000000 : OUT <= 2;  //187 / 64 = 2
    16'b10111011_01000001 : OUT <= 2;  //187 / 65 = 2
    16'b10111011_01000010 : OUT <= 2;  //187 / 66 = 2
    16'b10111011_01000011 : OUT <= 2;  //187 / 67 = 2
    16'b10111011_01000100 : OUT <= 2;  //187 / 68 = 2
    16'b10111011_01000101 : OUT <= 2;  //187 / 69 = 2
    16'b10111011_01000110 : OUT <= 2;  //187 / 70 = 2
    16'b10111011_01000111 : OUT <= 2;  //187 / 71 = 2
    16'b10111011_01001000 : OUT <= 2;  //187 / 72 = 2
    16'b10111011_01001001 : OUT <= 2;  //187 / 73 = 2
    16'b10111011_01001010 : OUT <= 2;  //187 / 74 = 2
    16'b10111011_01001011 : OUT <= 2;  //187 / 75 = 2
    16'b10111011_01001100 : OUT <= 2;  //187 / 76 = 2
    16'b10111011_01001101 : OUT <= 2;  //187 / 77 = 2
    16'b10111011_01001110 : OUT <= 2;  //187 / 78 = 2
    16'b10111011_01001111 : OUT <= 2;  //187 / 79 = 2
    16'b10111011_01010000 : OUT <= 2;  //187 / 80 = 2
    16'b10111011_01010001 : OUT <= 2;  //187 / 81 = 2
    16'b10111011_01010010 : OUT <= 2;  //187 / 82 = 2
    16'b10111011_01010011 : OUT <= 2;  //187 / 83 = 2
    16'b10111011_01010100 : OUT <= 2;  //187 / 84 = 2
    16'b10111011_01010101 : OUT <= 2;  //187 / 85 = 2
    16'b10111011_01010110 : OUT <= 2;  //187 / 86 = 2
    16'b10111011_01010111 : OUT <= 2;  //187 / 87 = 2
    16'b10111011_01011000 : OUT <= 2;  //187 / 88 = 2
    16'b10111011_01011001 : OUT <= 2;  //187 / 89 = 2
    16'b10111011_01011010 : OUT <= 2;  //187 / 90 = 2
    16'b10111011_01011011 : OUT <= 2;  //187 / 91 = 2
    16'b10111011_01011100 : OUT <= 2;  //187 / 92 = 2
    16'b10111011_01011101 : OUT <= 2;  //187 / 93 = 2
    16'b10111011_01011110 : OUT <= 1;  //187 / 94 = 1
    16'b10111011_01011111 : OUT <= 1;  //187 / 95 = 1
    16'b10111011_01100000 : OUT <= 1;  //187 / 96 = 1
    16'b10111011_01100001 : OUT <= 1;  //187 / 97 = 1
    16'b10111011_01100010 : OUT <= 1;  //187 / 98 = 1
    16'b10111011_01100011 : OUT <= 1;  //187 / 99 = 1
    16'b10111011_01100100 : OUT <= 1;  //187 / 100 = 1
    16'b10111011_01100101 : OUT <= 1;  //187 / 101 = 1
    16'b10111011_01100110 : OUT <= 1;  //187 / 102 = 1
    16'b10111011_01100111 : OUT <= 1;  //187 / 103 = 1
    16'b10111011_01101000 : OUT <= 1;  //187 / 104 = 1
    16'b10111011_01101001 : OUT <= 1;  //187 / 105 = 1
    16'b10111011_01101010 : OUT <= 1;  //187 / 106 = 1
    16'b10111011_01101011 : OUT <= 1;  //187 / 107 = 1
    16'b10111011_01101100 : OUT <= 1;  //187 / 108 = 1
    16'b10111011_01101101 : OUT <= 1;  //187 / 109 = 1
    16'b10111011_01101110 : OUT <= 1;  //187 / 110 = 1
    16'b10111011_01101111 : OUT <= 1;  //187 / 111 = 1
    16'b10111011_01110000 : OUT <= 1;  //187 / 112 = 1
    16'b10111011_01110001 : OUT <= 1;  //187 / 113 = 1
    16'b10111011_01110010 : OUT <= 1;  //187 / 114 = 1
    16'b10111011_01110011 : OUT <= 1;  //187 / 115 = 1
    16'b10111011_01110100 : OUT <= 1;  //187 / 116 = 1
    16'b10111011_01110101 : OUT <= 1;  //187 / 117 = 1
    16'b10111011_01110110 : OUT <= 1;  //187 / 118 = 1
    16'b10111011_01110111 : OUT <= 1;  //187 / 119 = 1
    16'b10111011_01111000 : OUT <= 1;  //187 / 120 = 1
    16'b10111011_01111001 : OUT <= 1;  //187 / 121 = 1
    16'b10111011_01111010 : OUT <= 1;  //187 / 122 = 1
    16'b10111011_01111011 : OUT <= 1;  //187 / 123 = 1
    16'b10111011_01111100 : OUT <= 1;  //187 / 124 = 1
    16'b10111011_01111101 : OUT <= 1;  //187 / 125 = 1
    16'b10111011_01111110 : OUT <= 1;  //187 / 126 = 1
    16'b10111011_01111111 : OUT <= 1;  //187 / 127 = 1
    16'b10111011_10000000 : OUT <= 1;  //187 / 128 = 1
    16'b10111011_10000001 : OUT <= 1;  //187 / 129 = 1
    16'b10111011_10000010 : OUT <= 1;  //187 / 130 = 1
    16'b10111011_10000011 : OUT <= 1;  //187 / 131 = 1
    16'b10111011_10000100 : OUT <= 1;  //187 / 132 = 1
    16'b10111011_10000101 : OUT <= 1;  //187 / 133 = 1
    16'b10111011_10000110 : OUT <= 1;  //187 / 134 = 1
    16'b10111011_10000111 : OUT <= 1;  //187 / 135 = 1
    16'b10111011_10001000 : OUT <= 1;  //187 / 136 = 1
    16'b10111011_10001001 : OUT <= 1;  //187 / 137 = 1
    16'b10111011_10001010 : OUT <= 1;  //187 / 138 = 1
    16'b10111011_10001011 : OUT <= 1;  //187 / 139 = 1
    16'b10111011_10001100 : OUT <= 1;  //187 / 140 = 1
    16'b10111011_10001101 : OUT <= 1;  //187 / 141 = 1
    16'b10111011_10001110 : OUT <= 1;  //187 / 142 = 1
    16'b10111011_10001111 : OUT <= 1;  //187 / 143 = 1
    16'b10111011_10010000 : OUT <= 1;  //187 / 144 = 1
    16'b10111011_10010001 : OUT <= 1;  //187 / 145 = 1
    16'b10111011_10010010 : OUT <= 1;  //187 / 146 = 1
    16'b10111011_10010011 : OUT <= 1;  //187 / 147 = 1
    16'b10111011_10010100 : OUT <= 1;  //187 / 148 = 1
    16'b10111011_10010101 : OUT <= 1;  //187 / 149 = 1
    16'b10111011_10010110 : OUT <= 1;  //187 / 150 = 1
    16'b10111011_10010111 : OUT <= 1;  //187 / 151 = 1
    16'b10111011_10011000 : OUT <= 1;  //187 / 152 = 1
    16'b10111011_10011001 : OUT <= 1;  //187 / 153 = 1
    16'b10111011_10011010 : OUT <= 1;  //187 / 154 = 1
    16'b10111011_10011011 : OUT <= 1;  //187 / 155 = 1
    16'b10111011_10011100 : OUT <= 1;  //187 / 156 = 1
    16'b10111011_10011101 : OUT <= 1;  //187 / 157 = 1
    16'b10111011_10011110 : OUT <= 1;  //187 / 158 = 1
    16'b10111011_10011111 : OUT <= 1;  //187 / 159 = 1
    16'b10111011_10100000 : OUT <= 1;  //187 / 160 = 1
    16'b10111011_10100001 : OUT <= 1;  //187 / 161 = 1
    16'b10111011_10100010 : OUT <= 1;  //187 / 162 = 1
    16'b10111011_10100011 : OUT <= 1;  //187 / 163 = 1
    16'b10111011_10100100 : OUT <= 1;  //187 / 164 = 1
    16'b10111011_10100101 : OUT <= 1;  //187 / 165 = 1
    16'b10111011_10100110 : OUT <= 1;  //187 / 166 = 1
    16'b10111011_10100111 : OUT <= 1;  //187 / 167 = 1
    16'b10111011_10101000 : OUT <= 1;  //187 / 168 = 1
    16'b10111011_10101001 : OUT <= 1;  //187 / 169 = 1
    16'b10111011_10101010 : OUT <= 1;  //187 / 170 = 1
    16'b10111011_10101011 : OUT <= 1;  //187 / 171 = 1
    16'b10111011_10101100 : OUT <= 1;  //187 / 172 = 1
    16'b10111011_10101101 : OUT <= 1;  //187 / 173 = 1
    16'b10111011_10101110 : OUT <= 1;  //187 / 174 = 1
    16'b10111011_10101111 : OUT <= 1;  //187 / 175 = 1
    16'b10111011_10110000 : OUT <= 1;  //187 / 176 = 1
    16'b10111011_10110001 : OUT <= 1;  //187 / 177 = 1
    16'b10111011_10110010 : OUT <= 1;  //187 / 178 = 1
    16'b10111011_10110011 : OUT <= 1;  //187 / 179 = 1
    16'b10111011_10110100 : OUT <= 1;  //187 / 180 = 1
    16'b10111011_10110101 : OUT <= 1;  //187 / 181 = 1
    16'b10111011_10110110 : OUT <= 1;  //187 / 182 = 1
    16'b10111011_10110111 : OUT <= 1;  //187 / 183 = 1
    16'b10111011_10111000 : OUT <= 1;  //187 / 184 = 1
    16'b10111011_10111001 : OUT <= 1;  //187 / 185 = 1
    16'b10111011_10111010 : OUT <= 1;  //187 / 186 = 1
    16'b10111011_10111011 : OUT <= 1;  //187 / 187 = 1
    16'b10111011_10111100 : OUT <= 0;  //187 / 188 = 0
    16'b10111011_10111101 : OUT <= 0;  //187 / 189 = 0
    16'b10111011_10111110 : OUT <= 0;  //187 / 190 = 0
    16'b10111011_10111111 : OUT <= 0;  //187 / 191 = 0
    16'b10111011_11000000 : OUT <= 0;  //187 / 192 = 0
    16'b10111011_11000001 : OUT <= 0;  //187 / 193 = 0
    16'b10111011_11000010 : OUT <= 0;  //187 / 194 = 0
    16'b10111011_11000011 : OUT <= 0;  //187 / 195 = 0
    16'b10111011_11000100 : OUT <= 0;  //187 / 196 = 0
    16'b10111011_11000101 : OUT <= 0;  //187 / 197 = 0
    16'b10111011_11000110 : OUT <= 0;  //187 / 198 = 0
    16'b10111011_11000111 : OUT <= 0;  //187 / 199 = 0
    16'b10111011_11001000 : OUT <= 0;  //187 / 200 = 0
    16'b10111011_11001001 : OUT <= 0;  //187 / 201 = 0
    16'b10111011_11001010 : OUT <= 0;  //187 / 202 = 0
    16'b10111011_11001011 : OUT <= 0;  //187 / 203 = 0
    16'b10111011_11001100 : OUT <= 0;  //187 / 204 = 0
    16'b10111011_11001101 : OUT <= 0;  //187 / 205 = 0
    16'b10111011_11001110 : OUT <= 0;  //187 / 206 = 0
    16'b10111011_11001111 : OUT <= 0;  //187 / 207 = 0
    16'b10111011_11010000 : OUT <= 0;  //187 / 208 = 0
    16'b10111011_11010001 : OUT <= 0;  //187 / 209 = 0
    16'b10111011_11010010 : OUT <= 0;  //187 / 210 = 0
    16'b10111011_11010011 : OUT <= 0;  //187 / 211 = 0
    16'b10111011_11010100 : OUT <= 0;  //187 / 212 = 0
    16'b10111011_11010101 : OUT <= 0;  //187 / 213 = 0
    16'b10111011_11010110 : OUT <= 0;  //187 / 214 = 0
    16'b10111011_11010111 : OUT <= 0;  //187 / 215 = 0
    16'b10111011_11011000 : OUT <= 0;  //187 / 216 = 0
    16'b10111011_11011001 : OUT <= 0;  //187 / 217 = 0
    16'b10111011_11011010 : OUT <= 0;  //187 / 218 = 0
    16'b10111011_11011011 : OUT <= 0;  //187 / 219 = 0
    16'b10111011_11011100 : OUT <= 0;  //187 / 220 = 0
    16'b10111011_11011101 : OUT <= 0;  //187 / 221 = 0
    16'b10111011_11011110 : OUT <= 0;  //187 / 222 = 0
    16'b10111011_11011111 : OUT <= 0;  //187 / 223 = 0
    16'b10111011_11100000 : OUT <= 0;  //187 / 224 = 0
    16'b10111011_11100001 : OUT <= 0;  //187 / 225 = 0
    16'b10111011_11100010 : OUT <= 0;  //187 / 226 = 0
    16'b10111011_11100011 : OUT <= 0;  //187 / 227 = 0
    16'b10111011_11100100 : OUT <= 0;  //187 / 228 = 0
    16'b10111011_11100101 : OUT <= 0;  //187 / 229 = 0
    16'b10111011_11100110 : OUT <= 0;  //187 / 230 = 0
    16'b10111011_11100111 : OUT <= 0;  //187 / 231 = 0
    16'b10111011_11101000 : OUT <= 0;  //187 / 232 = 0
    16'b10111011_11101001 : OUT <= 0;  //187 / 233 = 0
    16'b10111011_11101010 : OUT <= 0;  //187 / 234 = 0
    16'b10111011_11101011 : OUT <= 0;  //187 / 235 = 0
    16'b10111011_11101100 : OUT <= 0;  //187 / 236 = 0
    16'b10111011_11101101 : OUT <= 0;  //187 / 237 = 0
    16'b10111011_11101110 : OUT <= 0;  //187 / 238 = 0
    16'b10111011_11101111 : OUT <= 0;  //187 / 239 = 0
    16'b10111011_11110000 : OUT <= 0;  //187 / 240 = 0
    16'b10111011_11110001 : OUT <= 0;  //187 / 241 = 0
    16'b10111011_11110010 : OUT <= 0;  //187 / 242 = 0
    16'b10111011_11110011 : OUT <= 0;  //187 / 243 = 0
    16'b10111011_11110100 : OUT <= 0;  //187 / 244 = 0
    16'b10111011_11110101 : OUT <= 0;  //187 / 245 = 0
    16'b10111011_11110110 : OUT <= 0;  //187 / 246 = 0
    16'b10111011_11110111 : OUT <= 0;  //187 / 247 = 0
    16'b10111011_11111000 : OUT <= 0;  //187 / 248 = 0
    16'b10111011_11111001 : OUT <= 0;  //187 / 249 = 0
    16'b10111011_11111010 : OUT <= 0;  //187 / 250 = 0
    16'b10111011_11111011 : OUT <= 0;  //187 / 251 = 0
    16'b10111011_11111100 : OUT <= 0;  //187 / 252 = 0
    16'b10111011_11111101 : OUT <= 0;  //187 / 253 = 0
    16'b10111011_11111110 : OUT <= 0;  //187 / 254 = 0
    16'b10111011_11111111 : OUT <= 0;  //187 / 255 = 0
    16'b10111100_00000000 : OUT <= 0;  //188 / 0 = 0
    16'b10111100_00000001 : OUT <= 188;  //188 / 1 = 188
    16'b10111100_00000010 : OUT <= 94;  //188 / 2 = 94
    16'b10111100_00000011 : OUT <= 62;  //188 / 3 = 62
    16'b10111100_00000100 : OUT <= 47;  //188 / 4 = 47
    16'b10111100_00000101 : OUT <= 37;  //188 / 5 = 37
    16'b10111100_00000110 : OUT <= 31;  //188 / 6 = 31
    16'b10111100_00000111 : OUT <= 26;  //188 / 7 = 26
    16'b10111100_00001000 : OUT <= 23;  //188 / 8 = 23
    16'b10111100_00001001 : OUT <= 20;  //188 / 9 = 20
    16'b10111100_00001010 : OUT <= 18;  //188 / 10 = 18
    16'b10111100_00001011 : OUT <= 17;  //188 / 11 = 17
    16'b10111100_00001100 : OUT <= 15;  //188 / 12 = 15
    16'b10111100_00001101 : OUT <= 14;  //188 / 13 = 14
    16'b10111100_00001110 : OUT <= 13;  //188 / 14 = 13
    16'b10111100_00001111 : OUT <= 12;  //188 / 15 = 12
    16'b10111100_00010000 : OUT <= 11;  //188 / 16 = 11
    16'b10111100_00010001 : OUT <= 11;  //188 / 17 = 11
    16'b10111100_00010010 : OUT <= 10;  //188 / 18 = 10
    16'b10111100_00010011 : OUT <= 9;  //188 / 19 = 9
    16'b10111100_00010100 : OUT <= 9;  //188 / 20 = 9
    16'b10111100_00010101 : OUT <= 8;  //188 / 21 = 8
    16'b10111100_00010110 : OUT <= 8;  //188 / 22 = 8
    16'b10111100_00010111 : OUT <= 8;  //188 / 23 = 8
    16'b10111100_00011000 : OUT <= 7;  //188 / 24 = 7
    16'b10111100_00011001 : OUT <= 7;  //188 / 25 = 7
    16'b10111100_00011010 : OUT <= 7;  //188 / 26 = 7
    16'b10111100_00011011 : OUT <= 6;  //188 / 27 = 6
    16'b10111100_00011100 : OUT <= 6;  //188 / 28 = 6
    16'b10111100_00011101 : OUT <= 6;  //188 / 29 = 6
    16'b10111100_00011110 : OUT <= 6;  //188 / 30 = 6
    16'b10111100_00011111 : OUT <= 6;  //188 / 31 = 6
    16'b10111100_00100000 : OUT <= 5;  //188 / 32 = 5
    16'b10111100_00100001 : OUT <= 5;  //188 / 33 = 5
    16'b10111100_00100010 : OUT <= 5;  //188 / 34 = 5
    16'b10111100_00100011 : OUT <= 5;  //188 / 35 = 5
    16'b10111100_00100100 : OUT <= 5;  //188 / 36 = 5
    16'b10111100_00100101 : OUT <= 5;  //188 / 37 = 5
    16'b10111100_00100110 : OUT <= 4;  //188 / 38 = 4
    16'b10111100_00100111 : OUT <= 4;  //188 / 39 = 4
    16'b10111100_00101000 : OUT <= 4;  //188 / 40 = 4
    16'b10111100_00101001 : OUT <= 4;  //188 / 41 = 4
    16'b10111100_00101010 : OUT <= 4;  //188 / 42 = 4
    16'b10111100_00101011 : OUT <= 4;  //188 / 43 = 4
    16'b10111100_00101100 : OUT <= 4;  //188 / 44 = 4
    16'b10111100_00101101 : OUT <= 4;  //188 / 45 = 4
    16'b10111100_00101110 : OUT <= 4;  //188 / 46 = 4
    16'b10111100_00101111 : OUT <= 4;  //188 / 47 = 4
    16'b10111100_00110000 : OUT <= 3;  //188 / 48 = 3
    16'b10111100_00110001 : OUT <= 3;  //188 / 49 = 3
    16'b10111100_00110010 : OUT <= 3;  //188 / 50 = 3
    16'b10111100_00110011 : OUT <= 3;  //188 / 51 = 3
    16'b10111100_00110100 : OUT <= 3;  //188 / 52 = 3
    16'b10111100_00110101 : OUT <= 3;  //188 / 53 = 3
    16'b10111100_00110110 : OUT <= 3;  //188 / 54 = 3
    16'b10111100_00110111 : OUT <= 3;  //188 / 55 = 3
    16'b10111100_00111000 : OUT <= 3;  //188 / 56 = 3
    16'b10111100_00111001 : OUT <= 3;  //188 / 57 = 3
    16'b10111100_00111010 : OUT <= 3;  //188 / 58 = 3
    16'b10111100_00111011 : OUT <= 3;  //188 / 59 = 3
    16'b10111100_00111100 : OUT <= 3;  //188 / 60 = 3
    16'b10111100_00111101 : OUT <= 3;  //188 / 61 = 3
    16'b10111100_00111110 : OUT <= 3;  //188 / 62 = 3
    16'b10111100_00111111 : OUT <= 2;  //188 / 63 = 2
    16'b10111100_01000000 : OUT <= 2;  //188 / 64 = 2
    16'b10111100_01000001 : OUT <= 2;  //188 / 65 = 2
    16'b10111100_01000010 : OUT <= 2;  //188 / 66 = 2
    16'b10111100_01000011 : OUT <= 2;  //188 / 67 = 2
    16'b10111100_01000100 : OUT <= 2;  //188 / 68 = 2
    16'b10111100_01000101 : OUT <= 2;  //188 / 69 = 2
    16'b10111100_01000110 : OUT <= 2;  //188 / 70 = 2
    16'b10111100_01000111 : OUT <= 2;  //188 / 71 = 2
    16'b10111100_01001000 : OUT <= 2;  //188 / 72 = 2
    16'b10111100_01001001 : OUT <= 2;  //188 / 73 = 2
    16'b10111100_01001010 : OUT <= 2;  //188 / 74 = 2
    16'b10111100_01001011 : OUT <= 2;  //188 / 75 = 2
    16'b10111100_01001100 : OUT <= 2;  //188 / 76 = 2
    16'b10111100_01001101 : OUT <= 2;  //188 / 77 = 2
    16'b10111100_01001110 : OUT <= 2;  //188 / 78 = 2
    16'b10111100_01001111 : OUT <= 2;  //188 / 79 = 2
    16'b10111100_01010000 : OUT <= 2;  //188 / 80 = 2
    16'b10111100_01010001 : OUT <= 2;  //188 / 81 = 2
    16'b10111100_01010010 : OUT <= 2;  //188 / 82 = 2
    16'b10111100_01010011 : OUT <= 2;  //188 / 83 = 2
    16'b10111100_01010100 : OUT <= 2;  //188 / 84 = 2
    16'b10111100_01010101 : OUT <= 2;  //188 / 85 = 2
    16'b10111100_01010110 : OUT <= 2;  //188 / 86 = 2
    16'b10111100_01010111 : OUT <= 2;  //188 / 87 = 2
    16'b10111100_01011000 : OUT <= 2;  //188 / 88 = 2
    16'b10111100_01011001 : OUT <= 2;  //188 / 89 = 2
    16'b10111100_01011010 : OUT <= 2;  //188 / 90 = 2
    16'b10111100_01011011 : OUT <= 2;  //188 / 91 = 2
    16'b10111100_01011100 : OUT <= 2;  //188 / 92 = 2
    16'b10111100_01011101 : OUT <= 2;  //188 / 93 = 2
    16'b10111100_01011110 : OUT <= 2;  //188 / 94 = 2
    16'b10111100_01011111 : OUT <= 1;  //188 / 95 = 1
    16'b10111100_01100000 : OUT <= 1;  //188 / 96 = 1
    16'b10111100_01100001 : OUT <= 1;  //188 / 97 = 1
    16'b10111100_01100010 : OUT <= 1;  //188 / 98 = 1
    16'b10111100_01100011 : OUT <= 1;  //188 / 99 = 1
    16'b10111100_01100100 : OUT <= 1;  //188 / 100 = 1
    16'b10111100_01100101 : OUT <= 1;  //188 / 101 = 1
    16'b10111100_01100110 : OUT <= 1;  //188 / 102 = 1
    16'b10111100_01100111 : OUT <= 1;  //188 / 103 = 1
    16'b10111100_01101000 : OUT <= 1;  //188 / 104 = 1
    16'b10111100_01101001 : OUT <= 1;  //188 / 105 = 1
    16'b10111100_01101010 : OUT <= 1;  //188 / 106 = 1
    16'b10111100_01101011 : OUT <= 1;  //188 / 107 = 1
    16'b10111100_01101100 : OUT <= 1;  //188 / 108 = 1
    16'b10111100_01101101 : OUT <= 1;  //188 / 109 = 1
    16'b10111100_01101110 : OUT <= 1;  //188 / 110 = 1
    16'b10111100_01101111 : OUT <= 1;  //188 / 111 = 1
    16'b10111100_01110000 : OUT <= 1;  //188 / 112 = 1
    16'b10111100_01110001 : OUT <= 1;  //188 / 113 = 1
    16'b10111100_01110010 : OUT <= 1;  //188 / 114 = 1
    16'b10111100_01110011 : OUT <= 1;  //188 / 115 = 1
    16'b10111100_01110100 : OUT <= 1;  //188 / 116 = 1
    16'b10111100_01110101 : OUT <= 1;  //188 / 117 = 1
    16'b10111100_01110110 : OUT <= 1;  //188 / 118 = 1
    16'b10111100_01110111 : OUT <= 1;  //188 / 119 = 1
    16'b10111100_01111000 : OUT <= 1;  //188 / 120 = 1
    16'b10111100_01111001 : OUT <= 1;  //188 / 121 = 1
    16'b10111100_01111010 : OUT <= 1;  //188 / 122 = 1
    16'b10111100_01111011 : OUT <= 1;  //188 / 123 = 1
    16'b10111100_01111100 : OUT <= 1;  //188 / 124 = 1
    16'b10111100_01111101 : OUT <= 1;  //188 / 125 = 1
    16'b10111100_01111110 : OUT <= 1;  //188 / 126 = 1
    16'b10111100_01111111 : OUT <= 1;  //188 / 127 = 1
    16'b10111100_10000000 : OUT <= 1;  //188 / 128 = 1
    16'b10111100_10000001 : OUT <= 1;  //188 / 129 = 1
    16'b10111100_10000010 : OUT <= 1;  //188 / 130 = 1
    16'b10111100_10000011 : OUT <= 1;  //188 / 131 = 1
    16'b10111100_10000100 : OUT <= 1;  //188 / 132 = 1
    16'b10111100_10000101 : OUT <= 1;  //188 / 133 = 1
    16'b10111100_10000110 : OUT <= 1;  //188 / 134 = 1
    16'b10111100_10000111 : OUT <= 1;  //188 / 135 = 1
    16'b10111100_10001000 : OUT <= 1;  //188 / 136 = 1
    16'b10111100_10001001 : OUT <= 1;  //188 / 137 = 1
    16'b10111100_10001010 : OUT <= 1;  //188 / 138 = 1
    16'b10111100_10001011 : OUT <= 1;  //188 / 139 = 1
    16'b10111100_10001100 : OUT <= 1;  //188 / 140 = 1
    16'b10111100_10001101 : OUT <= 1;  //188 / 141 = 1
    16'b10111100_10001110 : OUT <= 1;  //188 / 142 = 1
    16'b10111100_10001111 : OUT <= 1;  //188 / 143 = 1
    16'b10111100_10010000 : OUT <= 1;  //188 / 144 = 1
    16'b10111100_10010001 : OUT <= 1;  //188 / 145 = 1
    16'b10111100_10010010 : OUT <= 1;  //188 / 146 = 1
    16'b10111100_10010011 : OUT <= 1;  //188 / 147 = 1
    16'b10111100_10010100 : OUT <= 1;  //188 / 148 = 1
    16'b10111100_10010101 : OUT <= 1;  //188 / 149 = 1
    16'b10111100_10010110 : OUT <= 1;  //188 / 150 = 1
    16'b10111100_10010111 : OUT <= 1;  //188 / 151 = 1
    16'b10111100_10011000 : OUT <= 1;  //188 / 152 = 1
    16'b10111100_10011001 : OUT <= 1;  //188 / 153 = 1
    16'b10111100_10011010 : OUT <= 1;  //188 / 154 = 1
    16'b10111100_10011011 : OUT <= 1;  //188 / 155 = 1
    16'b10111100_10011100 : OUT <= 1;  //188 / 156 = 1
    16'b10111100_10011101 : OUT <= 1;  //188 / 157 = 1
    16'b10111100_10011110 : OUT <= 1;  //188 / 158 = 1
    16'b10111100_10011111 : OUT <= 1;  //188 / 159 = 1
    16'b10111100_10100000 : OUT <= 1;  //188 / 160 = 1
    16'b10111100_10100001 : OUT <= 1;  //188 / 161 = 1
    16'b10111100_10100010 : OUT <= 1;  //188 / 162 = 1
    16'b10111100_10100011 : OUT <= 1;  //188 / 163 = 1
    16'b10111100_10100100 : OUT <= 1;  //188 / 164 = 1
    16'b10111100_10100101 : OUT <= 1;  //188 / 165 = 1
    16'b10111100_10100110 : OUT <= 1;  //188 / 166 = 1
    16'b10111100_10100111 : OUT <= 1;  //188 / 167 = 1
    16'b10111100_10101000 : OUT <= 1;  //188 / 168 = 1
    16'b10111100_10101001 : OUT <= 1;  //188 / 169 = 1
    16'b10111100_10101010 : OUT <= 1;  //188 / 170 = 1
    16'b10111100_10101011 : OUT <= 1;  //188 / 171 = 1
    16'b10111100_10101100 : OUT <= 1;  //188 / 172 = 1
    16'b10111100_10101101 : OUT <= 1;  //188 / 173 = 1
    16'b10111100_10101110 : OUT <= 1;  //188 / 174 = 1
    16'b10111100_10101111 : OUT <= 1;  //188 / 175 = 1
    16'b10111100_10110000 : OUT <= 1;  //188 / 176 = 1
    16'b10111100_10110001 : OUT <= 1;  //188 / 177 = 1
    16'b10111100_10110010 : OUT <= 1;  //188 / 178 = 1
    16'b10111100_10110011 : OUT <= 1;  //188 / 179 = 1
    16'b10111100_10110100 : OUT <= 1;  //188 / 180 = 1
    16'b10111100_10110101 : OUT <= 1;  //188 / 181 = 1
    16'b10111100_10110110 : OUT <= 1;  //188 / 182 = 1
    16'b10111100_10110111 : OUT <= 1;  //188 / 183 = 1
    16'b10111100_10111000 : OUT <= 1;  //188 / 184 = 1
    16'b10111100_10111001 : OUT <= 1;  //188 / 185 = 1
    16'b10111100_10111010 : OUT <= 1;  //188 / 186 = 1
    16'b10111100_10111011 : OUT <= 1;  //188 / 187 = 1
    16'b10111100_10111100 : OUT <= 1;  //188 / 188 = 1
    16'b10111100_10111101 : OUT <= 0;  //188 / 189 = 0
    16'b10111100_10111110 : OUT <= 0;  //188 / 190 = 0
    16'b10111100_10111111 : OUT <= 0;  //188 / 191 = 0
    16'b10111100_11000000 : OUT <= 0;  //188 / 192 = 0
    16'b10111100_11000001 : OUT <= 0;  //188 / 193 = 0
    16'b10111100_11000010 : OUT <= 0;  //188 / 194 = 0
    16'b10111100_11000011 : OUT <= 0;  //188 / 195 = 0
    16'b10111100_11000100 : OUT <= 0;  //188 / 196 = 0
    16'b10111100_11000101 : OUT <= 0;  //188 / 197 = 0
    16'b10111100_11000110 : OUT <= 0;  //188 / 198 = 0
    16'b10111100_11000111 : OUT <= 0;  //188 / 199 = 0
    16'b10111100_11001000 : OUT <= 0;  //188 / 200 = 0
    16'b10111100_11001001 : OUT <= 0;  //188 / 201 = 0
    16'b10111100_11001010 : OUT <= 0;  //188 / 202 = 0
    16'b10111100_11001011 : OUT <= 0;  //188 / 203 = 0
    16'b10111100_11001100 : OUT <= 0;  //188 / 204 = 0
    16'b10111100_11001101 : OUT <= 0;  //188 / 205 = 0
    16'b10111100_11001110 : OUT <= 0;  //188 / 206 = 0
    16'b10111100_11001111 : OUT <= 0;  //188 / 207 = 0
    16'b10111100_11010000 : OUT <= 0;  //188 / 208 = 0
    16'b10111100_11010001 : OUT <= 0;  //188 / 209 = 0
    16'b10111100_11010010 : OUT <= 0;  //188 / 210 = 0
    16'b10111100_11010011 : OUT <= 0;  //188 / 211 = 0
    16'b10111100_11010100 : OUT <= 0;  //188 / 212 = 0
    16'b10111100_11010101 : OUT <= 0;  //188 / 213 = 0
    16'b10111100_11010110 : OUT <= 0;  //188 / 214 = 0
    16'b10111100_11010111 : OUT <= 0;  //188 / 215 = 0
    16'b10111100_11011000 : OUT <= 0;  //188 / 216 = 0
    16'b10111100_11011001 : OUT <= 0;  //188 / 217 = 0
    16'b10111100_11011010 : OUT <= 0;  //188 / 218 = 0
    16'b10111100_11011011 : OUT <= 0;  //188 / 219 = 0
    16'b10111100_11011100 : OUT <= 0;  //188 / 220 = 0
    16'b10111100_11011101 : OUT <= 0;  //188 / 221 = 0
    16'b10111100_11011110 : OUT <= 0;  //188 / 222 = 0
    16'b10111100_11011111 : OUT <= 0;  //188 / 223 = 0
    16'b10111100_11100000 : OUT <= 0;  //188 / 224 = 0
    16'b10111100_11100001 : OUT <= 0;  //188 / 225 = 0
    16'b10111100_11100010 : OUT <= 0;  //188 / 226 = 0
    16'b10111100_11100011 : OUT <= 0;  //188 / 227 = 0
    16'b10111100_11100100 : OUT <= 0;  //188 / 228 = 0
    16'b10111100_11100101 : OUT <= 0;  //188 / 229 = 0
    16'b10111100_11100110 : OUT <= 0;  //188 / 230 = 0
    16'b10111100_11100111 : OUT <= 0;  //188 / 231 = 0
    16'b10111100_11101000 : OUT <= 0;  //188 / 232 = 0
    16'b10111100_11101001 : OUT <= 0;  //188 / 233 = 0
    16'b10111100_11101010 : OUT <= 0;  //188 / 234 = 0
    16'b10111100_11101011 : OUT <= 0;  //188 / 235 = 0
    16'b10111100_11101100 : OUT <= 0;  //188 / 236 = 0
    16'b10111100_11101101 : OUT <= 0;  //188 / 237 = 0
    16'b10111100_11101110 : OUT <= 0;  //188 / 238 = 0
    16'b10111100_11101111 : OUT <= 0;  //188 / 239 = 0
    16'b10111100_11110000 : OUT <= 0;  //188 / 240 = 0
    16'b10111100_11110001 : OUT <= 0;  //188 / 241 = 0
    16'b10111100_11110010 : OUT <= 0;  //188 / 242 = 0
    16'b10111100_11110011 : OUT <= 0;  //188 / 243 = 0
    16'b10111100_11110100 : OUT <= 0;  //188 / 244 = 0
    16'b10111100_11110101 : OUT <= 0;  //188 / 245 = 0
    16'b10111100_11110110 : OUT <= 0;  //188 / 246 = 0
    16'b10111100_11110111 : OUT <= 0;  //188 / 247 = 0
    16'b10111100_11111000 : OUT <= 0;  //188 / 248 = 0
    16'b10111100_11111001 : OUT <= 0;  //188 / 249 = 0
    16'b10111100_11111010 : OUT <= 0;  //188 / 250 = 0
    16'b10111100_11111011 : OUT <= 0;  //188 / 251 = 0
    16'b10111100_11111100 : OUT <= 0;  //188 / 252 = 0
    16'b10111100_11111101 : OUT <= 0;  //188 / 253 = 0
    16'b10111100_11111110 : OUT <= 0;  //188 / 254 = 0
    16'b10111100_11111111 : OUT <= 0;  //188 / 255 = 0
    16'b10111101_00000000 : OUT <= 0;  //189 / 0 = 0
    16'b10111101_00000001 : OUT <= 189;  //189 / 1 = 189
    16'b10111101_00000010 : OUT <= 94;  //189 / 2 = 94
    16'b10111101_00000011 : OUT <= 63;  //189 / 3 = 63
    16'b10111101_00000100 : OUT <= 47;  //189 / 4 = 47
    16'b10111101_00000101 : OUT <= 37;  //189 / 5 = 37
    16'b10111101_00000110 : OUT <= 31;  //189 / 6 = 31
    16'b10111101_00000111 : OUT <= 27;  //189 / 7 = 27
    16'b10111101_00001000 : OUT <= 23;  //189 / 8 = 23
    16'b10111101_00001001 : OUT <= 21;  //189 / 9 = 21
    16'b10111101_00001010 : OUT <= 18;  //189 / 10 = 18
    16'b10111101_00001011 : OUT <= 17;  //189 / 11 = 17
    16'b10111101_00001100 : OUT <= 15;  //189 / 12 = 15
    16'b10111101_00001101 : OUT <= 14;  //189 / 13 = 14
    16'b10111101_00001110 : OUT <= 13;  //189 / 14 = 13
    16'b10111101_00001111 : OUT <= 12;  //189 / 15 = 12
    16'b10111101_00010000 : OUT <= 11;  //189 / 16 = 11
    16'b10111101_00010001 : OUT <= 11;  //189 / 17 = 11
    16'b10111101_00010010 : OUT <= 10;  //189 / 18 = 10
    16'b10111101_00010011 : OUT <= 9;  //189 / 19 = 9
    16'b10111101_00010100 : OUT <= 9;  //189 / 20 = 9
    16'b10111101_00010101 : OUT <= 9;  //189 / 21 = 9
    16'b10111101_00010110 : OUT <= 8;  //189 / 22 = 8
    16'b10111101_00010111 : OUT <= 8;  //189 / 23 = 8
    16'b10111101_00011000 : OUT <= 7;  //189 / 24 = 7
    16'b10111101_00011001 : OUT <= 7;  //189 / 25 = 7
    16'b10111101_00011010 : OUT <= 7;  //189 / 26 = 7
    16'b10111101_00011011 : OUT <= 7;  //189 / 27 = 7
    16'b10111101_00011100 : OUT <= 6;  //189 / 28 = 6
    16'b10111101_00011101 : OUT <= 6;  //189 / 29 = 6
    16'b10111101_00011110 : OUT <= 6;  //189 / 30 = 6
    16'b10111101_00011111 : OUT <= 6;  //189 / 31 = 6
    16'b10111101_00100000 : OUT <= 5;  //189 / 32 = 5
    16'b10111101_00100001 : OUT <= 5;  //189 / 33 = 5
    16'b10111101_00100010 : OUT <= 5;  //189 / 34 = 5
    16'b10111101_00100011 : OUT <= 5;  //189 / 35 = 5
    16'b10111101_00100100 : OUT <= 5;  //189 / 36 = 5
    16'b10111101_00100101 : OUT <= 5;  //189 / 37 = 5
    16'b10111101_00100110 : OUT <= 4;  //189 / 38 = 4
    16'b10111101_00100111 : OUT <= 4;  //189 / 39 = 4
    16'b10111101_00101000 : OUT <= 4;  //189 / 40 = 4
    16'b10111101_00101001 : OUT <= 4;  //189 / 41 = 4
    16'b10111101_00101010 : OUT <= 4;  //189 / 42 = 4
    16'b10111101_00101011 : OUT <= 4;  //189 / 43 = 4
    16'b10111101_00101100 : OUT <= 4;  //189 / 44 = 4
    16'b10111101_00101101 : OUT <= 4;  //189 / 45 = 4
    16'b10111101_00101110 : OUT <= 4;  //189 / 46 = 4
    16'b10111101_00101111 : OUT <= 4;  //189 / 47 = 4
    16'b10111101_00110000 : OUT <= 3;  //189 / 48 = 3
    16'b10111101_00110001 : OUT <= 3;  //189 / 49 = 3
    16'b10111101_00110010 : OUT <= 3;  //189 / 50 = 3
    16'b10111101_00110011 : OUT <= 3;  //189 / 51 = 3
    16'b10111101_00110100 : OUT <= 3;  //189 / 52 = 3
    16'b10111101_00110101 : OUT <= 3;  //189 / 53 = 3
    16'b10111101_00110110 : OUT <= 3;  //189 / 54 = 3
    16'b10111101_00110111 : OUT <= 3;  //189 / 55 = 3
    16'b10111101_00111000 : OUT <= 3;  //189 / 56 = 3
    16'b10111101_00111001 : OUT <= 3;  //189 / 57 = 3
    16'b10111101_00111010 : OUT <= 3;  //189 / 58 = 3
    16'b10111101_00111011 : OUT <= 3;  //189 / 59 = 3
    16'b10111101_00111100 : OUT <= 3;  //189 / 60 = 3
    16'b10111101_00111101 : OUT <= 3;  //189 / 61 = 3
    16'b10111101_00111110 : OUT <= 3;  //189 / 62 = 3
    16'b10111101_00111111 : OUT <= 3;  //189 / 63 = 3
    16'b10111101_01000000 : OUT <= 2;  //189 / 64 = 2
    16'b10111101_01000001 : OUT <= 2;  //189 / 65 = 2
    16'b10111101_01000010 : OUT <= 2;  //189 / 66 = 2
    16'b10111101_01000011 : OUT <= 2;  //189 / 67 = 2
    16'b10111101_01000100 : OUT <= 2;  //189 / 68 = 2
    16'b10111101_01000101 : OUT <= 2;  //189 / 69 = 2
    16'b10111101_01000110 : OUT <= 2;  //189 / 70 = 2
    16'b10111101_01000111 : OUT <= 2;  //189 / 71 = 2
    16'b10111101_01001000 : OUT <= 2;  //189 / 72 = 2
    16'b10111101_01001001 : OUT <= 2;  //189 / 73 = 2
    16'b10111101_01001010 : OUT <= 2;  //189 / 74 = 2
    16'b10111101_01001011 : OUT <= 2;  //189 / 75 = 2
    16'b10111101_01001100 : OUT <= 2;  //189 / 76 = 2
    16'b10111101_01001101 : OUT <= 2;  //189 / 77 = 2
    16'b10111101_01001110 : OUT <= 2;  //189 / 78 = 2
    16'b10111101_01001111 : OUT <= 2;  //189 / 79 = 2
    16'b10111101_01010000 : OUT <= 2;  //189 / 80 = 2
    16'b10111101_01010001 : OUT <= 2;  //189 / 81 = 2
    16'b10111101_01010010 : OUT <= 2;  //189 / 82 = 2
    16'b10111101_01010011 : OUT <= 2;  //189 / 83 = 2
    16'b10111101_01010100 : OUT <= 2;  //189 / 84 = 2
    16'b10111101_01010101 : OUT <= 2;  //189 / 85 = 2
    16'b10111101_01010110 : OUT <= 2;  //189 / 86 = 2
    16'b10111101_01010111 : OUT <= 2;  //189 / 87 = 2
    16'b10111101_01011000 : OUT <= 2;  //189 / 88 = 2
    16'b10111101_01011001 : OUT <= 2;  //189 / 89 = 2
    16'b10111101_01011010 : OUT <= 2;  //189 / 90 = 2
    16'b10111101_01011011 : OUT <= 2;  //189 / 91 = 2
    16'b10111101_01011100 : OUT <= 2;  //189 / 92 = 2
    16'b10111101_01011101 : OUT <= 2;  //189 / 93 = 2
    16'b10111101_01011110 : OUT <= 2;  //189 / 94 = 2
    16'b10111101_01011111 : OUT <= 1;  //189 / 95 = 1
    16'b10111101_01100000 : OUT <= 1;  //189 / 96 = 1
    16'b10111101_01100001 : OUT <= 1;  //189 / 97 = 1
    16'b10111101_01100010 : OUT <= 1;  //189 / 98 = 1
    16'b10111101_01100011 : OUT <= 1;  //189 / 99 = 1
    16'b10111101_01100100 : OUT <= 1;  //189 / 100 = 1
    16'b10111101_01100101 : OUT <= 1;  //189 / 101 = 1
    16'b10111101_01100110 : OUT <= 1;  //189 / 102 = 1
    16'b10111101_01100111 : OUT <= 1;  //189 / 103 = 1
    16'b10111101_01101000 : OUT <= 1;  //189 / 104 = 1
    16'b10111101_01101001 : OUT <= 1;  //189 / 105 = 1
    16'b10111101_01101010 : OUT <= 1;  //189 / 106 = 1
    16'b10111101_01101011 : OUT <= 1;  //189 / 107 = 1
    16'b10111101_01101100 : OUT <= 1;  //189 / 108 = 1
    16'b10111101_01101101 : OUT <= 1;  //189 / 109 = 1
    16'b10111101_01101110 : OUT <= 1;  //189 / 110 = 1
    16'b10111101_01101111 : OUT <= 1;  //189 / 111 = 1
    16'b10111101_01110000 : OUT <= 1;  //189 / 112 = 1
    16'b10111101_01110001 : OUT <= 1;  //189 / 113 = 1
    16'b10111101_01110010 : OUT <= 1;  //189 / 114 = 1
    16'b10111101_01110011 : OUT <= 1;  //189 / 115 = 1
    16'b10111101_01110100 : OUT <= 1;  //189 / 116 = 1
    16'b10111101_01110101 : OUT <= 1;  //189 / 117 = 1
    16'b10111101_01110110 : OUT <= 1;  //189 / 118 = 1
    16'b10111101_01110111 : OUT <= 1;  //189 / 119 = 1
    16'b10111101_01111000 : OUT <= 1;  //189 / 120 = 1
    16'b10111101_01111001 : OUT <= 1;  //189 / 121 = 1
    16'b10111101_01111010 : OUT <= 1;  //189 / 122 = 1
    16'b10111101_01111011 : OUT <= 1;  //189 / 123 = 1
    16'b10111101_01111100 : OUT <= 1;  //189 / 124 = 1
    16'b10111101_01111101 : OUT <= 1;  //189 / 125 = 1
    16'b10111101_01111110 : OUT <= 1;  //189 / 126 = 1
    16'b10111101_01111111 : OUT <= 1;  //189 / 127 = 1
    16'b10111101_10000000 : OUT <= 1;  //189 / 128 = 1
    16'b10111101_10000001 : OUT <= 1;  //189 / 129 = 1
    16'b10111101_10000010 : OUT <= 1;  //189 / 130 = 1
    16'b10111101_10000011 : OUT <= 1;  //189 / 131 = 1
    16'b10111101_10000100 : OUT <= 1;  //189 / 132 = 1
    16'b10111101_10000101 : OUT <= 1;  //189 / 133 = 1
    16'b10111101_10000110 : OUT <= 1;  //189 / 134 = 1
    16'b10111101_10000111 : OUT <= 1;  //189 / 135 = 1
    16'b10111101_10001000 : OUT <= 1;  //189 / 136 = 1
    16'b10111101_10001001 : OUT <= 1;  //189 / 137 = 1
    16'b10111101_10001010 : OUT <= 1;  //189 / 138 = 1
    16'b10111101_10001011 : OUT <= 1;  //189 / 139 = 1
    16'b10111101_10001100 : OUT <= 1;  //189 / 140 = 1
    16'b10111101_10001101 : OUT <= 1;  //189 / 141 = 1
    16'b10111101_10001110 : OUT <= 1;  //189 / 142 = 1
    16'b10111101_10001111 : OUT <= 1;  //189 / 143 = 1
    16'b10111101_10010000 : OUT <= 1;  //189 / 144 = 1
    16'b10111101_10010001 : OUT <= 1;  //189 / 145 = 1
    16'b10111101_10010010 : OUT <= 1;  //189 / 146 = 1
    16'b10111101_10010011 : OUT <= 1;  //189 / 147 = 1
    16'b10111101_10010100 : OUT <= 1;  //189 / 148 = 1
    16'b10111101_10010101 : OUT <= 1;  //189 / 149 = 1
    16'b10111101_10010110 : OUT <= 1;  //189 / 150 = 1
    16'b10111101_10010111 : OUT <= 1;  //189 / 151 = 1
    16'b10111101_10011000 : OUT <= 1;  //189 / 152 = 1
    16'b10111101_10011001 : OUT <= 1;  //189 / 153 = 1
    16'b10111101_10011010 : OUT <= 1;  //189 / 154 = 1
    16'b10111101_10011011 : OUT <= 1;  //189 / 155 = 1
    16'b10111101_10011100 : OUT <= 1;  //189 / 156 = 1
    16'b10111101_10011101 : OUT <= 1;  //189 / 157 = 1
    16'b10111101_10011110 : OUT <= 1;  //189 / 158 = 1
    16'b10111101_10011111 : OUT <= 1;  //189 / 159 = 1
    16'b10111101_10100000 : OUT <= 1;  //189 / 160 = 1
    16'b10111101_10100001 : OUT <= 1;  //189 / 161 = 1
    16'b10111101_10100010 : OUT <= 1;  //189 / 162 = 1
    16'b10111101_10100011 : OUT <= 1;  //189 / 163 = 1
    16'b10111101_10100100 : OUT <= 1;  //189 / 164 = 1
    16'b10111101_10100101 : OUT <= 1;  //189 / 165 = 1
    16'b10111101_10100110 : OUT <= 1;  //189 / 166 = 1
    16'b10111101_10100111 : OUT <= 1;  //189 / 167 = 1
    16'b10111101_10101000 : OUT <= 1;  //189 / 168 = 1
    16'b10111101_10101001 : OUT <= 1;  //189 / 169 = 1
    16'b10111101_10101010 : OUT <= 1;  //189 / 170 = 1
    16'b10111101_10101011 : OUT <= 1;  //189 / 171 = 1
    16'b10111101_10101100 : OUT <= 1;  //189 / 172 = 1
    16'b10111101_10101101 : OUT <= 1;  //189 / 173 = 1
    16'b10111101_10101110 : OUT <= 1;  //189 / 174 = 1
    16'b10111101_10101111 : OUT <= 1;  //189 / 175 = 1
    16'b10111101_10110000 : OUT <= 1;  //189 / 176 = 1
    16'b10111101_10110001 : OUT <= 1;  //189 / 177 = 1
    16'b10111101_10110010 : OUT <= 1;  //189 / 178 = 1
    16'b10111101_10110011 : OUT <= 1;  //189 / 179 = 1
    16'b10111101_10110100 : OUT <= 1;  //189 / 180 = 1
    16'b10111101_10110101 : OUT <= 1;  //189 / 181 = 1
    16'b10111101_10110110 : OUT <= 1;  //189 / 182 = 1
    16'b10111101_10110111 : OUT <= 1;  //189 / 183 = 1
    16'b10111101_10111000 : OUT <= 1;  //189 / 184 = 1
    16'b10111101_10111001 : OUT <= 1;  //189 / 185 = 1
    16'b10111101_10111010 : OUT <= 1;  //189 / 186 = 1
    16'b10111101_10111011 : OUT <= 1;  //189 / 187 = 1
    16'b10111101_10111100 : OUT <= 1;  //189 / 188 = 1
    16'b10111101_10111101 : OUT <= 1;  //189 / 189 = 1
    16'b10111101_10111110 : OUT <= 0;  //189 / 190 = 0
    16'b10111101_10111111 : OUT <= 0;  //189 / 191 = 0
    16'b10111101_11000000 : OUT <= 0;  //189 / 192 = 0
    16'b10111101_11000001 : OUT <= 0;  //189 / 193 = 0
    16'b10111101_11000010 : OUT <= 0;  //189 / 194 = 0
    16'b10111101_11000011 : OUT <= 0;  //189 / 195 = 0
    16'b10111101_11000100 : OUT <= 0;  //189 / 196 = 0
    16'b10111101_11000101 : OUT <= 0;  //189 / 197 = 0
    16'b10111101_11000110 : OUT <= 0;  //189 / 198 = 0
    16'b10111101_11000111 : OUT <= 0;  //189 / 199 = 0
    16'b10111101_11001000 : OUT <= 0;  //189 / 200 = 0
    16'b10111101_11001001 : OUT <= 0;  //189 / 201 = 0
    16'b10111101_11001010 : OUT <= 0;  //189 / 202 = 0
    16'b10111101_11001011 : OUT <= 0;  //189 / 203 = 0
    16'b10111101_11001100 : OUT <= 0;  //189 / 204 = 0
    16'b10111101_11001101 : OUT <= 0;  //189 / 205 = 0
    16'b10111101_11001110 : OUT <= 0;  //189 / 206 = 0
    16'b10111101_11001111 : OUT <= 0;  //189 / 207 = 0
    16'b10111101_11010000 : OUT <= 0;  //189 / 208 = 0
    16'b10111101_11010001 : OUT <= 0;  //189 / 209 = 0
    16'b10111101_11010010 : OUT <= 0;  //189 / 210 = 0
    16'b10111101_11010011 : OUT <= 0;  //189 / 211 = 0
    16'b10111101_11010100 : OUT <= 0;  //189 / 212 = 0
    16'b10111101_11010101 : OUT <= 0;  //189 / 213 = 0
    16'b10111101_11010110 : OUT <= 0;  //189 / 214 = 0
    16'b10111101_11010111 : OUT <= 0;  //189 / 215 = 0
    16'b10111101_11011000 : OUT <= 0;  //189 / 216 = 0
    16'b10111101_11011001 : OUT <= 0;  //189 / 217 = 0
    16'b10111101_11011010 : OUT <= 0;  //189 / 218 = 0
    16'b10111101_11011011 : OUT <= 0;  //189 / 219 = 0
    16'b10111101_11011100 : OUT <= 0;  //189 / 220 = 0
    16'b10111101_11011101 : OUT <= 0;  //189 / 221 = 0
    16'b10111101_11011110 : OUT <= 0;  //189 / 222 = 0
    16'b10111101_11011111 : OUT <= 0;  //189 / 223 = 0
    16'b10111101_11100000 : OUT <= 0;  //189 / 224 = 0
    16'b10111101_11100001 : OUT <= 0;  //189 / 225 = 0
    16'b10111101_11100010 : OUT <= 0;  //189 / 226 = 0
    16'b10111101_11100011 : OUT <= 0;  //189 / 227 = 0
    16'b10111101_11100100 : OUT <= 0;  //189 / 228 = 0
    16'b10111101_11100101 : OUT <= 0;  //189 / 229 = 0
    16'b10111101_11100110 : OUT <= 0;  //189 / 230 = 0
    16'b10111101_11100111 : OUT <= 0;  //189 / 231 = 0
    16'b10111101_11101000 : OUT <= 0;  //189 / 232 = 0
    16'b10111101_11101001 : OUT <= 0;  //189 / 233 = 0
    16'b10111101_11101010 : OUT <= 0;  //189 / 234 = 0
    16'b10111101_11101011 : OUT <= 0;  //189 / 235 = 0
    16'b10111101_11101100 : OUT <= 0;  //189 / 236 = 0
    16'b10111101_11101101 : OUT <= 0;  //189 / 237 = 0
    16'b10111101_11101110 : OUT <= 0;  //189 / 238 = 0
    16'b10111101_11101111 : OUT <= 0;  //189 / 239 = 0
    16'b10111101_11110000 : OUT <= 0;  //189 / 240 = 0
    16'b10111101_11110001 : OUT <= 0;  //189 / 241 = 0
    16'b10111101_11110010 : OUT <= 0;  //189 / 242 = 0
    16'b10111101_11110011 : OUT <= 0;  //189 / 243 = 0
    16'b10111101_11110100 : OUT <= 0;  //189 / 244 = 0
    16'b10111101_11110101 : OUT <= 0;  //189 / 245 = 0
    16'b10111101_11110110 : OUT <= 0;  //189 / 246 = 0
    16'b10111101_11110111 : OUT <= 0;  //189 / 247 = 0
    16'b10111101_11111000 : OUT <= 0;  //189 / 248 = 0
    16'b10111101_11111001 : OUT <= 0;  //189 / 249 = 0
    16'b10111101_11111010 : OUT <= 0;  //189 / 250 = 0
    16'b10111101_11111011 : OUT <= 0;  //189 / 251 = 0
    16'b10111101_11111100 : OUT <= 0;  //189 / 252 = 0
    16'b10111101_11111101 : OUT <= 0;  //189 / 253 = 0
    16'b10111101_11111110 : OUT <= 0;  //189 / 254 = 0
    16'b10111101_11111111 : OUT <= 0;  //189 / 255 = 0
    16'b10111110_00000000 : OUT <= 0;  //190 / 0 = 0
    16'b10111110_00000001 : OUT <= 190;  //190 / 1 = 190
    16'b10111110_00000010 : OUT <= 95;  //190 / 2 = 95
    16'b10111110_00000011 : OUT <= 63;  //190 / 3 = 63
    16'b10111110_00000100 : OUT <= 47;  //190 / 4 = 47
    16'b10111110_00000101 : OUT <= 38;  //190 / 5 = 38
    16'b10111110_00000110 : OUT <= 31;  //190 / 6 = 31
    16'b10111110_00000111 : OUT <= 27;  //190 / 7 = 27
    16'b10111110_00001000 : OUT <= 23;  //190 / 8 = 23
    16'b10111110_00001001 : OUT <= 21;  //190 / 9 = 21
    16'b10111110_00001010 : OUT <= 19;  //190 / 10 = 19
    16'b10111110_00001011 : OUT <= 17;  //190 / 11 = 17
    16'b10111110_00001100 : OUT <= 15;  //190 / 12 = 15
    16'b10111110_00001101 : OUT <= 14;  //190 / 13 = 14
    16'b10111110_00001110 : OUT <= 13;  //190 / 14 = 13
    16'b10111110_00001111 : OUT <= 12;  //190 / 15 = 12
    16'b10111110_00010000 : OUT <= 11;  //190 / 16 = 11
    16'b10111110_00010001 : OUT <= 11;  //190 / 17 = 11
    16'b10111110_00010010 : OUT <= 10;  //190 / 18 = 10
    16'b10111110_00010011 : OUT <= 10;  //190 / 19 = 10
    16'b10111110_00010100 : OUT <= 9;  //190 / 20 = 9
    16'b10111110_00010101 : OUT <= 9;  //190 / 21 = 9
    16'b10111110_00010110 : OUT <= 8;  //190 / 22 = 8
    16'b10111110_00010111 : OUT <= 8;  //190 / 23 = 8
    16'b10111110_00011000 : OUT <= 7;  //190 / 24 = 7
    16'b10111110_00011001 : OUT <= 7;  //190 / 25 = 7
    16'b10111110_00011010 : OUT <= 7;  //190 / 26 = 7
    16'b10111110_00011011 : OUT <= 7;  //190 / 27 = 7
    16'b10111110_00011100 : OUT <= 6;  //190 / 28 = 6
    16'b10111110_00011101 : OUT <= 6;  //190 / 29 = 6
    16'b10111110_00011110 : OUT <= 6;  //190 / 30 = 6
    16'b10111110_00011111 : OUT <= 6;  //190 / 31 = 6
    16'b10111110_00100000 : OUT <= 5;  //190 / 32 = 5
    16'b10111110_00100001 : OUT <= 5;  //190 / 33 = 5
    16'b10111110_00100010 : OUT <= 5;  //190 / 34 = 5
    16'b10111110_00100011 : OUT <= 5;  //190 / 35 = 5
    16'b10111110_00100100 : OUT <= 5;  //190 / 36 = 5
    16'b10111110_00100101 : OUT <= 5;  //190 / 37 = 5
    16'b10111110_00100110 : OUT <= 5;  //190 / 38 = 5
    16'b10111110_00100111 : OUT <= 4;  //190 / 39 = 4
    16'b10111110_00101000 : OUT <= 4;  //190 / 40 = 4
    16'b10111110_00101001 : OUT <= 4;  //190 / 41 = 4
    16'b10111110_00101010 : OUT <= 4;  //190 / 42 = 4
    16'b10111110_00101011 : OUT <= 4;  //190 / 43 = 4
    16'b10111110_00101100 : OUT <= 4;  //190 / 44 = 4
    16'b10111110_00101101 : OUT <= 4;  //190 / 45 = 4
    16'b10111110_00101110 : OUT <= 4;  //190 / 46 = 4
    16'b10111110_00101111 : OUT <= 4;  //190 / 47 = 4
    16'b10111110_00110000 : OUT <= 3;  //190 / 48 = 3
    16'b10111110_00110001 : OUT <= 3;  //190 / 49 = 3
    16'b10111110_00110010 : OUT <= 3;  //190 / 50 = 3
    16'b10111110_00110011 : OUT <= 3;  //190 / 51 = 3
    16'b10111110_00110100 : OUT <= 3;  //190 / 52 = 3
    16'b10111110_00110101 : OUT <= 3;  //190 / 53 = 3
    16'b10111110_00110110 : OUT <= 3;  //190 / 54 = 3
    16'b10111110_00110111 : OUT <= 3;  //190 / 55 = 3
    16'b10111110_00111000 : OUT <= 3;  //190 / 56 = 3
    16'b10111110_00111001 : OUT <= 3;  //190 / 57 = 3
    16'b10111110_00111010 : OUT <= 3;  //190 / 58 = 3
    16'b10111110_00111011 : OUT <= 3;  //190 / 59 = 3
    16'b10111110_00111100 : OUT <= 3;  //190 / 60 = 3
    16'b10111110_00111101 : OUT <= 3;  //190 / 61 = 3
    16'b10111110_00111110 : OUT <= 3;  //190 / 62 = 3
    16'b10111110_00111111 : OUT <= 3;  //190 / 63 = 3
    16'b10111110_01000000 : OUT <= 2;  //190 / 64 = 2
    16'b10111110_01000001 : OUT <= 2;  //190 / 65 = 2
    16'b10111110_01000010 : OUT <= 2;  //190 / 66 = 2
    16'b10111110_01000011 : OUT <= 2;  //190 / 67 = 2
    16'b10111110_01000100 : OUT <= 2;  //190 / 68 = 2
    16'b10111110_01000101 : OUT <= 2;  //190 / 69 = 2
    16'b10111110_01000110 : OUT <= 2;  //190 / 70 = 2
    16'b10111110_01000111 : OUT <= 2;  //190 / 71 = 2
    16'b10111110_01001000 : OUT <= 2;  //190 / 72 = 2
    16'b10111110_01001001 : OUT <= 2;  //190 / 73 = 2
    16'b10111110_01001010 : OUT <= 2;  //190 / 74 = 2
    16'b10111110_01001011 : OUT <= 2;  //190 / 75 = 2
    16'b10111110_01001100 : OUT <= 2;  //190 / 76 = 2
    16'b10111110_01001101 : OUT <= 2;  //190 / 77 = 2
    16'b10111110_01001110 : OUT <= 2;  //190 / 78 = 2
    16'b10111110_01001111 : OUT <= 2;  //190 / 79 = 2
    16'b10111110_01010000 : OUT <= 2;  //190 / 80 = 2
    16'b10111110_01010001 : OUT <= 2;  //190 / 81 = 2
    16'b10111110_01010010 : OUT <= 2;  //190 / 82 = 2
    16'b10111110_01010011 : OUT <= 2;  //190 / 83 = 2
    16'b10111110_01010100 : OUT <= 2;  //190 / 84 = 2
    16'b10111110_01010101 : OUT <= 2;  //190 / 85 = 2
    16'b10111110_01010110 : OUT <= 2;  //190 / 86 = 2
    16'b10111110_01010111 : OUT <= 2;  //190 / 87 = 2
    16'b10111110_01011000 : OUT <= 2;  //190 / 88 = 2
    16'b10111110_01011001 : OUT <= 2;  //190 / 89 = 2
    16'b10111110_01011010 : OUT <= 2;  //190 / 90 = 2
    16'b10111110_01011011 : OUT <= 2;  //190 / 91 = 2
    16'b10111110_01011100 : OUT <= 2;  //190 / 92 = 2
    16'b10111110_01011101 : OUT <= 2;  //190 / 93 = 2
    16'b10111110_01011110 : OUT <= 2;  //190 / 94 = 2
    16'b10111110_01011111 : OUT <= 2;  //190 / 95 = 2
    16'b10111110_01100000 : OUT <= 1;  //190 / 96 = 1
    16'b10111110_01100001 : OUT <= 1;  //190 / 97 = 1
    16'b10111110_01100010 : OUT <= 1;  //190 / 98 = 1
    16'b10111110_01100011 : OUT <= 1;  //190 / 99 = 1
    16'b10111110_01100100 : OUT <= 1;  //190 / 100 = 1
    16'b10111110_01100101 : OUT <= 1;  //190 / 101 = 1
    16'b10111110_01100110 : OUT <= 1;  //190 / 102 = 1
    16'b10111110_01100111 : OUT <= 1;  //190 / 103 = 1
    16'b10111110_01101000 : OUT <= 1;  //190 / 104 = 1
    16'b10111110_01101001 : OUT <= 1;  //190 / 105 = 1
    16'b10111110_01101010 : OUT <= 1;  //190 / 106 = 1
    16'b10111110_01101011 : OUT <= 1;  //190 / 107 = 1
    16'b10111110_01101100 : OUT <= 1;  //190 / 108 = 1
    16'b10111110_01101101 : OUT <= 1;  //190 / 109 = 1
    16'b10111110_01101110 : OUT <= 1;  //190 / 110 = 1
    16'b10111110_01101111 : OUT <= 1;  //190 / 111 = 1
    16'b10111110_01110000 : OUT <= 1;  //190 / 112 = 1
    16'b10111110_01110001 : OUT <= 1;  //190 / 113 = 1
    16'b10111110_01110010 : OUT <= 1;  //190 / 114 = 1
    16'b10111110_01110011 : OUT <= 1;  //190 / 115 = 1
    16'b10111110_01110100 : OUT <= 1;  //190 / 116 = 1
    16'b10111110_01110101 : OUT <= 1;  //190 / 117 = 1
    16'b10111110_01110110 : OUT <= 1;  //190 / 118 = 1
    16'b10111110_01110111 : OUT <= 1;  //190 / 119 = 1
    16'b10111110_01111000 : OUT <= 1;  //190 / 120 = 1
    16'b10111110_01111001 : OUT <= 1;  //190 / 121 = 1
    16'b10111110_01111010 : OUT <= 1;  //190 / 122 = 1
    16'b10111110_01111011 : OUT <= 1;  //190 / 123 = 1
    16'b10111110_01111100 : OUT <= 1;  //190 / 124 = 1
    16'b10111110_01111101 : OUT <= 1;  //190 / 125 = 1
    16'b10111110_01111110 : OUT <= 1;  //190 / 126 = 1
    16'b10111110_01111111 : OUT <= 1;  //190 / 127 = 1
    16'b10111110_10000000 : OUT <= 1;  //190 / 128 = 1
    16'b10111110_10000001 : OUT <= 1;  //190 / 129 = 1
    16'b10111110_10000010 : OUT <= 1;  //190 / 130 = 1
    16'b10111110_10000011 : OUT <= 1;  //190 / 131 = 1
    16'b10111110_10000100 : OUT <= 1;  //190 / 132 = 1
    16'b10111110_10000101 : OUT <= 1;  //190 / 133 = 1
    16'b10111110_10000110 : OUT <= 1;  //190 / 134 = 1
    16'b10111110_10000111 : OUT <= 1;  //190 / 135 = 1
    16'b10111110_10001000 : OUT <= 1;  //190 / 136 = 1
    16'b10111110_10001001 : OUT <= 1;  //190 / 137 = 1
    16'b10111110_10001010 : OUT <= 1;  //190 / 138 = 1
    16'b10111110_10001011 : OUT <= 1;  //190 / 139 = 1
    16'b10111110_10001100 : OUT <= 1;  //190 / 140 = 1
    16'b10111110_10001101 : OUT <= 1;  //190 / 141 = 1
    16'b10111110_10001110 : OUT <= 1;  //190 / 142 = 1
    16'b10111110_10001111 : OUT <= 1;  //190 / 143 = 1
    16'b10111110_10010000 : OUT <= 1;  //190 / 144 = 1
    16'b10111110_10010001 : OUT <= 1;  //190 / 145 = 1
    16'b10111110_10010010 : OUT <= 1;  //190 / 146 = 1
    16'b10111110_10010011 : OUT <= 1;  //190 / 147 = 1
    16'b10111110_10010100 : OUT <= 1;  //190 / 148 = 1
    16'b10111110_10010101 : OUT <= 1;  //190 / 149 = 1
    16'b10111110_10010110 : OUT <= 1;  //190 / 150 = 1
    16'b10111110_10010111 : OUT <= 1;  //190 / 151 = 1
    16'b10111110_10011000 : OUT <= 1;  //190 / 152 = 1
    16'b10111110_10011001 : OUT <= 1;  //190 / 153 = 1
    16'b10111110_10011010 : OUT <= 1;  //190 / 154 = 1
    16'b10111110_10011011 : OUT <= 1;  //190 / 155 = 1
    16'b10111110_10011100 : OUT <= 1;  //190 / 156 = 1
    16'b10111110_10011101 : OUT <= 1;  //190 / 157 = 1
    16'b10111110_10011110 : OUT <= 1;  //190 / 158 = 1
    16'b10111110_10011111 : OUT <= 1;  //190 / 159 = 1
    16'b10111110_10100000 : OUT <= 1;  //190 / 160 = 1
    16'b10111110_10100001 : OUT <= 1;  //190 / 161 = 1
    16'b10111110_10100010 : OUT <= 1;  //190 / 162 = 1
    16'b10111110_10100011 : OUT <= 1;  //190 / 163 = 1
    16'b10111110_10100100 : OUT <= 1;  //190 / 164 = 1
    16'b10111110_10100101 : OUT <= 1;  //190 / 165 = 1
    16'b10111110_10100110 : OUT <= 1;  //190 / 166 = 1
    16'b10111110_10100111 : OUT <= 1;  //190 / 167 = 1
    16'b10111110_10101000 : OUT <= 1;  //190 / 168 = 1
    16'b10111110_10101001 : OUT <= 1;  //190 / 169 = 1
    16'b10111110_10101010 : OUT <= 1;  //190 / 170 = 1
    16'b10111110_10101011 : OUT <= 1;  //190 / 171 = 1
    16'b10111110_10101100 : OUT <= 1;  //190 / 172 = 1
    16'b10111110_10101101 : OUT <= 1;  //190 / 173 = 1
    16'b10111110_10101110 : OUT <= 1;  //190 / 174 = 1
    16'b10111110_10101111 : OUT <= 1;  //190 / 175 = 1
    16'b10111110_10110000 : OUT <= 1;  //190 / 176 = 1
    16'b10111110_10110001 : OUT <= 1;  //190 / 177 = 1
    16'b10111110_10110010 : OUT <= 1;  //190 / 178 = 1
    16'b10111110_10110011 : OUT <= 1;  //190 / 179 = 1
    16'b10111110_10110100 : OUT <= 1;  //190 / 180 = 1
    16'b10111110_10110101 : OUT <= 1;  //190 / 181 = 1
    16'b10111110_10110110 : OUT <= 1;  //190 / 182 = 1
    16'b10111110_10110111 : OUT <= 1;  //190 / 183 = 1
    16'b10111110_10111000 : OUT <= 1;  //190 / 184 = 1
    16'b10111110_10111001 : OUT <= 1;  //190 / 185 = 1
    16'b10111110_10111010 : OUT <= 1;  //190 / 186 = 1
    16'b10111110_10111011 : OUT <= 1;  //190 / 187 = 1
    16'b10111110_10111100 : OUT <= 1;  //190 / 188 = 1
    16'b10111110_10111101 : OUT <= 1;  //190 / 189 = 1
    16'b10111110_10111110 : OUT <= 1;  //190 / 190 = 1
    16'b10111110_10111111 : OUT <= 0;  //190 / 191 = 0
    16'b10111110_11000000 : OUT <= 0;  //190 / 192 = 0
    16'b10111110_11000001 : OUT <= 0;  //190 / 193 = 0
    16'b10111110_11000010 : OUT <= 0;  //190 / 194 = 0
    16'b10111110_11000011 : OUT <= 0;  //190 / 195 = 0
    16'b10111110_11000100 : OUT <= 0;  //190 / 196 = 0
    16'b10111110_11000101 : OUT <= 0;  //190 / 197 = 0
    16'b10111110_11000110 : OUT <= 0;  //190 / 198 = 0
    16'b10111110_11000111 : OUT <= 0;  //190 / 199 = 0
    16'b10111110_11001000 : OUT <= 0;  //190 / 200 = 0
    16'b10111110_11001001 : OUT <= 0;  //190 / 201 = 0
    16'b10111110_11001010 : OUT <= 0;  //190 / 202 = 0
    16'b10111110_11001011 : OUT <= 0;  //190 / 203 = 0
    16'b10111110_11001100 : OUT <= 0;  //190 / 204 = 0
    16'b10111110_11001101 : OUT <= 0;  //190 / 205 = 0
    16'b10111110_11001110 : OUT <= 0;  //190 / 206 = 0
    16'b10111110_11001111 : OUT <= 0;  //190 / 207 = 0
    16'b10111110_11010000 : OUT <= 0;  //190 / 208 = 0
    16'b10111110_11010001 : OUT <= 0;  //190 / 209 = 0
    16'b10111110_11010010 : OUT <= 0;  //190 / 210 = 0
    16'b10111110_11010011 : OUT <= 0;  //190 / 211 = 0
    16'b10111110_11010100 : OUT <= 0;  //190 / 212 = 0
    16'b10111110_11010101 : OUT <= 0;  //190 / 213 = 0
    16'b10111110_11010110 : OUT <= 0;  //190 / 214 = 0
    16'b10111110_11010111 : OUT <= 0;  //190 / 215 = 0
    16'b10111110_11011000 : OUT <= 0;  //190 / 216 = 0
    16'b10111110_11011001 : OUT <= 0;  //190 / 217 = 0
    16'b10111110_11011010 : OUT <= 0;  //190 / 218 = 0
    16'b10111110_11011011 : OUT <= 0;  //190 / 219 = 0
    16'b10111110_11011100 : OUT <= 0;  //190 / 220 = 0
    16'b10111110_11011101 : OUT <= 0;  //190 / 221 = 0
    16'b10111110_11011110 : OUT <= 0;  //190 / 222 = 0
    16'b10111110_11011111 : OUT <= 0;  //190 / 223 = 0
    16'b10111110_11100000 : OUT <= 0;  //190 / 224 = 0
    16'b10111110_11100001 : OUT <= 0;  //190 / 225 = 0
    16'b10111110_11100010 : OUT <= 0;  //190 / 226 = 0
    16'b10111110_11100011 : OUT <= 0;  //190 / 227 = 0
    16'b10111110_11100100 : OUT <= 0;  //190 / 228 = 0
    16'b10111110_11100101 : OUT <= 0;  //190 / 229 = 0
    16'b10111110_11100110 : OUT <= 0;  //190 / 230 = 0
    16'b10111110_11100111 : OUT <= 0;  //190 / 231 = 0
    16'b10111110_11101000 : OUT <= 0;  //190 / 232 = 0
    16'b10111110_11101001 : OUT <= 0;  //190 / 233 = 0
    16'b10111110_11101010 : OUT <= 0;  //190 / 234 = 0
    16'b10111110_11101011 : OUT <= 0;  //190 / 235 = 0
    16'b10111110_11101100 : OUT <= 0;  //190 / 236 = 0
    16'b10111110_11101101 : OUT <= 0;  //190 / 237 = 0
    16'b10111110_11101110 : OUT <= 0;  //190 / 238 = 0
    16'b10111110_11101111 : OUT <= 0;  //190 / 239 = 0
    16'b10111110_11110000 : OUT <= 0;  //190 / 240 = 0
    16'b10111110_11110001 : OUT <= 0;  //190 / 241 = 0
    16'b10111110_11110010 : OUT <= 0;  //190 / 242 = 0
    16'b10111110_11110011 : OUT <= 0;  //190 / 243 = 0
    16'b10111110_11110100 : OUT <= 0;  //190 / 244 = 0
    16'b10111110_11110101 : OUT <= 0;  //190 / 245 = 0
    16'b10111110_11110110 : OUT <= 0;  //190 / 246 = 0
    16'b10111110_11110111 : OUT <= 0;  //190 / 247 = 0
    16'b10111110_11111000 : OUT <= 0;  //190 / 248 = 0
    16'b10111110_11111001 : OUT <= 0;  //190 / 249 = 0
    16'b10111110_11111010 : OUT <= 0;  //190 / 250 = 0
    16'b10111110_11111011 : OUT <= 0;  //190 / 251 = 0
    16'b10111110_11111100 : OUT <= 0;  //190 / 252 = 0
    16'b10111110_11111101 : OUT <= 0;  //190 / 253 = 0
    16'b10111110_11111110 : OUT <= 0;  //190 / 254 = 0
    16'b10111110_11111111 : OUT <= 0;  //190 / 255 = 0
    16'b10111111_00000000 : OUT <= 0;  //191 / 0 = 0
    16'b10111111_00000001 : OUT <= 191;  //191 / 1 = 191
    16'b10111111_00000010 : OUT <= 95;  //191 / 2 = 95
    16'b10111111_00000011 : OUT <= 63;  //191 / 3 = 63
    16'b10111111_00000100 : OUT <= 47;  //191 / 4 = 47
    16'b10111111_00000101 : OUT <= 38;  //191 / 5 = 38
    16'b10111111_00000110 : OUT <= 31;  //191 / 6 = 31
    16'b10111111_00000111 : OUT <= 27;  //191 / 7 = 27
    16'b10111111_00001000 : OUT <= 23;  //191 / 8 = 23
    16'b10111111_00001001 : OUT <= 21;  //191 / 9 = 21
    16'b10111111_00001010 : OUT <= 19;  //191 / 10 = 19
    16'b10111111_00001011 : OUT <= 17;  //191 / 11 = 17
    16'b10111111_00001100 : OUT <= 15;  //191 / 12 = 15
    16'b10111111_00001101 : OUT <= 14;  //191 / 13 = 14
    16'b10111111_00001110 : OUT <= 13;  //191 / 14 = 13
    16'b10111111_00001111 : OUT <= 12;  //191 / 15 = 12
    16'b10111111_00010000 : OUT <= 11;  //191 / 16 = 11
    16'b10111111_00010001 : OUT <= 11;  //191 / 17 = 11
    16'b10111111_00010010 : OUT <= 10;  //191 / 18 = 10
    16'b10111111_00010011 : OUT <= 10;  //191 / 19 = 10
    16'b10111111_00010100 : OUT <= 9;  //191 / 20 = 9
    16'b10111111_00010101 : OUT <= 9;  //191 / 21 = 9
    16'b10111111_00010110 : OUT <= 8;  //191 / 22 = 8
    16'b10111111_00010111 : OUT <= 8;  //191 / 23 = 8
    16'b10111111_00011000 : OUT <= 7;  //191 / 24 = 7
    16'b10111111_00011001 : OUT <= 7;  //191 / 25 = 7
    16'b10111111_00011010 : OUT <= 7;  //191 / 26 = 7
    16'b10111111_00011011 : OUT <= 7;  //191 / 27 = 7
    16'b10111111_00011100 : OUT <= 6;  //191 / 28 = 6
    16'b10111111_00011101 : OUT <= 6;  //191 / 29 = 6
    16'b10111111_00011110 : OUT <= 6;  //191 / 30 = 6
    16'b10111111_00011111 : OUT <= 6;  //191 / 31 = 6
    16'b10111111_00100000 : OUT <= 5;  //191 / 32 = 5
    16'b10111111_00100001 : OUT <= 5;  //191 / 33 = 5
    16'b10111111_00100010 : OUT <= 5;  //191 / 34 = 5
    16'b10111111_00100011 : OUT <= 5;  //191 / 35 = 5
    16'b10111111_00100100 : OUT <= 5;  //191 / 36 = 5
    16'b10111111_00100101 : OUT <= 5;  //191 / 37 = 5
    16'b10111111_00100110 : OUT <= 5;  //191 / 38 = 5
    16'b10111111_00100111 : OUT <= 4;  //191 / 39 = 4
    16'b10111111_00101000 : OUT <= 4;  //191 / 40 = 4
    16'b10111111_00101001 : OUT <= 4;  //191 / 41 = 4
    16'b10111111_00101010 : OUT <= 4;  //191 / 42 = 4
    16'b10111111_00101011 : OUT <= 4;  //191 / 43 = 4
    16'b10111111_00101100 : OUT <= 4;  //191 / 44 = 4
    16'b10111111_00101101 : OUT <= 4;  //191 / 45 = 4
    16'b10111111_00101110 : OUT <= 4;  //191 / 46 = 4
    16'b10111111_00101111 : OUT <= 4;  //191 / 47 = 4
    16'b10111111_00110000 : OUT <= 3;  //191 / 48 = 3
    16'b10111111_00110001 : OUT <= 3;  //191 / 49 = 3
    16'b10111111_00110010 : OUT <= 3;  //191 / 50 = 3
    16'b10111111_00110011 : OUT <= 3;  //191 / 51 = 3
    16'b10111111_00110100 : OUT <= 3;  //191 / 52 = 3
    16'b10111111_00110101 : OUT <= 3;  //191 / 53 = 3
    16'b10111111_00110110 : OUT <= 3;  //191 / 54 = 3
    16'b10111111_00110111 : OUT <= 3;  //191 / 55 = 3
    16'b10111111_00111000 : OUT <= 3;  //191 / 56 = 3
    16'b10111111_00111001 : OUT <= 3;  //191 / 57 = 3
    16'b10111111_00111010 : OUT <= 3;  //191 / 58 = 3
    16'b10111111_00111011 : OUT <= 3;  //191 / 59 = 3
    16'b10111111_00111100 : OUT <= 3;  //191 / 60 = 3
    16'b10111111_00111101 : OUT <= 3;  //191 / 61 = 3
    16'b10111111_00111110 : OUT <= 3;  //191 / 62 = 3
    16'b10111111_00111111 : OUT <= 3;  //191 / 63 = 3
    16'b10111111_01000000 : OUT <= 2;  //191 / 64 = 2
    16'b10111111_01000001 : OUT <= 2;  //191 / 65 = 2
    16'b10111111_01000010 : OUT <= 2;  //191 / 66 = 2
    16'b10111111_01000011 : OUT <= 2;  //191 / 67 = 2
    16'b10111111_01000100 : OUT <= 2;  //191 / 68 = 2
    16'b10111111_01000101 : OUT <= 2;  //191 / 69 = 2
    16'b10111111_01000110 : OUT <= 2;  //191 / 70 = 2
    16'b10111111_01000111 : OUT <= 2;  //191 / 71 = 2
    16'b10111111_01001000 : OUT <= 2;  //191 / 72 = 2
    16'b10111111_01001001 : OUT <= 2;  //191 / 73 = 2
    16'b10111111_01001010 : OUT <= 2;  //191 / 74 = 2
    16'b10111111_01001011 : OUT <= 2;  //191 / 75 = 2
    16'b10111111_01001100 : OUT <= 2;  //191 / 76 = 2
    16'b10111111_01001101 : OUT <= 2;  //191 / 77 = 2
    16'b10111111_01001110 : OUT <= 2;  //191 / 78 = 2
    16'b10111111_01001111 : OUT <= 2;  //191 / 79 = 2
    16'b10111111_01010000 : OUT <= 2;  //191 / 80 = 2
    16'b10111111_01010001 : OUT <= 2;  //191 / 81 = 2
    16'b10111111_01010010 : OUT <= 2;  //191 / 82 = 2
    16'b10111111_01010011 : OUT <= 2;  //191 / 83 = 2
    16'b10111111_01010100 : OUT <= 2;  //191 / 84 = 2
    16'b10111111_01010101 : OUT <= 2;  //191 / 85 = 2
    16'b10111111_01010110 : OUT <= 2;  //191 / 86 = 2
    16'b10111111_01010111 : OUT <= 2;  //191 / 87 = 2
    16'b10111111_01011000 : OUT <= 2;  //191 / 88 = 2
    16'b10111111_01011001 : OUT <= 2;  //191 / 89 = 2
    16'b10111111_01011010 : OUT <= 2;  //191 / 90 = 2
    16'b10111111_01011011 : OUT <= 2;  //191 / 91 = 2
    16'b10111111_01011100 : OUT <= 2;  //191 / 92 = 2
    16'b10111111_01011101 : OUT <= 2;  //191 / 93 = 2
    16'b10111111_01011110 : OUT <= 2;  //191 / 94 = 2
    16'b10111111_01011111 : OUT <= 2;  //191 / 95 = 2
    16'b10111111_01100000 : OUT <= 1;  //191 / 96 = 1
    16'b10111111_01100001 : OUT <= 1;  //191 / 97 = 1
    16'b10111111_01100010 : OUT <= 1;  //191 / 98 = 1
    16'b10111111_01100011 : OUT <= 1;  //191 / 99 = 1
    16'b10111111_01100100 : OUT <= 1;  //191 / 100 = 1
    16'b10111111_01100101 : OUT <= 1;  //191 / 101 = 1
    16'b10111111_01100110 : OUT <= 1;  //191 / 102 = 1
    16'b10111111_01100111 : OUT <= 1;  //191 / 103 = 1
    16'b10111111_01101000 : OUT <= 1;  //191 / 104 = 1
    16'b10111111_01101001 : OUT <= 1;  //191 / 105 = 1
    16'b10111111_01101010 : OUT <= 1;  //191 / 106 = 1
    16'b10111111_01101011 : OUT <= 1;  //191 / 107 = 1
    16'b10111111_01101100 : OUT <= 1;  //191 / 108 = 1
    16'b10111111_01101101 : OUT <= 1;  //191 / 109 = 1
    16'b10111111_01101110 : OUT <= 1;  //191 / 110 = 1
    16'b10111111_01101111 : OUT <= 1;  //191 / 111 = 1
    16'b10111111_01110000 : OUT <= 1;  //191 / 112 = 1
    16'b10111111_01110001 : OUT <= 1;  //191 / 113 = 1
    16'b10111111_01110010 : OUT <= 1;  //191 / 114 = 1
    16'b10111111_01110011 : OUT <= 1;  //191 / 115 = 1
    16'b10111111_01110100 : OUT <= 1;  //191 / 116 = 1
    16'b10111111_01110101 : OUT <= 1;  //191 / 117 = 1
    16'b10111111_01110110 : OUT <= 1;  //191 / 118 = 1
    16'b10111111_01110111 : OUT <= 1;  //191 / 119 = 1
    16'b10111111_01111000 : OUT <= 1;  //191 / 120 = 1
    16'b10111111_01111001 : OUT <= 1;  //191 / 121 = 1
    16'b10111111_01111010 : OUT <= 1;  //191 / 122 = 1
    16'b10111111_01111011 : OUT <= 1;  //191 / 123 = 1
    16'b10111111_01111100 : OUT <= 1;  //191 / 124 = 1
    16'b10111111_01111101 : OUT <= 1;  //191 / 125 = 1
    16'b10111111_01111110 : OUT <= 1;  //191 / 126 = 1
    16'b10111111_01111111 : OUT <= 1;  //191 / 127 = 1
    16'b10111111_10000000 : OUT <= 1;  //191 / 128 = 1
    16'b10111111_10000001 : OUT <= 1;  //191 / 129 = 1
    16'b10111111_10000010 : OUT <= 1;  //191 / 130 = 1
    16'b10111111_10000011 : OUT <= 1;  //191 / 131 = 1
    16'b10111111_10000100 : OUT <= 1;  //191 / 132 = 1
    16'b10111111_10000101 : OUT <= 1;  //191 / 133 = 1
    16'b10111111_10000110 : OUT <= 1;  //191 / 134 = 1
    16'b10111111_10000111 : OUT <= 1;  //191 / 135 = 1
    16'b10111111_10001000 : OUT <= 1;  //191 / 136 = 1
    16'b10111111_10001001 : OUT <= 1;  //191 / 137 = 1
    16'b10111111_10001010 : OUT <= 1;  //191 / 138 = 1
    16'b10111111_10001011 : OUT <= 1;  //191 / 139 = 1
    16'b10111111_10001100 : OUT <= 1;  //191 / 140 = 1
    16'b10111111_10001101 : OUT <= 1;  //191 / 141 = 1
    16'b10111111_10001110 : OUT <= 1;  //191 / 142 = 1
    16'b10111111_10001111 : OUT <= 1;  //191 / 143 = 1
    16'b10111111_10010000 : OUT <= 1;  //191 / 144 = 1
    16'b10111111_10010001 : OUT <= 1;  //191 / 145 = 1
    16'b10111111_10010010 : OUT <= 1;  //191 / 146 = 1
    16'b10111111_10010011 : OUT <= 1;  //191 / 147 = 1
    16'b10111111_10010100 : OUT <= 1;  //191 / 148 = 1
    16'b10111111_10010101 : OUT <= 1;  //191 / 149 = 1
    16'b10111111_10010110 : OUT <= 1;  //191 / 150 = 1
    16'b10111111_10010111 : OUT <= 1;  //191 / 151 = 1
    16'b10111111_10011000 : OUT <= 1;  //191 / 152 = 1
    16'b10111111_10011001 : OUT <= 1;  //191 / 153 = 1
    16'b10111111_10011010 : OUT <= 1;  //191 / 154 = 1
    16'b10111111_10011011 : OUT <= 1;  //191 / 155 = 1
    16'b10111111_10011100 : OUT <= 1;  //191 / 156 = 1
    16'b10111111_10011101 : OUT <= 1;  //191 / 157 = 1
    16'b10111111_10011110 : OUT <= 1;  //191 / 158 = 1
    16'b10111111_10011111 : OUT <= 1;  //191 / 159 = 1
    16'b10111111_10100000 : OUT <= 1;  //191 / 160 = 1
    16'b10111111_10100001 : OUT <= 1;  //191 / 161 = 1
    16'b10111111_10100010 : OUT <= 1;  //191 / 162 = 1
    16'b10111111_10100011 : OUT <= 1;  //191 / 163 = 1
    16'b10111111_10100100 : OUT <= 1;  //191 / 164 = 1
    16'b10111111_10100101 : OUT <= 1;  //191 / 165 = 1
    16'b10111111_10100110 : OUT <= 1;  //191 / 166 = 1
    16'b10111111_10100111 : OUT <= 1;  //191 / 167 = 1
    16'b10111111_10101000 : OUT <= 1;  //191 / 168 = 1
    16'b10111111_10101001 : OUT <= 1;  //191 / 169 = 1
    16'b10111111_10101010 : OUT <= 1;  //191 / 170 = 1
    16'b10111111_10101011 : OUT <= 1;  //191 / 171 = 1
    16'b10111111_10101100 : OUT <= 1;  //191 / 172 = 1
    16'b10111111_10101101 : OUT <= 1;  //191 / 173 = 1
    16'b10111111_10101110 : OUT <= 1;  //191 / 174 = 1
    16'b10111111_10101111 : OUT <= 1;  //191 / 175 = 1
    16'b10111111_10110000 : OUT <= 1;  //191 / 176 = 1
    16'b10111111_10110001 : OUT <= 1;  //191 / 177 = 1
    16'b10111111_10110010 : OUT <= 1;  //191 / 178 = 1
    16'b10111111_10110011 : OUT <= 1;  //191 / 179 = 1
    16'b10111111_10110100 : OUT <= 1;  //191 / 180 = 1
    16'b10111111_10110101 : OUT <= 1;  //191 / 181 = 1
    16'b10111111_10110110 : OUT <= 1;  //191 / 182 = 1
    16'b10111111_10110111 : OUT <= 1;  //191 / 183 = 1
    16'b10111111_10111000 : OUT <= 1;  //191 / 184 = 1
    16'b10111111_10111001 : OUT <= 1;  //191 / 185 = 1
    16'b10111111_10111010 : OUT <= 1;  //191 / 186 = 1
    16'b10111111_10111011 : OUT <= 1;  //191 / 187 = 1
    16'b10111111_10111100 : OUT <= 1;  //191 / 188 = 1
    16'b10111111_10111101 : OUT <= 1;  //191 / 189 = 1
    16'b10111111_10111110 : OUT <= 1;  //191 / 190 = 1
    16'b10111111_10111111 : OUT <= 1;  //191 / 191 = 1
    16'b10111111_11000000 : OUT <= 0;  //191 / 192 = 0
    16'b10111111_11000001 : OUT <= 0;  //191 / 193 = 0
    16'b10111111_11000010 : OUT <= 0;  //191 / 194 = 0
    16'b10111111_11000011 : OUT <= 0;  //191 / 195 = 0
    16'b10111111_11000100 : OUT <= 0;  //191 / 196 = 0
    16'b10111111_11000101 : OUT <= 0;  //191 / 197 = 0
    16'b10111111_11000110 : OUT <= 0;  //191 / 198 = 0
    16'b10111111_11000111 : OUT <= 0;  //191 / 199 = 0
    16'b10111111_11001000 : OUT <= 0;  //191 / 200 = 0
    16'b10111111_11001001 : OUT <= 0;  //191 / 201 = 0
    16'b10111111_11001010 : OUT <= 0;  //191 / 202 = 0
    16'b10111111_11001011 : OUT <= 0;  //191 / 203 = 0
    16'b10111111_11001100 : OUT <= 0;  //191 / 204 = 0
    16'b10111111_11001101 : OUT <= 0;  //191 / 205 = 0
    16'b10111111_11001110 : OUT <= 0;  //191 / 206 = 0
    16'b10111111_11001111 : OUT <= 0;  //191 / 207 = 0
    16'b10111111_11010000 : OUT <= 0;  //191 / 208 = 0
    16'b10111111_11010001 : OUT <= 0;  //191 / 209 = 0
    16'b10111111_11010010 : OUT <= 0;  //191 / 210 = 0
    16'b10111111_11010011 : OUT <= 0;  //191 / 211 = 0
    16'b10111111_11010100 : OUT <= 0;  //191 / 212 = 0
    16'b10111111_11010101 : OUT <= 0;  //191 / 213 = 0
    16'b10111111_11010110 : OUT <= 0;  //191 / 214 = 0
    16'b10111111_11010111 : OUT <= 0;  //191 / 215 = 0
    16'b10111111_11011000 : OUT <= 0;  //191 / 216 = 0
    16'b10111111_11011001 : OUT <= 0;  //191 / 217 = 0
    16'b10111111_11011010 : OUT <= 0;  //191 / 218 = 0
    16'b10111111_11011011 : OUT <= 0;  //191 / 219 = 0
    16'b10111111_11011100 : OUT <= 0;  //191 / 220 = 0
    16'b10111111_11011101 : OUT <= 0;  //191 / 221 = 0
    16'b10111111_11011110 : OUT <= 0;  //191 / 222 = 0
    16'b10111111_11011111 : OUT <= 0;  //191 / 223 = 0
    16'b10111111_11100000 : OUT <= 0;  //191 / 224 = 0
    16'b10111111_11100001 : OUT <= 0;  //191 / 225 = 0
    16'b10111111_11100010 : OUT <= 0;  //191 / 226 = 0
    16'b10111111_11100011 : OUT <= 0;  //191 / 227 = 0
    16'b10111111_11100100 : OUT <= 0;  //191 / 228 = 0
    16'b10111111_11100101 : OUT <= 0;  //191 / 229 = 0
    16'b10111111_11100110 : OUT <= 0;  //191 / 230 = 0
    16'b10111111_11100111 : OUT <= 0;  //191 / 231 = 0
    16'b10111111_11101000 : OUT <= 0;  //191 / 232 = 0
    16'b10111111_11101001 : OUT <= 0;  //191 / 233 = 0
    16'b10111111_11101010 : OUT <= 0;  //191 / 234 = 0
    16'b10111111_11101011 : OUT <= 0;  //191 / 235 = 0
    16'b10111111_11101100 : OUT <= 0;  //191 / 236 = 0
    16'b10111111_11101101 : OUT <= 0;  //191 / 237 = 0
    16'b10111111_11101110 : OUT <= 0;  //191 / 238 = 0
    16'b10111111_11101111 : OUT <= 0;  //191 / 239 = 0
    16'b10111111_11110000 : OUT <= 0;  //191 / 240 = 0
    16'b10111111_11110001 : OUT <= 0;  //191 / 241 = 0
    16'b10111111_11110010 : OUT <= 0;  //191 / 242 = 0
    16'b10111111_11110011 : OUT <= 0;  //191 / 243 = 0
    16'b10111111_11110100 : OUT <= 0;  //191 / 244 = 0
    16'b10111111_11110101 : OUT <= 0;  //191 / 245 = 0
    16'b10111111_11110110 : OUT <= 0;  //191 / 246 = 0
    16'b10111111_11110111 : OUT <= 0;  //191 / 247 = 0
    16'b10111111_11111000 : OUT <= 0;  //191 / 248 = 0
    16'b10111111_11111001 : OUT <= 0;  //191 / 249 = 0
    16'b10111111_11111010 : OUT <= 0;  //191 / 250 = 0
    16'b10111111_11111011 : OUT <= 0;  //191 / 251 = 0
    16'b10111111_11111100 : OUT <= 0;  //191 / 252 = 0
    16'b10111111_11111101 : OUT <= 0;  //191 / 253 = 0
    16'b10111111_11111110 : OUT <= 0;  //191 / 254 = 0
    16'b10111111_11111111 : OUT <= 0;  //191 / 255 = 0
    16'b11000000_00000000 : OUT <= 0;  //192 / 0 = 0
    16'b11000000_00000001 : OUT <= 192;  //192 / 1 = 192
    16'b11000000_00000010 : OUT <= 96;  //192 / 2 = 96
    16'b11000000_00000011 : OUT <= 64;  //192 / 3 = 64
    16'b11000000_00000100 : OUT <= 48;  //192 / 4 = 48
    16'b11000000_00000101 : OUT <= 38;  //192 / 5 = 38
    16'b11000000_00000110 : OUT <= 32;  //192 / 6 = 32
    16'b11000000_00000111 : OUT <= 27;  //192 / 7 = 27
    16'b11000000_00001000 : OUT <= 24;  //192 / 8 = 24
    16'b11000000_00001001 : OUT <= 21;  //192 / 9 = 21
    16'b11000000_00001010 : OUT <= 19;  //192 / 10 = 19
    16'b11000000_00001011 : OUT <= 17;  //192 / 11 = 17
    16'b11000000_00001100 : OUT <= 16;  //192 / 12 = 16
    16'b11000000_00001101 : OUT <= 14;  //192 / 13 = 14
    16'b11000000_00001110 : OUT <= 13;  //192 / 14 = 13
    16'b11000000_00001111 : OUT <= 12;  //192 / 15 = 12
    16'b11000000_00010000 : OUT <= 12;  //192 / 16 = 12
    16'b11000000_00010001 : OUT <= 11;  //192 / 17 = 11
    16'b11000000_00010010 : OUT <= 10;  //192 / 18 = 10
    16'b11000000_00010011 : OUT <= 10;  //192 / 19 = 10
    16'b11000000_00010100 : OUT <= 9;  //192 / 20 = 9
    16'b11000000_00010101 : OUT <= 9;  //192 / 21 = 9
    16'b11000000_00010110 : OUT <= 8;  //192 / 22 = 8
    16'b11000000_00010111 : OUT <= 8;  //192 / 23 = 8
    16'b11000000_00011000 : OUT <= 8;  //192 / 24 = 8
    16'b11000000_00011001 : OUT <= 7;  //192 / 25 = 7
    16'b11000000_00011010 : OUT <= 7;  //192 / 26 = 7
    16'b11000000_00011011 : OUT <= 7;  //192 / 27 = 7
    16'b11000000_00011100 : OUT <= 6;  //192 / 28 = 6
    16'b11000000_00011101 : OUT <= 6;  //192 / 29 = 6
    16'b11000000_00011110 : OUT <= 6;  //192 / 30 = 6
    16'b11000000_00011111 : OUT <= 6;  //192 / 31 = 6
    16'b11000000_00100000 : OUT <= 6;  //192 / 32 = 6
    16'b11000000_00100001 : OUT <= 5;  //192 / 33 = 5
    16'b11000000_00100010 : OUT <= 5;  //192 / 34 = 5
    16'b11000000_00100011 : OUT <= 5;  //192 / 35 = 5
    16'b11000000_00100100 : OUT <= 5;  //192 / 36 = 5
    16'b11000000_00100101 : OUT <= 5;  //192 / 37 = 5
    16'b11000000_00100110 : OUT <= 5;  //192 / 38 = 5
    16'b11000000_00100111 : OUT <= 4;  //192 / 39 = 4
    16'b11000000_00101000 : OUT <= 4;  //192 / 40 = 4
    16'b11000000_00101001 : OUT <= 4;  //192 / 41 = 4
    16'b11000000_00101010 : OUT <= 4;  //192 / 42 = 4
    16'b11000000_00101011 : OUT <= 4;  //192 / 43 = 4
    16'b11000000_00101100 : OUT <= 4;  //192 / 44 = 4
    16'b11000000_00101101 : OUT <= 4;  //192 / 45 = 4
    16'b11000000_00101110 : OUT <= 4;  //192 / 46 = 4
    16'b11000000_00101111 : OUT <= 4;  //192 / 47 = 4
    16'b11000000_00110000 : OUT <= 4;  //192 / 48 = 4
    16'b11000000_00110001 : OUT <= 3;  //192 / 49 = 3
    16'b11000000_00110010 : OUT <= 3;  //192 / 50 = 3
    16'b11000000_00110011 : OUT <= 3;  //192 / 51 = 3
    16'b11000000_00110100 : OUT <= 3;  //192 / 52 = 3
    16'b11000000_00110101 : OUT <= 3;  //192 / 53 = 3
    16'b11000000_00110110 : OUT <= 3;  //192 / 54 = 3
    16'b11000000_00110111 : OUT <= 3;  //192 / 55 = 3
    16'b11000000_00111000 : OUT <= 3;  //192 / 56 = 3
    16'b11000000_00111001 : OUT <= 3;  //192 / 57 = 3
    16'b11000000_00111010 : OUT <= 3;  //192 / 58 = 3
    16'b11000000_00111011 : OUT <= 3;  //192 / 59 = 3
    16'b11000000_00111100 : OUT <= 3;  //192 / 60 = 3
    16'b11000000_00111101 : OUT <= 3;  //192 / 61 = 3
    16'b11000000_00111110 : OUT <= 3;  //192 / 62 = 3
    16'b11000000_00111111 : OUT <= 3;  //192 / 63 = 3
    16'b11000000_01000000 : OUT <= 3;  //192 / 64 = 3
    16'b11000000_01000001 : OUT <= 2;  //192 / 65 = 2
    16'b11000000_01000010 : OUT <= 2;  //192 / 66 = 2
    16'b11000000_01000011 : OUT <= 2;  //192 / 67 = 2
    16'b11000000_01000100 : OUT <= 2;  //192 / 68 = 2
    16'b11000000_01000101 : OUT <= 2;  //192 / 69 = 2
    16'b11000000_01000110 : OUT <= 2;  //192 / 70 = 2
    16'b11000000_01000111 : OUT <= 2;  //192 / 71 = 2
    16'b11000000_01001000 : OUT <= 2;  //192 / 72 = 2
    16'b11000000_01001001 : OUT <= 2;  //192 / 73 = 2
    16'b11000000_01001010 : OUT <= 2;  //192 / 74 = 2
    16'b11000000_01001011 : OUT <= 2;  //192 / 75 = 2
    16'b11000000_01001100 : OUT <= 2;  //192 / 76 = 2
    16'b11000000_01001101 : OUT <= 2;  //192 / 77 = 2
    16'b11000000_01001110 : OUT <= 2;  //192 / 78 = 2
    16'b11000000_01001111 : OUT <= 2;  //192 / 79 = 2
    16'b11000000_01010000 : OUT <= 2;  //192 / 80 = 2
    16'b11000000_01010001 : OUT <= 2;  //192 / 81 = 2
    16'b11000000_01010010 : OUT <= 2;  //192 / 82 = 2
    16'b11000000_01010011 : OUT <= 2;  //192 / 83 = 2
    16'b11000000_01010100 : OUT <= 2;  //192 / 84 = 2
    16'b11000000_01010101 : OUT <= 2;  //192 / 85 = 2
    16'b11000000_01010110 : OUT <= 2;  //192 / 86 = 2
    16'b11000000_01010111 : OUT <= 2;  //192 / 87 = 2
    16'b11000000_01011000 : OUT <= 2;  //192 / 88 = 2
    16'b11000000_01011001 : OUT <= 2;  //192 / 89 = 2
    16'b11000000_01011010 : OUT <= 2;  //192 / 90 = 2
    16'b11000000_01011011 : OUT <= 2;  //192 / 91 = 2
    16'b11000000_01011100 : OUT <= 2;  //192 / 92 = 2
    16'b11000000_01011101 : OUT <= 2;  //192 / 93 = 2
    16'b11000000_01011110 : OUT <= 2;  //192 / 94 = 2
    16'b11000000_01011111 : OUT <= 2;  //192 / 95 = 2
    16'b11000000_01100000 : OUT <= 2;  //192 / 96 = 2
    16'b11000000_01100001 : OUT <= 1;  //192 / 97 = 1
    16'b11000000_01100010 : OUT <= 1;  //192 / 98 = 1
    16'b11000000_01100011 : OUT <= 1;  //192 / 99 = 1
    16'b11000000_01100100 : OUT <= 1;  //192 / 100 = 1
    16'b11000000_01100101 : OUT <= 1;  //192 / 101 = 1
    16'b11000000_01100110 : OUT <= 1;  //192 / 102 = 1
    16'b11000000_01100111 : OUT <= 1;  //192 / 103 = 1
    16'b11000000_01101000 : OUT <= 1;  //192 / 104 = 1
    16'b11000000_01101001 : OUT <= 1;  //192 / 105 = 1
    16'b11000000_01101010 : OUT <= 1;  //192 / 106 = 1
    16'b11000000_01101011 : OUT <= 1;  //192 / 107 = 1
    16'b11000000_01101100 : OUT <= 1;  //192 / 108 = 1
    16'b11000000_01101101 : OUT <= 1;  //192 / 109 = 1
    16'b11000000_01101110 : OUT <= 1;  //192 / 110 = 1
    16'b11000000_01101111 : OUT <= 1;  //192 / 111 = 1
    16'b11000000_01110000 : OUT <= 1;  //192 / 112 = 1
    16'b11000000_01110001 : OUT <= 1;  //192 / 113 = 1
    16'b11000000_01110010 : OUT <= 1;  //192 / 114 = 1
    16'b11000000_01110011 : OUT <= 1;  //192 / 115 = 1
    16'b11000000_01110100 : OUT <= 1;  //192 / 116 = 1
    16'b11000000_01110101 : OUT <= 1;  //192 / 117 = 1
    16'b11000000_01110110 : OUT <= 1;  //192 / 118 = 1
    16'b11000000_01110111 : OUT <= 1;  //192 / 119 = 1
    16'b11000000_01111000 : OUT <= 1;  //192 / 120 = 1
    16'b11000000_01111001 : OUT <= 1;  //192 / 121 = 1
    16'b11000000_01111010 : OUT <= 1;  //192 / 122 = 1
    16'b11000000_01111011 : OUT <= 1;  //192 / 123 = 1
    16'b11000000_01111100 : OUT <= 1;  //192 / 124 = 1
    16'b11000000_01111101 : OUT <= 1;  //192 / 125 = 1
    16'b11000000_01111110 : OUT <= 1;  //192 / 126 = 1
    16'b11000000_01111111 : OUT <= 1;  //192 / 127 = 1
    16'b11000000_10000000 : OUT <= 1;  //192 / 128 = 1
    16'b11000000_10000001 : OUT <= 1;  //192 / 129 = 1
    16'b11000000_10000010 : OUT <= 1;  //192 / 130 = 1
    16'b11000000_10000011 : OUT <= 1;  //192 / 131 = 1
    16'b11000000_10000100 : OUT <= 1;  //192 / 132 = 1
    16'b11000000_10000101 : OUT <= 1;  //192 / 133 = 1
    16'b11000000_10000110 : OUT <= 1;  //192 / 134 = 1
    16'b11000000_10000111 : OUT <= 1;  //192 / 135 = 1
    16'b11000000_10001000 : OUT <= 1;  //192 / 136 = 1
    16'b11000000_10001001 : OUT <= 1;  //192 / 137 = 1
    16'b11000000_10001010 : OUT <= 1;  //192 / 138 = 1
    16'b11000000_10001011 : OUT <= 1;  //192 / 139 = 1
    16'b11000000_10001100 : OUT <= 1;  //192 / 140 = 1
    16'b11000000_10001101 : OUT <= 1;  //192 / 141 = 1
    16'b11000000_10001110 : OUT <= 1;  //192 / 142 = 1
    16'b11000000_10001111 : OUT <= 1;  //192 / 143 = 1
    16'b11000000_10010000 : OUT <= 1;  //192 / 144 = 1
    16'b11000000_10010001 : OUT <= 1;  //192 / 145 = 1
    16'b11000000_10010010 : OUT <= 1;  //192 / 146 = 1
    16'b11000000_10010011 : OUT <= 1;  //192 / 147 = 1
    16'b11000000_10010100 : OUT <= 1;  //192 / 148 = 1
    16'b11000000_10010101 : OUT <= 1;  //192 / 149 = 1
    16'b11000000_10010110 : OUT <= 1;  //192 / 150 = 1
    16'b11000000_10010111 : OUT <= 1;  //192 / 151 = 1
    16'b11000000_10011000 : OUT <= 1;  //192 / 152 = 1
    16'b11000000_10011001 : OUT <= 1;  //192 / 153 = 1
    16'b11000000_10011010 : OUT <= 1;  //192 / 154 = 1
    16'b11000000_10011011 : OUT <= 1;  //192 / 155 = 1
    16'b11000000_10011100 : OUT <= 1;  //192 / 156 = 1
    16'b11000000_10011101 : OUT <= 1;  //192 / 157 = 1
    16'b11000000_10011110 : OUT <= 1;  //192 / 158 = 1
    16'b11000000_10011111 : OUT <= 1;  //192 / 159 = 1
    16'b11000000_10100000 : OUT <= 1;  //192 / 160 = 1
    16'b11000000_10100001 : OUT <= 1;  //192 / 161 = 1
    16'b11000000_10100010 : OUT <= 1;  //192 / 162 = 1
    16'b11000000_10100011 : OUT <= 1;  //192 / 163 = 1
    16'b11000000_10100100 : OUT <= 1;  //192 / 164 = 1
    16'b11000000_10100101 : OUT <= 1;  //192 / 165 = 1
    16'b11000000_10100110 : OUT <= 1;  //192 / 166 = 1
    16'b11000000_10100111 : OUT <= 1;  //192 / 167 = 1
    16'b11000000_10101000 : OUT <= 1;  //192 / 168 = 1
    16'b11000000_10101001 : OUT <= 1;  //192 / 169 = 1
    16'b11000000_10101010 : OUT <= 1;  //192 / 170 = 1
    16'b11000000_10101011 : OUT <= 1;  //192 / 171 = 1
    16'b11000000_10101100 : OUT <= 1;  //192 / 172 = 1
    16'b11000000_10101101 : OUT <= 1;  //192 / 173 = 1
    16'b11000000_10101110 : OUT <= 1;  //192 / 174 = 1
    16'b11000000_10101111 : OUT <= 1;  //192 / 175 = 1
    16'b11000000_10110000 : OUT <= 1;  //192 / 176 = 1
    16'b11000000_10110001 : OUT <= 1;  //192 / 177 = 1
    16'b11000000_10110010 : OUT <= 1;  //192 / 178 = 1
    16'b11000000_10110011 : OUT <= 1;  //192 / 179 = 1
    16'b11000000_10110100 : OUT <= 1;  //192 / 180 = 1
    16'b11000000_10110101 : OUT <= 1;  //192 / 181 = 1
    16'b11000000_10110110 : OUT <= 1;  //192 / 182 = 1
    16'b11000000_10110111 : OUT <= 1;  //192 / 183 = 1
    16'b11000000_10111000 : OUT <= 1;  //192 / 184 = 1
    16'b11000000_10111001 : OUT <= 1;  //192 / 185 = 1
    16'b11000000_10111010 : OUT <= 1;  //192 / 186 = 1
    16'b11000000_10111011 : OUT <= 1;  //192 / 187 = 1
    16'b11000000_10111100 : OUT <= 1;  //192 / 188 = 1
    16'b11000000_10111101 : OUT <= 1;  //192 / 189 = 1
    16'b11000000_10111110 : OUT <= 1;  //192 / 190 = 1
    16'b11000000_10111111 : OUT <= 1;  //192 / 191 = 1
    16'b11000000_11000000 : OUT <= 1;  //192 / 192 = 1
    16'b11000000_11000001 : OUT <= 0;  //192 / 193 = 0
    16'b11000000_11000010 : OUT <= 0;  //192 / 194 = 0
    16'b11000000_11000011 : OUT <= 0;  //192 / 195 = 0
    16'b11000000_11000100 : OUT <= 0;  //192 / 196 = 0
    16'b11000000_11000101 : OUT <= 0;  //192 / 197 = 0
    16'b11000000_11000110 : OUT <= 0;  //192 / 198 = 0
    16'b11000000_11000111 : OUT <= 0;  //192 / 199 = 0
    16'b11000000_11001000 : OUT <= 0;  //192 / 200 = 0
    16'b11000000_11001001 : OUT <= 0;  //192 / 201 = 0
    16'b11000000_11001010 : OUT <= 0;  //192 / 202 = 0
    16'b11000000_11001011 : OUT <= 0;  //192 / 203 = 0
    16'b11000000_11001100 : OUT <= 0;  //192 / 204 = 0
    16'b11000000_11001101 : OUT <= 0;  //192 / 205 = 0
    16'b11000000_11001110 : OUT <= 0;  //192 / 206 = 0
    16'b11000000_11001111 : OUT <= 0;  //192 / 207 = 0
    16'b11000000_11010000 : OUT <= 0;  //192 / 208 = 0
    16'b11000000_11010001 : OUT <= 0;  //192 / 209 = 0
    16'b11000000_11010010 : OUT <= 0;  //192 / 210 = 0
    16'b11000000_11010011 : OUT <= 0;  //192 / 211 = 0
    16'b11000000_11010100 : OUT <= 0;  //192 / 212 = 0
    16'b11000000_11010101 : OUT <= 0;  //192 / 213 = 0
    16'b11000000_11010110 : OUT <= 0;  //192 / 214 = 0
    16'b11000000_11010111 : OUT <= 0;  //192 / 215 = 0
    16'b11000000_11011000 : OUT <= 0;  //192 / 216 = 0
    16'b11000000_11011001 : OUT <= 0;  //192 / 217 = 0
    16'b11000000_11011010 : OUT <= 0;  //192 / 218 = 0
    16'b11000000_11011011 : OUT <= 0;  //192 / 219 = 0
    16'b11000000_11011100 : OUT <= 0;  //192 / 220 = 0
    16'b11000000_11011101 : OUT <= 0;  //192 / 221 = 0
    16'b11000000_11011110 : OUT <= 0;  //192 / 222 = 0
    16'b11000000_11011111 : OUT <= 0;  //192 / 223 = 0
    16'b11000000_11100000 : OUT <= 0;  //192 / 224 = 0
    16'b11000000_11100001 : OUT <= 0;  //192 / 225 = 0
    16'b11000000_11100010 : OUT <= 0;  //192 / 226 = 0
    16'b11000000_11100011 : OUT <= 0;  //192 / 227 = 0
    16'b11000000_11100100 : OUT <= 0;  //192 / 228 = 0
    16'b11000000_11100101 : OUT <= 0;  //192 / 229 = 0
    16'b11000000_11100110 : OUT <= 0;  //192 / 230 = 0
    16'b11000000_11100111 : OUT <= 0;  //192 / 231 = 0
    16'b11000000_11101000 : OUT <= 0;  //192 / 232 = 0
    16'b11000000_11101001 : OUT <= 0;  //192 / 233 = 0
    16'b11000000_11101010 : OUT <= 0;  //192 / 234 = 0
    16'b11000000_11101011 : OUT <= 0;  //192 / 235 = 0
    16'b11000000_11101100 : OUT <= 0;  //192 / 236 = 0
    16'b11000000_11101101 : OUT <= 0;  //192 / 237 = 0
    16'b11000000_11101110 : OUT <= 0;  //192 / 238 = 0
    16'b11000000_11101111 : OUT <= 0;  //192 / 239 = 0
    16'b11000000_11110000 : OUT <= 0;  //192 / 240 = 0
    16'b11000000_11110001 : OUT <= 0;  //192 / 241 = 0
    16'b11000000_11110010 : OUT <= 0;  //192 / 242 = 0
    16'b11000000_11110011 : OUT <= 0;  //192 / 243 = 0
    16'b11000000_11110100 : OUT <= 0;  //192 / 244 = 0
    16'b11000000_11110101 : OUT <= 0;  //192 / 245 = 0
    16'b11000000_11110110 : OUT <= 0;  //192 / 246 = 0
    16'b11000000_11110111 : OUT <= 0;  //192 / 247 = 0
    16'b11000000_11111000 : OUT <= 0;  //192 / 248 = 0
    16'b11000000_11111001 : OUT <= 0;  //192 / 249 = 0
    16'b11000000_11111010 : OUT <= 0;  //192 / 250 = 0
    16'b11000000_11111011 : OUT <= 0;  //192 / 251 = 0
    16'b11000000_11111100 : OUT <= 0;  //192 / 252 = 0
    16'b11000000_11111101 : OUT <= 0;  //192 / 253 = 0
    16'b11000000_11111110 : OUT <= 0;  //192 / 254 = 0
    16'b11000000_11111111 : OUT <= 0;  //192 / 255 = 0
    16'b11000001_00000000 : OUT <= 0;  //193 / 0 = 0
    16'b11000001_00000001 : OUT <= 193;  //193 / 1 = 193
    16'b11000001_00000010 : OUT <= 96;  //193 / 2 = 96
    16'b11000001_00000011 : OUT <= 64;  //193 / 3 = 64
    16'b11000001_00000100 : OUT <= 48;  //193 / 4 = 48
    16'b11000001_00000101 : OUT <= 38;  //193 / 5 = 38
    16'b11000001_00000110 : OUT <= 32;  //193 / 6 = 32
    16'b11000001_00000111 : OUT <= 27;  //193 / 7 = 27
    16'b11000001_00001000 : OUT <= 24;  //193 / 8 = 24
    16'b11000001_00001001 : OUT <= 21;  //193 / 9 = 21
    16'b11000001_00001010 : OUT <= 19;  //193 / 10 = 19
    16'b11000001_00001011 : OUT <= 17;  //193 / 11 = 17
    16'b11000001_00001100 : OUT <= 16;  //193 / 12 = 16
    16'b11000001_00001101 : OUT <= 14;  //193 / 13 = 14
    16'b11000001_00001110 : OUT <= 13;  //193 / 14 = 13
    16'b11000001_00001111 : OUT <= 12;  //193 / 15 = 12
    16'b11000001_00010000 : OUT <= 12;  //193 / 16 = 12
    16'b11000001_00010001 : OUT <= 11;  //193 / 17 = 11
    16'b11000001_00010010 : OUT <= 10;  //193 / 18 = 10
    16'b11000001_00010011 : OUT <= 10;  //193 / 19 = 10
    16'b11000001_00010100 : OUT <= 9;  //193 / 20 = 9
    16'b11000001_00010101 : OUT <= 9;  //193 / 21 = 9
    16'b11000001_00010110 : OUT <= 8;  //193 / 22 = 8
    16'b11000001_00010111 : OUT <= 8;  //193 / 23 = 8
    16'b11000001_00011000 : OUT <= 8;  //193 / 24 = 8
    16'b11000001_00011001 : OUT <= 7;  //193 / 25 = 7
    16'b11000001_00011010 : OUT <= 7;  //193 / 26 = 7
    16'b11000001_00011011 : OUT <= 7;  //193 / 27 = 7
    16'b11000001_00011100 : OUT <= 6;  //193 / 28 = 6
    16'b11000001_00011101 : OUT <= 6;  //193 / 29 = 6
    16'b11000001_00011110 : OUT <= 6;  //193 / 30 = 6
    16'b11000001_00011111 : OUT <= 6;  //193 / 31 = 6
    16'b11000001_00100000 : OUT <= 6;  //193 / 32 = 6
    16'b11000001_00100001 : OUT <= 5;  //193 / 33 = 5
    16'b11000001_00100010 : OUT <= 5;  //193 / 34 = 5
    16'b11000001_00100011 : OUT <= 5;  //193 / 35 = 5
    16'b11000001_00100100 : OUT <= 5;  //193 / 36 = 5
    16'b11000001_00100101 : OUT <= 5;  //193 / 37 = 5
    16'b11000001_00100110 : OUT <= 5;  //193 / 38 = 5
    16'b11000001_00100111 : OUT <= 4;  //193 / 39 = 4
    16'b11000001_00101000 : OUT <= 4;  //193 / 40 = 4
    16'b11000001_00101001 : OUT <= 4;  //193 / 41 = 4
    16'b11000001_00101010 : OUT <= 4;  //193 / 42 = 4
    16'b11000001_00101011 : OUT <= 4;  //193 / 43 = 4
    16'b11000001_00101100 : OUT <= 4;  //193 / 44 = 4
    16'b11000001_00101101 : OUT <= 4;  //193 / 45 = 4
    16'b11000001_00101110 : OUT <= 4;  //193 / 46 = 4
    16'b11000001_00101111 : OUT <= 4;  //193 / 47 = 4
    16'b11000001_00110000 : OUT <= 4;  //193 / 48 = 4
    16'b11000001_00110001 : OUT <= 3;  //193 / 49 = 3
    16'b11000001_00110010 : OUT <= 3;  //193 / 50 = 3
    16'b11000001_00110011 : OUT <= 3;  //193 / 51 = 3
    16'b11000001_00110100 : OUT <= 3;  //193 / 52 = 3
    16'b11000001_00110101 : OUT <= 3;  //193 / 53 = 3
    16'b11000001_00110110 : OUT <= 3;  //193 / 54 = 3
    16'b11000001_00110111 : OUT <= 3;  //193 / 55 = 3
    16'b11000001_00111000 : OUT <= 3;  //193 / 56 = 3
    16'b11000001_00111001 : OUT <= 3;  //193 / 57 = 3
    16'b11000001_00111010 : OUT <= 3;  //193 / 58 = 3
    16'b11000001_00111011 : OUT <= 3;  //193 / 59 = 3
    16'b11000001_00111100 : OUT <= 3;  //193 / 60 = 3
    16'b11000001_00111101 : OUT <= 3;  //193 / 61 = 3
    16'b11000001_00111110 : OUT <= 3;  //193 / 62 = 3
    16'b11000001_00111111 : OUT <= 3;  //193 / 63 = 3
    16'b11000001_01000000 : OUT <= 3;  //193 / 64 = 3
    16'b11000001_01000001 : OUT <= 2;  //193 / 65 = 2
    16'b11000001_01000010 : OUT <= 2;  //193 / 66 = 2
    16'b11000001_01000011 : OUT <= 2;  //193 / 67 = 2
    16'b11000001_01000100 : OUT <= 2;  //193 / 68 = 2
    16'b11000001_01000101 : OUT <= 2;  //193 / 69 = 2
    16'b11000001_01000110 : OUT <= 2;  //193 / 70 = 2
    16'b11000001_01000111 : OUT <= 2;  //193 / 71 = 2
    16'b11000001_01001000 : OUT <= 2;  //193 / 72 = 2
    16'b11000001_01001001 : OUT <= 2;  //193 / 73 = 2
    16'b11000001_01001010 : OUT <= 2;  //193 / 74 = 2
    16'b11000001_01001011 : OUT <= 2;  //193 / 75 = 2
    16'b11000001_01001100 : OUT <= 2;  //193 / 76 = 2
    16'b11000001_01001101 : OUT <= 2;  //193 / 77 = 2
    16'b11000001_01001110 : OUT <= 2;  //193 / 78 = 2
    16'b11000001_01001111 : OUT <= 2;  //193 / 79 = 2
    16'b11000001_01010000 : OUT <= 2;  //193 / 80 = 2
    16'b11000001_01010001 : OUT <= 2;  //193 / 81 = 2
    16'b11000001_01010010 : OUT <= 2;  //193 / 82 = 2
    16'b11000001_01010011 : OUT <= 2;  //193 / 83 = 2
    16'b11000001_01010100 : OUT <= 2;  //193 / 84 = 2
    16'b11000001_01010101 : OUT <= 2;  //193 / 85 = 2
    16'b11000001_01010110 : OUT <= 2;  //193 / 86 = 2
    16'b11000001_01010111 : OUT <= 2;  //193 / 87 = 2
    16'b11000001_01011000 : OUT <= 2;  //193 / 88 = 2
    16'b11000001_01011001 : OUT <= 2;  //193 / 89 = 2
    16'b11000001_01011010 : OUT <= 2;  //193 / 90 = 2
    16'b11000001_01011011 : OUT <= 2;  //193 / 91 = 2
    16'b11000001_01011100 : OUT <= 2;  //193 / 92 = 2
    16'b11000001_01011101 : OUT <= 2;  //193 / 93 = 2
    16'b11000001_01011110 : OUT <= 2;  //193 / 94 = 2
    16'b11000001_01011111 : OUT <= 2;  //193 / 95 = 2
    16'b11000001_01100000 : OUT <= 2;  //193 / 96 = 2
    16'b11000001_01100001 : OUT <= 1;  //193 / 97 = 1
    16'b11000001_01100010 : OUT <= 1;  //193 / 98 = 1
    16'b11000001_01100011 : OUT <= 1;  //193 / 99 = 1
    16'b11000001_01100100 : OUT <= 1;  //193 / 100 = 1
    16'b11000001_01100101 : OUT <= 1;  //193 / 101 = 1
    16'b11000001_01100110 : OUT <= 1;  //193 / 102 = 1
    16'b11000001_01100111 : OUT <= 1;  //193 / 103 = 1
    16'b11000001_01101000 : OUT <= 1;  //193 / 104 = 1
    16'b11000001_01101001 : OUT <= 1;  //193 / 105 = 1
    16'b11000001_01101010 : OUT <= 1;  //193 / 106 = 1
    16'b11000001_01101011 : OUT <= 1;  //193 / 107 = 1
    16'b11000001_01101100 : OUT <= 1;  //193 / 108 = 1
    16'b11000001_01101101 : OUT <= 1;  //193 / 109 = 1
    16'b11000001_01101110 : OUT <= 1;  //193 / 110 = 1
    16'b11000001_01101111 : OUT <= 1;  //193 / 111 = 1
    16'b11000001_01110000 : OUT <= 1;  //193 / 112 = 1
    16'b11000001_01110001 : OUT <= 1;  //193 / 113 = 1
    16'b11000001_01110010 : OUT <= 1;  //193 / 114 = 1
    16'b11000001_01110011 : OUT <= 1;  //193 / 115 = 1
    16'b11000001_01110100 : OUT <= 1;  //193 / 116 = 1
    16'b11000001_01110101 : OUT <= 1;  //193 / 117 = 1
    16'b11000001_01110110 : OUT <= 1;  //193 / 118 = 1
    16'b11000001_01110111 : OUT <= 1;  //193 / 119 = 1
    16'b11000001_01111000 : OUT <= 1;  //193 / 120 = 1
    16'b11000001_01111001 : OUT <= 1;  //193 / 121 = 1
    16'b11000001_01111010 : OUT <= 1;  //193 / 122 = 1
    16'b11000001_01111011 : OUT <= 1;  //193 / 123 = 1
    16'b11000001_01111100 : OUT <= 1;  //193 / 124 = 1
    16'b11000001_01111101 : OUT <= 1;  //193 / 125 = 1
    16'b11000001_01111110 : OUT <= 1;  //193 / 126 = 1
    16'b11000001_01111111 : OUT <= 1;  //193 / 127 = 1
    16'b11000001_10000000 : OUT <= 1;  //193 / 128 = 1
    16'b11000001_10000001 : OUT <= 1;  //193 / 129 = 1
    16'b11000001_10000010 : OUT <= 1;  //193 / 130 = 1
    16'b11000001_10000011 : OUT <= 1;  //193 / 131 = 1
    16'b11000001_10000100 : OUT <= 1;  //193 / 132 = 1
    16'b11000001_10000101 : OUT <= 1;  //193 / 133 = 1
    16'b11000001_10000110 : OUT <= 1;  //193 / 134 = 1
    16'b11000001_10000111 : OUT <= 1;  //193 / 135 = 1
    16'b11000001_10001000 : OUT <= 1;  //193 / 136 = 1
    16'b11000001_10001001 : OUT <= 1;  //193 / 137 = 1
    16'b11000001_10001010 : OUT <= 1;  //193 / 138 = 1
    16'b11000001_10001011 : OUT <= 1;  //193 / 139 = 1
    16'b11000001_10001100 : OUT <= 1;  //193 / 140 = 1
    16'b11000001_10001101 : OUT <= 1;  //193 / 141 = 1
    16'b11000001_10001110 : OUT <= 1;  //193 / 142 = 1
    16'b11000001_10001111 : OUT <= 1;  //193 / 143 = 1
    16'b11000001_10010000 : OUT <= 1;  //193 / 144 = 1
    16'b11000001_10010001 : OUT <= 1;  //193 / 145 = 1
    16'b11000001_10010010 : OUT <= 1;  //193 / 146 = 1
    16'b11000001_10010011 : OUT <= 1;  //193 / 147 = 1
    16'b11000001_10010100 : OUT <= 1;  //193 / 148 = 1
    16'b11000001_10010101 : OUT <= 1;  //193 / 149 = 1
    16'b11000001_10010110 : OUT <= 1;  //193 / 150 = 1
    16'b11000001_10010111 : OUT <= 1;  //193 / 151 = 1
    16'b11000001_10011000 : OUT <= 1;  //193 / 152 = 1
    16'b11000001_10011001 : OUT <= 1;  //193 / 153 = 1
    16'b11000001_10011010 : OUT <= 1;  //193 / 154 = 1
    16'b11000001_10011011 : OUT <= 1;  //193 / 155 = 1
    16'b11000001_10011100 : OUT <= 1;  //193 / 156 = 1
    16'b11000001_10011101 : OUT <= 1;  //193 / 157 = 1
    16'b11000001_10011110 : OUT <= 1;  //193 / 158 = 1
    16'b11000001_10011111 : OUT <= 1;  //193 / 159 = 1
    16'b11000001_10100000 : OUT <= 1;  //193 / 160 = 1
    16'b11000001_10100001 : OUT <= 1;  //193 / 161 = 1
    16'b11000001_10100010 : OUT <= 1;  //193 / 162 = 1
    16'b11000001_10100011 : OUT <= 1;  //193 / 163 = 1
    16'b11000001_10100100 : OUT <= 1;  //193 / 164 = 1
    16'b11000001_10100101 : OUT <= 1;  //193 / 165 = 1
    16'b11000001_10100110 : OUT <= 1;  //193 / 166 = 1
    16'b11000001_10100111 : OUT <= 1;  //193 / 167 = 1
    16'b11000001_10101000 : OUT <= 1;  //193 / 168 = 1
    16'b11000001_10101001 : OUT <= 1;  //193 / 169 = 1
    16'b11000001_10101010 : OUT <= 1;  //193 / 170 = 1
    16'b11000001_10101011 : OUT <= 1;  //193 / 171 = 1
    16'b11000001_10101100 : OUT <= 1;  //193 / 172 = 1
    16'b11000001_10101101 : OUT <= 1;  //193 / 173 = 1
    16'b11000001_10101110 : OUT <= 1;  //193 / 174 = 1
    16'b11000001_10101111 : OUT <= 1;  //193 / 175 = 1
    16'b11000001_10110000 : OUT <= 1;  //193 / 176 = 1
    16'b11000001_10110001 : OUT <= 1;  //193 / 177 = 1
    16'b11000001_10110010 : OUT <= 1;  //193 / 178 = 1
    16'b11000001_10110011 : OUT <= 1;  //193 / 179 = 1
    16'b11000001_10110100 : OUT <= 1;  //193 / 180 = 1
    16'b11000001_10110101 : OUT <= 1;  //193 / 181 = 1
    16'b11000001_10110110 : OUT <= 1;  //193 / 182 = 1
    16'b11000001_10110111 : OUT <= 1;  //193 / 183 = 1
    16'b11000001_10111000 : OUT <= 1;  //193 / 184 = 1
    16'b11000001_10111001 : OUT <= 1;  //193 / 185 = 1
    16'b11000001_10111010 : OUT <= 1;  //193 / 186 = 1
    16'b11000001_10111011 : OUT <= 1;  //193 / 187 = 1
    16'b11000001_10111100 : OUT <= 1;  //193 / 188 = 1
    16'b11000001_10111101 : OUT <= 1;  //193 / 189 = 1
    16'b11000001_10111110 : OUT <= 1;  //193 / 190 = 1
    16'b11000001_10111111 : OUT <= 1;  //193 / 191 = 1
    16'b11000001_11000000 : OUT <= 1;  //193 / 192 = 1
    16'b11000001_11000001 : OUT <= 1;  //193 / 193 = 1
    16'b11000001_11000010 : OUT <= 0;  //193 / 194 = 0
    16'b11000001_11000011 : OUT <= 0;  //193 / 195 = 0
    16'b11000001_11000100 : OUT <= 0;  //193 / 196 = 0
    16'b11000001_11000101 : OUT <= 0;  //193 / 197 = 0
    16'b11000001_11000110 : OUT <= 0;  //193 / 198 = 0
    16'b11000001_11000111 : OUT <= 0;  //193 / 199 = 0
    16'b11000001_11001000 : OUT <= 0;  //193 / 200 = 0
    16'b11000001_11001001 : OUT <= 0;  //193 / 201 = 0
    16'b11000001_11001010 : OUT <= 0;  //193 / 202 = 0
    16'b11000001_11001011 : OUT <= 0;  //193 / 203 = 0
    16'b11000001_11001100 : OUT <= 0;  //193 / 204 = 0
    16'b11000001_11001101 : OUT <= 0;  //193 / 205 = 0
    16'b11000001_11001110 : OUT <= 0;  //193 / 206 = 0
    16'b11000001_11001111 : OUT <= 0;  //193 / 207 = 0
    16'b11000001_11010000 : OUT <= 0;  //193 / 208 = 0
    16'b11000001_11010001 : OUT <= 0;  //193 / 209 = 0
    16'b11000001_11010010 : OUT <= 0;  //193 / 210 = 0
    16'b11000001_11010011 : OUT <= 0;  //193 / 211 = 0
    16'b11000001_11010100 : OUT <= 0;  //193 / 212 = 0
    16'b11000001_11010101 : OUT <= 0;  //193 / 213 = 0
    16'b11000001_11010110 : OUT <= 0;  //193 / 214 = 0
    16'b11000001_11010111 : OUT <= 0;  //193 / 215 = 0
    16'b11000001_11011000 : OUT <= 0;  //193 / 216 = 0
    16'b11000001_11011001 : OUT <= 0;  //193 / 217 = 0
    16'b11000001_11011010 : OUT <= 0;  //193 / 218 = 0
    16'b11000001_11011011 : OUT <= 0;  //193 / 219 = 0
    16'b11000001_11011100 : OUT <= 0;  //193 / 220 = 0
    16'b11000001_11011101 : OUT <= 0;  //193 / 221 = 0
    16'b11000001_11011110 : OUT <= 0;  //193 / 222 = 0
    16'b11000001_11011111 : OUT <= 0;  //193 / 223 = 0
    16'b11000001_11100000 : OUT <= 0;  //193 / 224 = 0
    16'b11000001_11100001 : OUT <= 0;  //193 / 225 = 0
    16'b11000001_11100010 : OUT <= 0;  //193 / 226 = 0
    16'b11000001_11100011 : OUT <= 0;  //193 / 227 = 0
    16'b11000001_11100100 : OUT <= 0;  //193 / 228 = 0
    16'b11000001_11100101 : OUT <= 0;  //193 / 229 = 0
    16'b11000001_11100110 : OUT <= 0;  //193 / 230 = 0
    16'b11000001_11100111 : OUT <= 0;  //193 / 231 = 0
    16'b11000001_11101000 : OUT <= 0;  //193 / 232 = 0
    16'b11000001_11101001 : OUT <= 0;  //193 / 233 = 0
    16'b11000001_11101010 : OUT <= 0;  //193 / 234 = 0
    16'b11000001_11101011 : OUT <= 0;  //193 / 235 = 0
    16'b11000001_11101100 : OUT <= 0;  //193 / 236 = 0
    16'b11000001_11101101 : OUT <= 0;  //193 / 237 = 0
    16'b11000001_11101110 : OUT <= 0;  //193 / 238 = 0
    16'b11000001_11101111 : OUT <= 0;  //193 / 239 = 0
    16'b11000001_11110000 : OUT <= 0;  //193 / 240 = 0
    16'b11000001_11110001 : OUT <= 0;  //193 / 241 = 0
    16'b11000001_11110010 : OUT <= 0;  //193 / 242 = 0
    16'b11000001_11110011 : OUT <= 0;  //193 / 243 = 0
    16'b11000001_11110100 : OUT <= 0;  //193 / 244 = 0
    16'b11000001_11110101 : OUT <= 0;  //193 / 245 = 0
    16'b11000001_11110110 : OUT <= 0;  //193 / 246 = 0
    16'b11000001_11110111 : OUT <= 0;  //193 / 247 = 0
    16'b11000001_11111000 : OUT <= 0;  //193 / 248 = 0
    16'b11000001_11111001 : OUT <= 0;  //193 / 249 = 0
    16'b11000001_11111010 : OUT <= 0;  //193 / 250 = 0
    16'b11000001_11111011 : OUT <= 0;  //193 / 251 = 0
    16'b11000001_11111100 : OUT <= 0;  //193 / 252 = 0
    16'b11000001_11111101 : OUT <= 0;  //193 / 253 = 0
    16'b11000001_11111110 : OUT <= 0;  //193 / 254 = 0
    16'b11000001_11111111 : OUT <= 0;  //193 / 255 = 0
    16'b11000010_00000000 : OUT <= 0;  //194 / 0 = 0
    16'b11000010_00000001 : OUT <= 194;  //194 / 1 = 194
    16'b11000010_00000010 : OUT <= 97;  //194 / 2 = 97
    16'b11000010_00000011 : OUT <= 64;  //194 / 3 = 64
    16'b11000010_00000100 : OUT <= 48;  //194 / 4 = 48
    16'b11000010_00000101 : OUT <= 38;  //194 / 5 = 38
    16'b11000010_00000110 : OUT <= 32;  //194 / 6 = 32
    16'b11000010_00000111 : OUT <= 27;  //194 / 7 = 27
    16'b11000010_00001000 : OUT <= 24;  //194 / 8 = 24
    16'b11000010_00001001 : OUT <= 21;  //194 / 9 = 21
    16'b11000010_00001010 : OUT <= 19;  //194 / 10 = 19
    16'b11000010_00001011 : OUT <= 17;  //194 / 11 = 17
    16'b11000010_00001100 : OUT <= 16;  //194 / 12 = 16
    16'b11000010_00001101 : OUT <= 14;  //194 / 13 = 14
    16'b11000010_00001110 : OUT <= 13;  //194 / 14 = 13
    16'b11000010_00001111 : OUT <= 12;  //194 / 15 = 12
    16'b11000010_00010000 : OUT <= 12;  //194 / 16 = 12
    16'b11000010_00010001 : OUT <= 11;  //194 / 17 = 11
    16'b11000010_00010010 : OUT <= 10;  //194 / 18 = 10
    16'b11000010_00010011 : OUT <= 10;  //194 / 19 = 10
    16'b11000010_00010100 : OUT <= 9;  //194 / 20 = 9
    16'b11000010_00010101 : OUT <= 9;  //194 / 21 = 9
    16'b11000010_00010110 : OUT <= 8;  //194 / 22 = 8
    16'b11000010_00010111 : OUT <= 8;  //194 / 23 = 8
    16'b11000010_00011000 : OUT <= 8;  //194 / 24 = 8
    16'b11000010_00011001 : OUT <= 7;  //194 / 25 = 7
    16'b11000010_00011010 : OUT <= 7;  //194 / 26 = 7
    16'b11000010_00011011 : OUT <= 7;  //194 / 27 = 7
    16'b11000010_00011100 : OUT <= 6;  //194 / 28 = 6
    16'b11000010_00011101 : OUT <= 6;  //194 / 29 = 6
    16'b11000010_00011110 : OUT <= 6;  //194 / 30 = 6
    16'b11000010_00011111 : OUT <= 6;  //194 / 31 = 6
    16'b11000010_00100000 : OUT <= 6;  //194 / 32 = 6
    16'b11000010_00100001 : OUT <= 5;  //194 / 33 = 5
    16'b11000010_00100010 : OUT <= 5;  //194 / 34 = 5
    16'b11000010_00100011 : OUT <= 5;  //194 / 35 = 5
    16'b11000010_00100100 : OUT <= 5;  //194 / 36 = 5
    16'b11000010_00100101 : OUT <= 5;  //194 / 37 = 5
    16'b11000010_00100110 : OUT <= 5;  //194 / 38 = 5
    16'b11000010_00100111 : OUT <= 4;  //194 / 39 = 4
    16'b11000010_00101000 : OUT <= 4;  //194 / 40 = 4
    16'b11000010_00101001 : OUT <= 4;  //194 / 41 = 4
    16'b11000010_00101010 : OUT <= 4;  //194 / 42 = 4
    16'b11000010_00101011 : OUT <= 4;  //194 / 43 = 4
    16'b11000010_00101100 : OUT <= 4;  //194 / 44 = 4
    16'b11000010_00101101 : OUT <= 4;  //194 / 45 = 4
    16'b11000010_00101110 : OUT <= 4;  //194 / 46 = 4
    16'b11000010_00101111 : OUT <= 4;  //194 / 47 = 4
    16'b11000010_00110000 : OUT <= 4;  //194 / 48 = 4
    16'b11000010_00110001 : OUT <= 3;  //194 / 49 = 3
    16'b11000010_00110010 : OUT <= 3;  //194 / 50 = 3
    16'b11000010_00110011 : OUT <= 3;  //194 / 51 = 3
    16'b11000010_00110100 : OUT <= 3;  //194 / 52 = 3
    16'b11000010_00110101 : OUT <= 3;  //194 / 53 = 3
    16'b11000010_00110110 : OUT <= 3;  //194 / 54 = 3
    16'b11000010_00110111 : OUT <= 3;  //194 / 55 = 3
    16'b11000010_00111000 : OUT <= 3;  //194 / 56 = 3
    16'b11000010_00111001 : OUT <= 3;  //194 / 57 = 3
    16'b11000010_00111010 : OUT <= 3;  //194 / 58 = 3
    16'b11000010_00111011 : OUT <= 3;  //194 / 59 = 3
    16'b11000010_00111100 : OUT <= 3;  //194 / 60 = 3
    16'b11000010_00111101 : OUT <= 3;  //194 / 61 = 3
    16'b11000010_00111110 : OUT <= 3;  //194 / 62 = 3
    16'b11000010_00111111 : OUT <= 3;  //194 / 63 = 3
    16'b11000010_01000000 : OUT <= 3;  //194 / 64 = 3
    16'b11000010_01000001 : OUT <= 2;  //194 / 65 = 2
    16'b11000010_01000010 : OUT <= 2;  //194 / 66 = 2
    16'b11000010_01000011 : OUT <= 2;  //194 / 67 = 2
    16'b11000010_01000100 : OUT <= 2;  //194 / 68 = 2
    16'b11000010_01000101 : OUT <= 2;  //194 / 69 = 2
    16'b11000010_01000110 : OUT <= 2;  //194 / 70 = 2
    16'b11000010_01000111 : OUT <= 2;  //194 / 71 = 2
    16'b11000010_01001000 : OUT <= 2;  //194 / 72 = 2
    16'b11000010_01001001 : OUT <= 2;  //194 / 73 = 2
    16'b11000010_01001010 : OUT <= 2;  //194 / 74 = 2
    16'b11000010_01001011 : OUT <= 2;  //194 / 75 = 2
    16'b11000010_01001100 : OUT <= 2;  //194 / 76 = 2
    16'b11000010_01001101 : OUT <= 2;  //194 / 77 = 2
    16'b11000010_01001110 : OUT <= 2;  //194 / 78 = 2
    16'b11000010_01001111 : OUT <= 2;  //194 / 79 = 2
    16'b11000010_01010000 : OUT <= 2;  //194 / 80 = 2
    16'b11000010_01010001 : OUT <= 2;  //194 / 81 = 2
    16'b11000010_01010010 : OUT <= 2;  //194 / 82 = 2
    16'b11000010_01010011 : OUT <= 2;  //194 / 83 = 2
    16'b11000010_01010100 : OUT <= 2;  //194 / 84 = 2
    16'b11000010_01010101 : OUT <= 2;  //194 / 85 = 2
    16'b11000010_01010110 : OUT <= 2;  //194 / 86 = 2
    16'b11000010_01010111 : OUT <= 2;  //194 / 87 = 2
    16'b11000010_01011000 : OUT <= 2;  //194 / 88 = 2
    16'b11000010_01011001 : OUT <= 2;  //194 / 89 = 2
    16'b11000010_01011010 : OUT <= 2;  //194 / 90 = 2
    16'b11000010_01011011 : OUT <= 2;  //194 / 91 = 2
    16'b11000010_01011100 : OUT <= 2;  //194 / 92 = 2
    16'b11000010_01011101 : OUT <= 2;  //194 / 93 = 2
    16'b11000010_01011110 : OUT <= 2;  //194 / 94 = 2
    16'b11000010_01011111 : OUT <= 2;  //194 / 95 = 2
    16'b11000010_01100000 : OUT <= 2;  //194 / 96 = 2
    16'b11000010_01100001 : OUT <= 2;  //194 / 97 = 2
    16'b11000010_01100010 : OUT <= 1;  //194 / 98 = 1
    16'b11000010_01100011 : OUT <= 1;  //194 / 99 = 1
    16'b11000010_01100100 : OUT <= 1;  //194 / 100 = 1
    16'b11000010_01100101 : OUT <= 1;  //194 / 101 = 1
    16'b11000010_01100110 : OUT <= 1;  //194 / 102 = 1
    16'b11000010_01100111 : OUT <= 1;  //194 / 103 = 1
    16'b11000010_01101000 : OUT <= 1;  //194 / 104 = 1
    16'b11000010_01101001 : OUT <= 1;  //194 / 105 = 1
    16'b11000010_01101010 : OUT <= 1;  //194 / 106 = 1
    16'b11000010_01101011 : OUT <= 1;  //194 / 107 = 1
    16'b11000010_01101100 : OUT <= 1;  //194 / 108 = 1
    16'b11000010_01101101 : OUT <= 1;  //194 / 109 = 1
    16'b11000010_01101110 : OUT <= 1;  //194 / 110 = 1
    16'b11000010_01101111 : OUT <= 1;  //194 / 111 = 1
    16'b11000010_01110000 : OUT <= 1;  //194 / 112 = 1
    16'b11000010_01110001 : OUT <= 1;  //194 / 113 = 1
    16'b11000010_01110010 : OUT <= 1;  //194 / 114 = 1
    16'b11000010_01110011 : OUT <= 1;  //194 / 115 = 1
    16'b11000010_01110100 : OUT <= 1;  //194 / 116 = 1
    16'b11000010_01110101 : OUT <= 1;  //194 / 117 = 1
    16'b11000010_01110110 : OUT <= 1;  //194 / 118 = 1
    16'b11000010_01110111 : OUT <= 1;  //194 / 119 = 1
    16'b11000010_01111000 : OUT <= 1;  //194 / 120 = 1
    16'b11000010_01111001 : OUT <= 1;  //194 / 121 = 1
    16'b11000010_01111010 : OUT <= 1;  //194 / 122 = 1
    16'b11000010_01111011 : OUT <= 1;  //194 / 123 = 1
    16'b11000010_01111100 : OUT <= 1;  //194 / 124 = 1
    16'b11000010_01111101 : OUT <= 1;  //194 / 125 = 1
    16'b11000010_01111110 : OUT <= 1;  //194 / 126 = 1
    16'b11000010_01111111 : OUT <= 1;  //194 / 127 = 1
    16'b11000010_10000000 : OUT <= 1;  //194 / 128 = 1
    16'b11000010_10000001 : OUT <= 1;  //194 / 129 = 1
    16'b11000010_10000010 : OUT <= 1;  //194 / 130 = 1
    16'b11000010_10000011 : OUT <= 1;  //194 / 131 = 1
    16'b11000010_10000100 : OUT <= 1;  //194 / 132 = 1
    16'b11000010_10000101 : OUT <= 1;  //194 / 133 = 1
    16'b11000010_10000110 : OUT <= 1;  //194 / 134 = 1
    16'b11000010_10000111 : OUT <= 1;  //194 / 135 = 1
    16'b11000010_10001000 : OUT <= 1;  //194 / 136 = 1
    16'b11000010_10001001 : OUT <= 1;  //194 / 137 = 1
    16'b11000010_10001010 : OUT <= 1;  //194 / 138 = 1
    16'b11000010_10001011 : OUT <= 1;  //194 / 139 = 1
    16'b11000010_10001100 : OUT <= 1;  //194 / 140 = 1
    16'b11000010_10001101 : OUT <= 1;  //194 / 141 = 1
    16'b11000010_10001110 : OUT <= 1;  //194 / 142 = 1
    16'b11000010_10001111 : OUT <= 1;  //194 / 143 = 1
    16'b11000010_10010000 : OUT <= 1;  //194 / 144 = 1
    16'b11000010_10010001 : OUT <= 1;  //194 / 145 = 1
    16'b11000010_10010010 : OUT <= 1;  //194 / 146 = 1
    16'b11000010_10010011 : OUT <= 1;  //194 / 147 = 1
    16'b11000010_10010100 : OUT <= 1;  //194 / 148 = 1
    16'b11000010_10010101 : OUT <= 1;  //194 / 149 = 1
    16'b11000010_10010110 : OUT <= 1;  //194 / 150 = 1
    16'b11000010_10010111 : OUT <= 1;  //194 / 151 = 1
    16'b11000010_10011000 : OUT <= 1;  //194 / 152 = 1
    16'b11000010_10011001 : OUT <= 1;  //194 / 153 = 1
    16'b11000010_10011010 : OUT <= 1;  //194 / 154 = 1
    16'b11000010_10011011 : OUT <= 1;  //194 / 155 = 1
    16'b11000010_10011100 : OUT <= 1;  //194 / 156 = 1
    16'b11000010_10011101 : OUT <= 1;  //194 / 157 = 1
    16'b11000010_10011110 : OUT <= 1;  //194 / 158 = 1
    16'b11000010_10011111 : OUT <= 1;  //194 / 159 = 1
    16'b11000010_10100000 : OUT <= 1;  //194 / 160 = 1
    16'b11000010_10100001 : OUT <= 1;  //194 / 161 = 1
    16'b11000010_10100010 : OUT <= 1;  //194 / 162 = 1
    16'b11000010_10100011 : OUT <= 1;  //194 / 163 = 1
    16'b11000010_10100100 : OUT <= 1;  //194 / 164 = 1
    16'b11000010_10100101 : OUT <= 1;  //194 / 165 = 1
    16'b11000010_10100110 : OUT <= 1;  //194 / 166 = 1
    16'b11000010_10100111 : OUT <= 1;  //194 / 167 = 1
    16'b11000010_10101000 : OUT <= 1;  //194 / 168 = 1
    16'b11000010_10101001 : OUT <= 1;  //194 / 169 = 1
    16'b11000010_10101010 : OUT <= 1;  //194 / 170 = 1
    16'b11000010_10101011 : OUT <= 1;  //194 / 171 = 1
    16'b11000010_10101100 : OUT <= 1;  //194 / 172 = 1
    16'b11000010_10101101 : OUT <= 1;  //194 / 173 = 1
    16'b11000010_10101110 : OUT <= 1;  //194 / 174 = 1
    16'b11000010_10101111 : OUT <= 1;  //194 / 175 = 1
    16'b11000010_10110000 : OUT <= 1;  //194 / 176 = 1
    16'b11000010_10110001 : OUT <= 1;  //194 / 177 = 1
    16'b11000010_10110010 : OUT <= 1;  //194 / 178 = 1
    16'b11000010_10110011 : OUT <= 1;  //194 / 179 = 1
    16'b11000010_10110100 : OUT <= 1;  //194 / 180 = 1
    16'b11000010_10110101 : OUT <= 1;  //194 / 181 = 1
    16'b11000010_10110110 : OUT <= 1;  //194 / 182 = 1
    16'b11000010_10110111 : OUT <= 1;  //194 / 183 = 1
    16'b11000010_10111000 : OUT <= 1;  //194 / 184 = 1
    16'b11000010_10111001 : OUT <= 1;  //194 / 185 = 1
    16'b11000010_10111010 : OUT <= 1;  //194 / 186 = 1
    16'b11000010_10111011 : OUT <= 1;  //194 / 187 = 1
    16'b11000010_10111100 : OUT <= 1;  //194 / 188 = 1
    16'b11000010_10111101 : OUT <= 1;  //194 / 189 = 1
    16'b11000010_10111110 : OUT <= 1;  //194 / 190 = 1
    16'b11000010_10111111 : OUT <= 1;  //194 / 191 = 1
    16'b11000010_11000000 : OUT <= 1;  //194 / 192 = 1
    16'b11000010_11000001 : OUT <= 1;  //194 / 193 = 1
    16'b11000010_11000010 : OUT <= 1;  //194 / 194 = 1
    16'b11000010_11000011 : OUT <= 0;  //194 / 195 = 0
    16'b11000010_11000100 : OUT <= 0;  //194 / 196 = 0
    16'b11000010_11000101 : OUT <= 0;  //194 / 197 = 0
    16'b11000010_11000110 : OUT <= 0;  //194 / 198 = 0
    16'b11000010_11000111 : OUT <= 0;  //194 / 199 = 0
    16'b11000010_11001000 : OUT <= 0;  //194 / 200 = 0
    16'b11000010_11001001 : OUT <= 0;  //194 / 201 = 0
    16'b11000010_11001010 : OUT <= 0;  //194 / 202 = 0
    16'b11000010_11001011 : OUT <= 0;  //194 / 203 = 0
    16'b11000010_11001100 : OUT <= 0;  //194 / 204 = 0
    16'b11000010_11001101 : OUT <= 0;  //194 / 205 = 0
    16'b11000010_11001110 : OUT <= 0;  //194 / 206 = 0
    16'b11000010_11001111 : OUT <= 0;  //194 / 207 = 0
    16'b11000010_11010000 : OUT <= 0;  //194 / 208 = 0
    16'b11000010_11010001 : OUT <= 0;  //194 / 209 = 0
    16'b11000010_11010010 : OUT <= 0;  //194 / 210 = 0
    16'b11000010_11010011 : OUT <= 0;  //194 / 211 = 0
    16'b11000010_11010100 : OUT <= 0;  //194 / 212 = 0
    16'b11000010_11010101 : OUT <= 0;  //194 / 213 = 0
    16'b11000010_11010110 : OUT <= 0;  //194 / 214 = 0
    16'b11000010_11010111 : OUT <= 0;  //194 / 215 = 0
    16'b11000010_11011000 : OUT <= 0;  //194 / 216 = 0
    16'b11000010_11011001 : OUT <= 0;  //194 / 217 = 0
    16'b11000010_11011010 : OUT <= 0;  //194 / 218 = 0
    16'b11000010_11011011 : OUT <= 0;  //194 / 219 = 0
    16'b11000010_11011100 : OUT <= 0;  //194 / 220 = 0
    16'b11000010_11011101 : OUT <= 0;  //194 / 221 = 0
    16'b11000010_11011110 : OUT <= 0;  //194 / 222 = 0
    16'b11000010_11011111 : OUT <= 0;  //194 / 223 = 0
    16'b11000010_11100000 : OUT <= 0;  //194 / 224 = 0
    16'b11000010_11100001 : OUT <= 0;  //194 / 225 = 0
    16'b11000010_11100010 : OUT <= 0;  //194 / 226 = 0
    16'b11000010_11100011 : OUT <= 0;  //194 / 227 = 0
    16'b11000010_11100100 : OUT <= 0;  //194 / 228 = 0
    16'b11000010_11100101 : OUT <= 0;  //194 / 229 = 0
    16'b11000010_11100110 : OUT <= 0;  //194 / 230 = 0
    16'b11000010_11100111 : OUT <= 0;  //194 / 231 = 0
    16'b11000010_11101000 : OUT <= 0;  //194 / 232 = 0
    16'b11000010_11101001 : OUT <= 0;  //194 / 233 = 0
    16'b11000010_11101010 : OUT <= 0;  //194 / 234 = 0
    16'b11000010_11101011 : OUT <= 0;  //194 / 235 = 0
    16'b11000010_11101100 : OUT <= 0;  //194 / 236 = 0
    16'b11000010_11101101 : OUT <= 0;  //194 / 237 = 0
    16'b11000010_11101110 : OUT <= 0;  //194 / 238 = 0
    16'b11000010_11101111 : OUT <= 0;  //194 / 239 = 0
    16'b11000010_11110000 : OUT <= 0;  //194 / 240 = 0
    16'b11000010_11110001 : OUT <= 0;  //194 / 241 = 0
    16'b11000010_11110010 : OUT <= 0;  //194 / 242 = 0
    16'b11000010_11110011 : OUT <= 0;  //194 / 243 = 0
    16'b11000010_11110100 : OUT <= 0;  //194 / 244 = 0
    16'b11000010_11110101 : OUT <= 0;  //194 / 245 = 0
    16'b11000010_11110110 : OUT <= 0;  //194 / 246 = 0
    16'b11000010_11110111 : OUT <= 0;  //194 / 247 = 0
    16'b11000010_11111000 : OUT <= 0;  //194 / 248 = 0
    16'b11000010_11111001 : OUT <= 0;  //194 / 249 = 0
    16'b11000010_11111010 : OUT <= 0;  //194 / 250 = 0
    16'b11000010_11111011 : OUT <= 0;  //194 / 251 = 0
    16'b11000010_11111100 : OUT <= 0;  //194 / 252 = 0
    16'b11000010_11111101 : OUT <= 0;  //194 / 253 = 0
    16'b11000010_11111110 : OUT <= 0;  //194 / 254 = 0
    16'b11000010_11111111 : OUT <= 0;  //194 / 255 = 0
    16'b11000011_00000000 : OUT <= 0;  //195 / 0 = 0
    16'b11000011_00000001 : OUT <= 195;  //195 / 1 = 195
    16'b11000011_00000010 : OUT <= 97;  //195 / 2 = 97
    16'b11000011_00000011 : OUT <= 65;  //195 / 3 = 65
    16'b11000011_00000100 : OUT <= 48;  //195 / 4 = 48
    16'b11000011_00000101 : OUT <= 39;  //195 / 5 = 39
    16'b11000011_00000110 : OUT <= 32;  //195 / 6 = 32
    16'b11000011_00000111 : OUT <= 27;  //195 / 7 = 27
    16'b11000011_00001000 : OUT <= 24;  //195 / 8 = 24
    16'b11000011_00001001 : OUT <= 21;  //195 / 9 = 21
    16'b11000011_00001010 : OUT <= 19;  //195 / 10 = 19
    16'b11000011_00001011 : OUT <= 17;  //195 / 11 = 17
    16'b11000011_00001100 : OUT <= 16;  //195 / 12 = 16
    16'b11000011_00001101 : OUT <= 15;  //195 / 13 = 15
    16'b11000011_00001110 : OUT <= 13;  //195 / 14 = 13
    16'b11000011_00001111 : OUT <= 13;  //195 / 15 = 13
    16'b11000011_00010000 : OUT <= 12;  //195 / 16 = 12
    16'b11000011_00010001 : OUT <= 11;  //195 / 17 = 11
    16'b11000011_00010010 : OUT <= 10;  //195 / 18 = 10
    16'b11000011_00010011 : OUT <= 10;  //195 / 19 = 10
    16'b11000011_00010100 : OUT <= 9;  //195 / 20 = 9
    16'b11000011_00010101 : OUT <= 9;  //195 / 21 = 9
    16'b11000011_00010110 : OUT <= 8;  //195 / 22 = 8
    16'b11000011_00010111 : OUT <= 8;  //195 / 23 = 8
    16'b11000011_00011000 : OUT <= 8;  //195 / 24 = 8
    16'b11000011_00011001 : OUT <= 7;  //195 / 25 = 7
    16'b11000011_00011010 : OUT <= 7;  //195 / 26 = 7
    16'b11000011_00011011 : OUT <= 7;  //195 / 27 = 7
    16'b11000011_00011100 : OUT <= 6;  //195 / 28 = 6
    16'b11000011_00011101 : OUT <= 6;  //195 / 29 = 6
    16'b11000011_00011110 : OUT <= 6;  //195 / 30 = 6
    16'b11000011_00011111 : OUT <= 6;  //195 / 31 = 6
    16'b11000011_00100000 : OUT <= 6;  //195 / 32 = 6
    16'b11000011_00100001 : OUT <= 5;  //195 / 33 = 5
    16'b11000011_00100010 : OUT <= 5;  //195 / 34 = 5
    16'b11000011_00100011 : OUT <= 5;  //195 / 35 = 5
    16'b11000011_00100100 : OUT <= 5;  //195 / 36 = 5
    16'b11000011_00100101 : OUT <= 5;  //195 / 37 = 5
    16'b11000011_00100110 : OUT <= 5;  //195 / 38 = 5
    16'b11000011_00100111 : OUT <= 5;  //195 / 39 = 5
    16'b11000011_00101000 : OUT <= 4;  //195 / 40 = 4
    16'b11000011_00101001 : OUT <= 4;  //195 / 41 = 4
    16'b11000011_00101010 : OUT <= 4;  //195 / 42 = 4
    16'b11000011_00101011 : OUT <= 4;  //195 / 43 = 4
    16'b11000011_00101100 : OUT <= 4;  //195 / 44 = 4
    16'b11000011_00101101 : OUT <= 4;  //195 / 45 = 4
    16'b11000011_00101110 : OUT <= 4;  //195 / 46 = 4
    16'b11000011_00101111 : OUT <= 4;  //195 / 47 = 4
    16'b11000011_00110000 : OUT <= 4;  //195 / 48 = 4
    16'b11000011_00110001 : OUT <= 3;  //195 / 49 = 3
    16'b11000011_00110010 : OUT <= 3;  //195 / 50 = 3
    16'b11000011_00110011 : OUT <= 3;  //195 / 51 = 3
    16'b11000011_00110100 : OUT <= 3;  //195 / 52 = 3
    16'b11000011_00110101 : OUT <= 3;  //195 / 53 = 3
    16'b11000011_00110110 : OUT <= 3;  //195 / 54 = 3
    16'b11000011_00110111 : OUT <= 3;  //195 / 55 = 3
    16'b11000011_00111000 : OUT <= 3;  //195 / 56 = 3
    16'b11000011_00111001 : OUT <= 3;  //195 / 57 = 3
    16'b11000011_00111010 : OUT <= 3;  //195 / 58 = 3
    16'b11000011_00111011 : OUT <= 3;  //195 / 59 = 3
    16'b11000011_00111100 : OUT <= 3;  //195 / 60 = 3
    16'b11000011_00111101 : OUT <= 3;  //195 / 61 = 3
    16'b11000011_00111110 : OUT <= 3;  //195 / 62 = 3
    16'b11000011_00111111 : OUT <= 3;  //195 / 63 = 3
    16'b11000011_01000000 : OUT <= 3;  //195 / 64 = 3
    16'b11000011_01000001 : OUT <= 3;  //195 / 65 = 3
    16'b11000011_01000010 : OUT <= 2;  //195 / 66 = 2
    16'b11000011_01000011 : OUT <= 2;  //195 / 67 = 2
    16'b11000011_01000100 : OUT <= 2;  //195 / 68 = 2
    16'b11000011_01000101 : OUT <= 2;  //195 / 69 = 2
    16'b11000011_01000110 : OUT <= 2;  //195 / 70 = 2
    16'b11000011_01000111 : OUT <= 2;  //195 / 71 = 2
    16'b11000011_01001000 : OUT <= 2;  //195 / 72 = 2
    16'b11000011_01001001 : OUT <= 2;  //195 / 73 = 2
    16'b11000011_01001010 : OUT <= 2;  //195 / 74 = 2
    16'b11000011_01001011 : OUT <= 2;  //195 / 75 = 2
    16'b11000011_01001100 : OUT <= 2;  //195 / 76 = 2
    16'b11000011_01001101 : OUT <= 2;  //195 / 77 = 2
    16'b11000011_01001110 : OUT <= 2;  //195 / 78 = 2
    16'b11000011_01001111 : OUT <= 2;  //195 / 79 = 2
    16'b11000011_01010000 : OUT <= 2;  //195 / 80 = 2
    16'b11000011_01010001 : OUT <= 2;  //195 / 81 = 2
    16'b11000011_01010010 : OUT <= 2;  //195 / 82 = 2
    16'b11000011_01010011 : OUT <= 2;  //195 / 83 = 2
    16'b11000011_01010100 : OUT <= 2;  //195 / 84 = 2
    16'b11000011_01010101 : OUT <= 2;  //195 / 85 = 2
    16'b11000011_01010110 : OUT <= 2;  //195 / 86 = 2
    16'b11000011_01010111 : OUT <= 2;  //195 / 87 = 2
    16'b11000011_01011000 : OUT <= 2;  //195 / 88 = 2
    16'b11000011_01011001 : OUT <= 2;  //195 / 89 = 2
    16'b11000011_01011010 : OUT <= 2;  //195 / 90 = 2
    16'b11000011_01011011 : OUT <= 2;  //195 / 91 = 2
    16'b11000011_01011100 : OUT <= 2;  //195 / 92 = 2
    16'b11000011_01011101 : OUT <= 2;  //195 / 93 = 2
    16'b11000011_01011110 : OUT <= 2;  //195 / 94 = 2
    16'b11000011_01011111 : OUT <= 2;  //195 / 95 = 2
    16'b11000011_01100000 : OUT <= 2;  //195 / 96 = 2
    16'b11000011_01100001 : OUT <= 2;  //195 / 97 = 2
    16'b11000011_01100010 : OUT <= 1;  //195 / 98 = 1
    16'b11000011_01100011 : OUT <= 1;  //195 / 99 = 1
    16'b11000011_01100100 : OUT <= 1;  //195 / 100 = 1
    16'b11000011_01100101 : OUT <= 1;  //195 / 101 = 1
    16'b11000011_01100110 : OUT <= 1;  //195 / 102 = 1
    16'b11000011_01100111 : OUT <= 1;  //195 / 103 = 1
    16'b11000011_01101000 : OUT <= 1;  //195 / 104 = 1
    16'b11000011_01101001 : OUT <= 1;  //195 / 105 = 1
    16'b11000011_01101010 : OUT <= 1;  //195 / 106 = 1
    16'b11000011_01101011 : OUT <= 1;  //195 / 107 = 1
    16'b11000011_01101100 : OUT <= 1;  //195 / 108 = 1
    16'b11000011_01101101 : OUT <= 1;  //195 / 109 = 1
    16'b11000011_01101110 : OUT <= 1;  //195 / 110 = 1
    16'b11000011_01101111 : OUT <= 1;  //195 / 111 = 1
    16'b11000011_01110000 : OUT <= 1;  //195 / 112 = 1
    16'b11000011_01110001 : OUT <= 1;  //195 / 113 = 1
    16'b11000011_01110010 : OUT <= 1;  //195 / 114 = 1
    16'b11000011_01110011 : OUT <= 1;  //195 / 115 = 1
    16'b11000011_01110100 : OUT <= 1;  //195 / 116 = 1
    16'b11000011_01110101 : OUT <= 1;  //195 / 117 = 1
    16'b11000011_01110110 : OUT <= 1;  //195 / 118 = 1
    16'b11000011_01110111 : OUT <= 1;  //195 / 119 = 1
    16'b11000011_01111000 : OUT <= 1;  //195 / 120 = 1
    16'b11000011_01111001 : OUT <= 1;  //195 / 121 = 1
    16'b11000011_01111010 : OUT <= 1;  //195 / 122 = 1
    16'b11000011_01111011 : OUT <= 1;  //195 / 123 = 1
    16'b11000011_01111100 : OUT <= 1;  //195 / 124 = 1
    16'b11000011_01111101 : OUT <= 1;  //195 / 125 = 1
    16'b11000011_01111110 : OUT <= 1;  //195 / 126 = 1
    16'b11000011_01111111 : OUT <= 1;  //195 / 127 = 1
    16'b11000011_10000000 : OUT <= 1;  //195 / 128 = 1
    16'b11000011_10000001 : OUT <= 1;  //195 / 129 = 1
    16'b11000011_10000010 : OUT <= 1;  //195 / 130 = 1
    16'b11000011_10000011 : OUT <= 1;  //195 / 131 = 1
    16'b11000011_10000100 : OUT <= 1;  //195 / 132 = 1
    16'b11000011_10000101 : OUT <= 1;  //195 / 133 = 1
    16'b11000011_10000110 : OUT <= 1;  //195 / 134 = 1
    16'b11000011_10000111 : OUT <= 1;  //195 / 135 = 1
    16'b11000011_10001000 : OUT <= 1;  //195 / 136 = 1
    16'b11000011_10001001 : OUT <= 1;  //195 / 137 = 1
    16'b11000011_10001010 : OUT <= 1;  //195 / 138 = 1
    16'b11000011_10001011 : OUT <= 1;  //195 / 139 = 1
    16'b11000011_10001100 : OUT <= 1;  //195 / 140 = 1
    16'b11000011_10001101 : OUT <= 1;  //195 / 141 = 1
    16'b11000011_10001110 : OUT <= 1;  //195 / 142 = 1
    16'b11000011_10001111 : OUT <= 1;  //195 / 143 = 1
    16'b11000011_10010000 : OUT <= 1;  //195 / 144 = 1
    16'b11000011_10010001 : OUT <= 1;  //195 / 145 = 1
    16'b11000011_10010010 : OUT <= 1;  //195 / 146 = 1
    16'b11000011_10010011 : OUT <= 1;  //195 / 147 = 1
    16'b11000011_10010100 : OUT <= 1;  //195 / 148 = 1
    16'b11000011_10010101 : OUT <= 1;  //195 / 149 = 1
    16'b11000011_10010110 : OUT <= 1;  //195 / 150 = 1
    16'b11000011_10010111 : OUT <= 1;  //195 / 151 = 1
    16'b11000011_10011000 : OUT <= 1;  //195 / 152 = 1
    16'b11000011_10011001 : OUT <= 1;  //195 / 153 = 1
    16'b11000011_10011010 : OUT <= 1;  //195 / 154 = 1
    16'b11000011_10011011 : OUT <= 1;  //195 / 155 = 1
    16'b11000011_10011100 : OUT <= 1;  //195 / 156 = 1
    16'b11000011_10011101 : OUT <= 1;  //195 / 157 = 1
    16'b11000011_10011110 : OUT <= 1;  //195 / 158 = 1
    16'b11000011_10011111 : OUT <= 1;  //195 / 159 = 1
    16'b11000011_10100000 : OUT <= 1;  //195 / 160 = 1
    16'b11000011_10100001 : OUT <= 1;  //195 / 161 = 1
    16'b11000011_10100010 : OUT <= 1;  //195 / 162 = 1
    16'b11000011_10100011 : OUT <= 1;  //195 / 163 = 1
    16'b11000011_10100100 : OUT <= 1;  //195 / 164 = 1
    16'b11000011_10100101 : OUT <= 1;  //195 / 165 = 1
    16'b11000011_10100110 : OUT <= 1;  //195 / 166 = 1
    16'b11000011_10100111 : OUT <= 1;  //195 / 167 = 1
    16'b11000011_10101000 : OUT <= 1;  //195 / 168 = 1
    16'b11000011_10101001 : OUT <= 1;  //195 / 169 = 1
    16'b11000011_10101010 : OUT <= 1;  //195 / 170 = 1
    16'b11000011_10101011 : OUT <= 1;  //195 / 171 = 1
    16'b11000011_10101100 : OUT <= 1;  //195 / 172 = 1
    16'b11000011_10101101 : OUT <= 1;  //195 / 173 = 1
    16'b11000011_10101110 : OUT <= 1;  //195 / 174 = 1
    16'b11000011_10101111 : OUT <= 1;  //195 / 175 = 1
    16'b11000011_10110000 : OUT <= 1;  //195 / 176 = 1
    16'b11000011_10110001 : OUT <= 1;  //195 / 177 = 1
    16'b11000011_10110010 : OUT <= 1;  //195 / 178 = 1
    16'b11000011_10110011 : OUT <= 1;  //195 / 179 = 1
    16'b11000011_10110100 : OUT <= 1;  //195 / 180 = 1
    16'b11000011_10110101 : OUT <= 1;  //195 / 181 = 1
    16'b11000011_10110110 : OUT <= 1;  //195 / 182 = 1
    16'b11000011_10110111 : OUT <= 1;  //195 / 183 = 1
    16'b11000011_10111000 : OUT <= 1;  //195 / 184 = 1
    16'b11000011_10111001 : OUT <= 1;  //195 / 185 = 1
    16'b11000011_10111010 : OUT <= 1;  //195 / 186 = 1
    16'b11000011_10111011 : OUT <= 1;  //195 / 187 = 1
    16'b11000011_10111100 : OUT <= 1;  //195 / 188 = 1
    16'b11000011_10111101 : OUT <= 1;  //195 / 189 = 1
    16'b11000011_10111110 : OUT <= 1;  //195 / 190 = 1
    16'b11000011_10111111 : OUT <= 1;  //195 / 191 = 1
    16'b11000011_11000000 : OUT <= 1;  //195 / 192 = 1
    16'b11000011_11000001 : OUT <= 1;  //195 / 193 = 1
    16'b11000011_11000010 : OUT <= 1;  //195 / 194 = 1
    16'b11000011_11000011 : OUT <= 1;  //195 / 195 = 1
    16'b11000011_11000100 : OUT <= 0;  //195 / 196 = 0
    16'b11000011_11000101 : OUT <= 0;  //195 / 197 = 0
    16'b11000011_11000110 : OUT <= 0;  //195 / 198 = 0
    16'b11000011_11000111 : OUT <= 0;  //195 / 199 = 0
    16'b11000011_11001000 : OUT <= 0;  //195 / 200 = 0
    16'b11000011_11001001 : OUT <= 0;  //195 / 201 = 0
    16'b11000011_11001010 : OUT <= 0;  //195 / 202 = 0
    16'b11000011_11001011 : OUT <= 0;  //195 / 203 = 0
    16'b11000011_11001100 : OUT <= 0;  //195 / 204 = 0
    16'b11000011_11001101 : OUT <= 0;  //195 / 205 = 0
    16'b11000011_11001110 : OUT <= 0;  //195 / 206 = 0
    16'b11000011_11001111 : OUT <= 0;  //195 / 207 = 0
    16'b11000011_11010000 : OUT <= 0;  //195 / 208 = 0
    16'b11000011_11010001 : OUT <= 0;  //195 / 209 = 0
    16'b11000011_11010010 : OUT <= 0;  //195 / 210 = 0
    16'b11000011_11010011 : OUT <= 0;  //195 / 211 = 0
    16'b11000011_11010100 : OUT <= 0;  //195 / 212 = 0
    16'b11000011_11010101 : OUT <= 0;  //195 / 213 = 0
    16'b11000011_11010110 : OUT <= 0;  //195 / 214 = 0
    16'b11000011_11010111 : OUT <= 0;  //195 / 215 = 0
    16'b11000011_11011000 : OUT <= 0;  //195 / 216 = 0
    16'b11000011_11011001 : OUT <= 0;  //195 / 217 = 0
    16'b11000011_11011010 : OUT <= 0;  //195 / 218 = 0
    16'b11000011_11011011 : OUT <= 0;  //195 / 219 = 0
    16'b11000011_11011100 : OUT <= 0;  //195 / 220 = 0
    16'b11000011_11011101 : OUT <= 0;  //195 / 221 = 0
    16'b11000011_11011110 : OUT <= 0;  //195 / 222 = 0
    16'b11000011_11011111 : OUT <= 0;  //195 / 223 = 0
    16'b11000011_11100000 : OUT <= 0;  //195 / 224 = 0
    16'b11000011_11100001 : OUT <= 0;  //195 / 225 = 0
    16'b11000011_11100010 : OUT <= 0;  //195 / 226 = 0
    16'b11000011_11100011 : OUT <= 0;  //195 / 227 = 0
    16'b11000011_11100100 : OUT <= 0;  //195 / 228 = 0
    16'b11000011_11100101 : OUT <= 0;  //195 / 229 = 0
    16'b11000011_11100110 : OUT <= 0;  //195 / 230 = 0
    16'b11000011_11100111 : OUT <= 0;  //195 / 231 = 0
    16'b11000011_11101000 : OUT <= 0;  //195 / 232 = 0
    16'b11000011_11101001 : OUT <= 0;  //195 / 233 = 0
    16'b11000011_11101010 : OUT <= 0;  //195 / 234 = 0
    16'b11000011_11101011 : OUT <= 0;  //195 / 235 = 0
    16'b11000011_11101100 : OUT <= 0;  //195 / 236 = 0
    16'b11000011_11101101 : OUT <= 0;  //195 / 237 = 0
    16'b11000011_11101110 : OUT <= 0;  //195 / 238 = 0
    16'b11000011_11101111 : OUT <= 0;  //195 / 239 = 0
    16'b11000011_11110000 : OUT <= 0;  //195 / 240 = 0
    16'b11000011_11110001 : OUT <= 0;  //195 / 241 = 0
    16'b11000011_11110010 : OUT <= 0;  //195 / 242 = 0
    16'b11000011_11110011 : OUT <= 0;  //195 / 243 = 0
    16'b11000011_11110100 : OUT <= 0;  //195 / 244 = 0
    16'b11000011_11110101 : OUT <= 0;  //195 / 245 = 0
    16'b11000011_11110110 : OUT <= 0;  //195 / 246 = 0
    16'b11000011_11110111 : OUT <= 0;  //195 / 247 = 0
    16'b11000011_11111000 : OUT <= 0;  //195 / 248 = 0
    16'b11000011_11111001 : OUT <= 0;  //195 / 249 = 0
    16'b11000011_11111010 : OUT <= 0;  //195 / 250 = 0
    16'b11000011_11111011 : OUT <= 0;  //195 / 251 = 0
    16'b11000011_11111100 : OUT <= 0;  //195 / 252 = 0
    16'b11000011_11111101 : OUT <= 0;  //195 / 253 = 0
    16'b11000011_11111110 : OUT <= 0;  //195 / 254 = 0
    16'b11000011_11111111 : OUT <= 0;  //195 / 255 = 0
    16'b11000100_00000000 : OUT <= 0;  //196 / 0 = 0
    16'b11000100_00000001 : OUT <= 196;  //196 / 1 = 196
    16'b11000100_00000010 : OUT <= 98;  //196 / 2 = 98
    16'b11000100_00000011 : OUT <= 65;  //196 / 3 = 65
    16'b11000100_00000100 : OUT <= 49;  //196 / 4 = 49
    16'b11000100_00000101 : OUT <= 39;  //196 / 5 = 39
    16'b11000100_00000110 : OUT <= 32;  //196 / 6 = 32
    16'b11000100_00000111 : OUT <= 28;  //196 / 7 = 28
    16'b11000100_00001000 : OUT <= 24;  //196 / 8 = 24
    16'b11000100_00001001 : OUT <= 21;  //196 / 9 = 21
    16'b11000100_00001010 : OUT <= 19;  //196 / 10 = 19
    16'b11000100_00001011 : OUT <= 17;  //196 / 11 = 17
    16'b11000100_00001100 : OUT <= 16;  //196 / 12 = 16
    16'b11000100_00001101 : OUT <= 15;  //196 / 13 = 15
    16'b11000100_00001110 : OUT <= 14;  //196 / 14 = 14
    16'b11000100_00001111 : OUT <= 13;  //196 / 15 = 13
    16'b11000100_00010000 : OUT <= 12;  //196 / 16 = 12
    16'b11000100_00010001 : OUT <= 11;  //196 / 17 = 11
    16'b11000100_00010010 : OUT <= 10;  //196 / 18 = 10
    16'b11000100_00010011 : OUT <= 10;  //196 / 19 = 10
    16'b11000100_00010100 : OUT <= 9;  //196 / 20 = 9
    16'b11000100_00010101 : OUT <= 9;  //196 / 21 = 9
    16'b11000100_00010110 : OUT <= 8;  //196 / 22 = 8
    16'b11000100_00010111 : OUT <= 8;  //196 / 23 = 8
    16'b11000100_00011000 : OUT <= 8;  //196 / 24 = 8
    16'b11000100_00011001 : OUT <= 7;  //196 / 25 = 7
    16'b11000100_00011010 : OUT <= 7;  //196 / 26 = 7
    16'b11000100_00011011 : OUT <= 7;  //196 / 27 = 7
    16'b11000100_00011100 : OUT <= 7;  //196 / 28 = 7
    16'b11000100_00011101 : OUT <= 6;  //196 / 29 = 6
    16'b11000100_00011110 : OUT <= 6;  //196 / 30 = 6
    16'b11000100_00011111 : OUT <= 6;  //196 / 31 = 6
    16'b11000100_00100000 : OUT <= 6;  //196 / 32 = 6
    16'b11000100_00100001 : OUT <= 5;  //196 / 33 = 5
    16'b11000100_00100010 : OUT <= 5;  //196 / 34 = 5
    16'b11000100_00100011 : OUT <= 5;  //196 / 35 = 5
    16'b11000100_00100100 : OUT <= 5;  //196 / 36 = 5
    16'b11000100_00100101 : OUT <= 5;  //196 / 37 = 5
    16'b11000100_00100110 : OUT <= 5;  //196 / 38 = 5
    16'b11000100_00100111 : OUT <= 5;  //196 / 39 = 5
    16'b11000100_00101000 : OUT <= 4;  //196 / 40 = 4
    16'b11000100_00101001 : OUT <= 4;  //196 / 41 = 4
    16'b11000100_00101010 : OUT <= 4;  //196 / 42 = 4
    16'b11000100_00101011 : OUT <= 4;  //196 / 43 = 4
    16'b11000100_00101100 : OUT <= 4;  //196 / 44 = 4
    16'b11000100_00101101 : OUT <= 4;  //196 / 45 = 4
    16'b11000100_00101110 : OUT <= 4;  //196 / 46 = 4
    16'b11000100_00101111 : OUT <= 4;  //196 / 47 = 4
    16'b11000100_00110000 : OUT <= 4;  //196 / 48 = 4
    16'b11000100_00110001 : OUT <= 4;  //196 / 49 = 4
    16'b11000100_00110010 : OUT <= 3;  //196 / 50 = 3
    16'b11000100_00110011 : OUT <= 3;  //196 / 51 = 3
    16'b11000100_00110100 : OUT <= 3;  //196 / 52 = 3
    16'b11000100_00110101 : OUT <= 3;  //196 / 53 = 3
    16'b11000100_00110110 : OUT <= 3;  //196 / 54 = 3
    16'b11000100_00110111 : OUT <= 3;  //196 / 55 = 3
    16'b11000100_00111000 : OUT <= 3;  //196 / 56 = 3
    16'b11000100_00111001 : OUT <= 3;  //196 / 57 = 3
    16'b11000100_00111010 : OUT <= 3;  //196 / 58 = 3
    16'b11000100_00111011 : OUT <= 3;  //196 / 59 = 3
    16'b11000100_00111100 : OUT <= 3;  //196 / 60 = 3
    16'b11000100_00111101 : OUT <= 3;  //196 / 61 = 3
    16'b11000100_00111110 : OUT <= 3;  //196 / 62 = 3
    16'b11000100_00111111 : OUT <= 3;  //196 / 63 = 3
    16'b11000100_01000000 : OUT <= 3;  //196 / 64 = 3
    16'b11000100_01000001 : OUT <= 3;  //196 / 65 = 3
    16'b11000100_01000010 : OUT <= 2;  //196 / 66 = 2
    16'b11000100_01000011 : OUT <= 2;  //196 / 67 = 2
    16'b11000100_01000100 : OUT <= 2;  //196 / 68 = 2
    16'b11000100_01000101 : OUT <= 2;  //196 / 69 = 2
    16'b11000100_01000110 : OUT <= 2;  //196 / 70 = 2
    16'b11000100_01000111 : OUT <= 2;  //196 / 71 = 2
    16'b11000100_01001000 : OUT <= 2;  //196 / 72 = 2
    16'b11000100_01001001 : OUT <= 2;  //196 / 73 = 2
    16'b11000100_01001010 : OUT <= 2;  //196 / 74 = 2
    16'b11000100_01001011 : OUT <= 2;  //196 / 75 = 2
    16'b11000100_01001100 : OUT <= 2;  //196 / 76 = 2
    16'b11000100_01001101 : OUT <= 2;  //196 / 77 = 2
    16'b11000100_01001110 : OUT <= 2;  //196 / 78 = 2
    16'b11000100_01001111 : OUT <= 2;  //196 / 79 = 2
    16'b11000100_01010000 : OUT <= 2;  //196 / 80 = 2
    16'b11000100_01010001 : OUT <= 2;  //196 / 81 = 2
    16'b11000100_01010010 : OUT <= 2;  //196 / 82 = 2
    16'b11000100_01010011 : OUT <= 2;  //196 / 83 = 2
    16'b11000100_01010100 : OUT <= 2;  //196 / 84 = 2
    16'b11000100_01010101 : OUT <= 2;  //196 / 85 = 2
    16'b11000100_01010110 : OUT <= 2;  //196 / 86 = 2
    16'b11000100_01010111 : OUT <= 2;  //196 / 87 = 2
    16'b11000100_01011000 : OUT <= 2;  //196 / 88 = 2
    16'b11000100_01011001 : OUT <= 2;  //196 / 89 = 2
    16'b11000100_01011010 : OUT <= 2;  //196 / 90 = 2
    16'b11000100_01011011 : OUT <= 2;  //196 / 91 = 2
    16'b11000100_01011100 : OUT <= 2;  //196 / 92 = 2
    16'b11000100_01011101 : OUT <= 2;  //196 / 93 = 2
    16'b11000100_01011110 : OUT <= 2;  //196 / 94 = 2
    16'b11000100_01011111 : OUT <= 2;  //196 / 95 = 2
    16'b11000100_01100000 : OUT <= 2;  //196 / 96 = 2
    16'b11000100_01100001 : OUT <= 2;  //196 / 97 = 2
    16'b11000100_01100010 : OUT <= 2;  //196 / 98 = 2
    16'b11000100_01100011 : OUT <= 1;  //196 / 99 = 1
    16'b11000100_01100100 : OUT <= 1;  //196 / 100 = 1
    16'b11000100_01100101 : OUT <= 1;  //196 / 101 = 1
    16'b11000100_01100110 : OUT <= 1;  //196 / 102 = 1
    16'b11000100_01100111 : OUT <= 1;  //196 / 103 = 1
    16'b11000100_01101000 : OUT <= 1;  //196 / 104 = 1
    16'b11000100_01101001 : OUT <= 1;  //196 / 105 = 1
    16'b11000100_01101010 : OUT <= 1;  //196 / 106 = 1
    16'b11000100_01101011 : OUT <= 1;  //196 / 107 = 1
    16'b11000100_01101100 : OUT <= 1;  //196 / 108 = 1
    16'b11000100_01101101 : OUT <= 1;  //196 / 109 = 1
    16'b11000100_01101110 : OUT <= 1;  //196 / 110 = 1
    16'b11000100_01101111 : OUT <= 1;  //196 / 111 = 1
    16'b11000100_01110000 : OUT <= 1;  //196 / 112 = 1
    16'b11000100_01110001 : OUT <= 1;  //196 / 113 = 1
    16'b11000100_01110010 : OUT <= 1;  //196 / 114 = 1
    16'b11000100_01110011 : OUT <= 1;  //196 / 115 = 1
    16'b11000100_01110100 : OUT <= 1;  //196 / 116 = 1
    16'b11000100_01110101 : OUT <= 1;  //196 / 117 = 1
    16'b11000100_01110110 : OUT <= 1;  //196 / 118 = 1
    16'b11000100_01110111 : OUT <= 1;  //196 / 119 = 1
    16'b11000100_01111000 : OUT <= 1;  //196 / 120 = 1
    16'b11000100_01111001 : OUT <= 1;  //196 / 121 = 1
    16'b11000100_01111010 : OUT <= 1;  //196 / 122 = 1
    16'b11000100_01111011 : OUT <= 1;  //196 / 123 = 1
    16'b11000100_01111100 : OUT <= 1;  //196 / 124 = 1
    16'b11000100_01111101 : OUT <= 1;  //196 / 125 = 1
    16'b11000100_01111110 : OUT <= 1;  //196 / 126 = 1
    16'b11000100_01111111 : OUT <= 1;  //196 / 127 = 1
    16'b11000100_10000000 : OUT <= 1;  //196 / 128 = 1
    16'b11000100_10000001 : OUT <= 1;  //196 / 129 = 1
    16'b11000100_10000010 : OUT <= 1;  //196 / 130 = 1
    16'b11000100_10000011 : OUT <= 1;  //196 / 131 = 1
    16'b11000100_10000100 : OUT <= 1;  //196 / 132 = 1
    16'b11000100_10000101 : OUT <= 1;  //196 / 133 = 1
    16'b11000100_10000110 : OUT <= 1;  //196 / 134 = 1
    16'b11000100_10000111 : OUT <= 1;  //196 / 135 = 1
    16'b11000100_10001000 : OUT <= 1;  //196 / 136 = 1
    16'b11000100_10001001 : OUT <= 1;  //196 / 137 = 1
    16'b11000100_10001010 : OUT <= 1;  //196 / 138 = 1
    16'b11000100_10001011 : OUT <= 1;  //196 / 139 = 1
    16'b11000100_10001100 : OUT <= 1;  //196 / 140 = 1
    16'b11000100_10001101 : OUT <= 1;  //196 / 141 = 1
    16'b11000100_10001110 : OUT <= 1;  //196 / 142 = 1
    16'b11000100_10001111 : OUT <= 1;  //196 / 143 = 1
    16'b11000100_10010000 : OUT <= 1;  //196 / 144 = 1
    16'b11000100_10010001 : OUT <= 1;  //196 / 145 = 1
    16'b11000100_10010010 : OUT <= 1;  //196 / 146 = 1
    16'b11000100_10010011 : OUT <= 1;  //196 / 147 = 1
    16'b11000100_10010100 : OUT <= 1;  //196 / 148 = 1
    16'b11000100_10010101 : OUT <= 1;  //196 / 149 = 1
    16'b11000100_10010110 : OUT <= 1;  //196 / 150 = 1
    16'b11000100_10010111 : OUT <= 1;  //196 / 151 = 1
    16'b11000100_10011000 : OUT <= 1;  //196 / 152 = 1
    16'b11000100_10011001 : OUT <= 1;  //196 / 153 = 1
    16'b11000100_10011010 : OUT <= 1;  //196 / 154 = 1
    16'b11000100_10011011 : OUT <= 1;  //196 / 155 = 1
    16'b11000100_10011100 : OUT <= 1;  //196 / 156 = 1
    16'b11000100_10011101 : OUT <= 1;  //196 / 157 = 1
    16'b11000100_10011110 : OUT <= 1;  //196 / 158 = 1
    16'b11000100_10011111 : OUT <= 1;  //196 / 159 = 1
    16'b11000100_10100000 : OUT <= 1;  //196 / 160 = 1
    16'b11000100_10100001 : OUT <= 1;  //196 / 161 = 1
    16'b11000100_10100010 : OUT <= 1;  //196 / 162 = 1
    16'b11000100_10100011 : OUT <= 1;  //196 / 163 = 1
    16'b11000100_10100100 : OUT <= 1;  //196 / 164 = 1
    16'b11000100_10100101 : OUT <= 1;  //196 / 165 = 1
    16'b11000100_10100110 : OUT <= 1;  //196 / 166 = 1
    16'b11000100_10100111 : OUT <= 1;  //196 / 167 = 1
    16'b11000100_10101000 : OUT <= 1;  //196 / 168 = 1
    16'b11000100_10101001 : OUT <= 1;  //196 / 169 = 1
    16'b11000100_10101010 : OUT <= 1;  //196 / 170 = 1
    16'b11000100_10101011 : OUT <= 1;  //196 / 171 = 1
    16'b11000100_10101100 : OUT <= 1;  //196 / 172 = 1
    16'b11000100_10101101 : OUT <= 1;  //196 / 173 = 1
    16'b11000100_10101110 : OUT <= 1;  //196 / 174 = 1
    16'b11000100_10101111 : OUT <= 1;  //196 / 175 = 1
    16'b11000100_10110000 : OUT <= 1;  //196 / 176 = 1
    16'b11000100_10110001 : OUT <= 1;  //196 / 177 = 1
    16'b11000100_10110010 : OUT <= 1;  //196 / 178 = 1
    16'b11000100_10110011 : OUT <= 1;  //196 / 179 = 1
    16'b11000100_10110100 : OUT <= 1;  //196 / 180 = 1
    16'b11000100_10110101 : OUT <= 1;  //196 / 181 = 1
    16'b11000100_10110110 : OUT <= 1;  //196 / 182 = 1
    16'b11000100_10110111 : OUT <= 1;  //196 / 183 = 1
    16'b11000100_10111000 : OUT <= 1;  //196 / 184 = 1
    16'b11000100_10111001 : OUT <= 1;  //196 / 185 = 1
    16'b11000100_10111010 : OUT <= 1;  //196 / 186 = 1
    16'b11000100_10111011 : OUT <= 1;  //196 / 187 = 1
    16'b11000100_10111100 : OUT <= 1;  //196 / 188 = 1
    16'b11000100_10111101 : OUT <= 1;  //196 / 189 = 1
    16'b11000100_10111110 : OUT <= 1;  //196 / 190 = 1
    16'b11000100_10111111 : OUT <= 1;  //196 / 191 = 1
    16'b11000100_11000000 : OUT <= 1;  //196 / 192 = 1
    16'b11000100_11000001 : OUT <= 1;  //196 / 193 = 1
    16'b11000100_11000010 : OUT <= 1;  //196 / 194 = 1
    16'b11000100_11000011 : OUT <= 1;  //196 / 195 = 1
    16'b11000100_11000100 : OUT <= 1;  //196 / 196 = 1
    16'b11000100_11000101 : OUT <= 0;  //196 / 197 = 0
    16'b11000100_11000110 : OUT <= 0;  //196 / 198 = 0
    16'b11000100_11000111 : OUT <= 0;  //196 / 199 = 0
    16'b11000100_11001000 : OUT <= 0;  //196 / 200 = 0
    16'b11000100_11001001 : OUT <= 0;  //196 / 201 = 0
    16'b11000100_11001010 : OUT <= 0;  //196 / 202 = 0
    16'b11000100_11001011 : OUT <= 0;  //196 / 203 = 0
    16'b11000100_11001100 : OUT <= 0;  //196 / 204 = 0
    16'b11000100_11001101 : OUT <= 0;  //196 / 205 = 0
    16'b11000100_11001110 : OUT <= 0;  //196 / 206 = 0
    16'b11000100_11001111 : OUT <= 0;  //196 / 207 = 0
    16'b11000100_11010000 : OUT <= 0;  //196 / 208 = 0
    16'b11000100_11010001 : OUT <= 0;  //196 / 209 = 0
    16'b11000100_11010010 : OUT <= 0;  //196 / 210 = 0
    16'b11000100_11010011 : OUT <= 0;  //196 / 211 = 0
    16'b11000100_11010100 : OUT <= 0;  //196 / 212 = 0
    16'b11000100_11010101 : OUT <= 0;  //196 / 213 = 0
    16'b11000100_11010110 : OUT <= 0;  //196 / 214 = 0
    16'b11000100_11010111 : OUT <= 0;  //196 / 215 = 0
    16'b11000100_11011000 : OUT <= 0;  //196 / 216 = 0
    16'b11000100_11011001 : OUT <= 0;  //196 / 217 = 0
    16'b11000100_11011010 : OUT <= 0;  //196 / 218 = 0
    16'b11000100_11011011 : OUT <= 0;  //196 / 219 = 0
    16'b11000100_11011100 : OUT <= 0;  //196 / 220 = 0
    16'b11000100_11011101 : OUT <= 0;  //196 / 221 = 0
    16'b11000100_11011110 : OUT <= 0;  //196 / 222 = 0
    16'b11000100_11011111 : OUT <= 0;  //196 / 223 = 0
    16'b11000100_11100000 : OUT <= 0;  //196 / 224 = 0
    16'b11000100_11100001 : OUT <= 0;  //196 / 225 = 0
    16'b11000100_11100010 : OUT <= 0;  //196 / 226 = 0
    16'b11000100_11100011 : OUT <= 0;  //196 / 227 = 0
    16'b11000100_11100100 : OUT <= 0;  //196 / 228 = 0
    16'b11000100_11100101 : OUT <= 0;  //196 / 229 = 0
    16'b11000100_11100110 : OUT <= 0;  //196 / 230 = 0
    16'b11000100_11100111 : OUT <= 0;  //196 / 231 = 0
    16'b11000100_11101000 : OUT <= 0;  //196 / 232 = 0
    16'b11000100_11101001 : OUT <= 0;  //196 / 233 = 0
    16'b11000100_11101010 : OUT <= 0;  //196 / 234 = 0
    16'b11000100_11101011 : OUT <= 0;  //196 / 235 = 0
    16'b11000100_11101100 : OUT <= 0;  //196 / 236 = 0
    16'b11000100_11101101 : OUT <= 0;  //196 / 237 = 0
    16'b11000100_11101110 : OUT <= 0;  //196 / 238 = 0
    16'b11000100_11101111 : OUT <= 0;  //196 / 239 = 0
    16'b11000100_11110000 : OUT <= 0;  //196 / 240 = 0
    16'b11000100_11110001 : OUT <= 0;  //196 / 241 = 0
    16'b11000100_11110010 : OUT <= 0;  //196 / 242 = 0
    16'b11000100_11110011 : OUT <= 0;  //196 / 243 = 0
    16'b11000100_11110100 : OUT <= 0;  //196 / 244 = 0
    16'b11000100_11110101 : OUT <= 0;  //196 / 245 = 0
    16'b11000100_11110110 : OUT <= 0;  //196 / 246 = 0
    16'b11000100_11110111 : OUT <= 0;  //196 / 247 = 0
    16'b11000100_11111000 : OUT <= 0;  //196 / 248 = 0
    16'b11000100_11111001 : OUT <= 0;  //196 / 249 = 0
    16'b11000100_11111010 : OUT <= 0;  //196 / 250 = 0
    16'b11000100_11111011 : OUT <= 0;  //196 / 251 = 0
    16'b11000100_11111100 : OUT <= 0;  //196 / 252 = 0
    16'b11000100_11111101 : OUT <= 0;  //196 / 253 = 0
    16'b11000100_11111110 : OUT <= 0;  //196 / 254 = 0
    16'b11000100_11111111 : OUT <= 0;  //196 / 255 = 0
    16'b11000101_00000000 : OUT <= 0;  //197 / 0 = 0
    16'b11000101_00000001 : OUT <= 197;  //197 / 1 = 197
    16'b11000101_00000010 : OUT <= 98;  //197 / 2 = 98
    16'b11000101_00000011 : OUT <= 65;  //197 / 3 = 65
    16'b11000101_00000100 : OUT <= 49;  //197 / 4 = 49
    16'b11000101_00000101 : OUT <= 39;  //197 / 5 = 39
    16'b11000101_00000110 : OUT <= 32;  //197 / 6 = 32
    16'b11000101_00000111 : OUT <= 28;  //197 / 7 = 28
    16'b11000101_00001000 : OUT <= 24;  //197 / 8 = 24
    16'b11000101_00001001 : OUT <= 21;  //197 / 9 = 21
    16'b11000101_00001010 : OUT <= 19;  //197 / 10 = 19
    16'b11000101_00001011 : OUT <= 17;  //197 / 11 = 17
    16'b11000101_00001100 : OUT <= 16;  //197 / 12 = 16
    16'b11000101_00001101 : OUT <= 15;  //197 / 13 = 15
    16'b11000101_00001110 : OUT <= 14;  //197 / 14 = 14
    16'b11000101_00001111 : OUT <= 13;  //197 / 15 = 13
    16'b11000101_00010000 : OUT <= 12;  //197 / 16 = 12
    16'b11000101_00010001 : OUT <= 11;  //197 / 17 = 11
    16'b11000101_00010010 : OUT <= 10;  //197 / 18 = 10
    16'b11000101_00010011 : OUT <= 10;  //197 / 19 = 10
    16'b11000101_00010100 : OUT <= 9;  //197 / 20 = 9
    16'b11000101_00010101 : OUT <= 9;  //197 / 21 = 9
    16'b11000101_00010110 : OUT <= 8;  //197 / 22 = 8
    16'b11000101_00010111 : OUT <= 8;  //197 / 23 = 8
    16'b11000101_00011000 : OUT <= 8;  //197 / 24 = 8
    16'b11000101_00011001 : OUT <= 7;  //197 / 25 = 7
    16'b11000101_00011010 : OUT <= 7;  //197 / 26 = 7
    16'b11000101_00011011 : OUT <= 7;  //197 / 27 = 7
    16'b11000101_00011100 : OUT <= 7;  //197 / 28 = 7
    16'b11000101_00011101 : OUT <= 6;  //197 / 29 = 6
    16'b11000101_00011110 : OUT <= 6;  //197 / 30 = 6
    16'b11000101_00011111 : OUT <= 6;  //197 / 31 = 6
    16'b11000101_00100000 : OUT <= 6;  //197 / 32 = 6
    16'b11000101_00100001 : OUT <= 5;  //197 / 33 = 5
    16'b11000101_00100010 : OUT <= 5;  //197 / 34 = 5
    16'b11000101_00100011 : OUT <= 5;  //197 / 35 = 5
    16'b11000101_00100100 : OUT <= 5;  //197 / 36 = 5
    16'b11000101_00100101 : OUT <= 5;  //197 / 37 = 5
    16'b11000101_00100110 : OUT <= 5;  //197 / 38 = 5
    16'b11000101_00100111 : OUT <= 5;  //197 / 39 = 5
    16'b11000101_00101000 : OUT <= 4;  //197 / 40 = 4
    16'b11000101_00101001 : OUT <= 4;  //197 / 41 = 4
    16'b11000101_00101010 : OUT <= 4;  //197 / 42 = 4
    16'b11000101_00101011 : OUT <= 4;  //197 / 43 = 4
    16'b11000101_00101100 : OUT <= 4;  //197 / 44 = 4
    16'b11000101_00101101 : OUT <= 4;  //197 / 45 = 4
    16'b11000101_00101110 : OUT <= 4;  //197 / 46 = 4
    16'b11000101_00101111 : OUT <= 4;  //197 / 47 = 4
    16'b11000101_00110000 : OUT <= 4;  //197 / 48 = 4
    16'b11000101_00110001 : OUT <= 4;  //197 / 49 = 4
    16'b11000101_00110010 : OUT <= 3;  //197 / 50 = 3
    16'b11000101_00110011 : OUT <= 3;  //197 / 51 = 3
    16'b11000101_00110100 : OUT <= 3;  //197 / 52 = 3
    16'b11000101_00110101 : OUT <= 3;  //197 / 53 = 3
    16'b11000101_00110110 : OUT <= 3;  //197 / 54 = 3
    16'b11000101_00110111 : OUT <= 3;  //197 / 55 = 3
    16'b11000101_00111000 : OUT <= 3;  //197 / 56 = 3
    16'b11000101_00111001 : OUT <= 3;  //197 / 57 = 3
    16'b11000101_00111010 : OUT <= 3;  //197 / 58 = 3
    16'b11000101_00111011 : OUT <= 3;  //197 / 59 = 3
    16'b11000101_00111100 : OUT <= 3;  //197 / 60 = 3
    16'b11000101_00111101 : OUT <= 3;  //197 / 61 = 3
    16'b11000101_00111110 : OUT <= 3;  //197 / 62 = 3
    16'b11000101_00111111 : OUT <= 3;  //197 / 63 = 3
    16'b11000101_01000000 : OUT <= 3;  //197 / 64 = 3
    16'b11000101_01000001 : OUT <= 3;  //197 / 65 = 3
    16'b11000101_01000010 : OUT <= 2;  //197 / 66 = 2
    16'b11000101_01000011 : OUT <= 2;  //197 / 67 = 2
    16'b11000101_01000100 : OUT <= 2;  //197 / 68 = 2
    16'b11000101_01000101 : OUT <= 2;  //197 / 69 = 2
    16'b11000101_01000110 : OUT <= 2;  //197 / 70 = 2
    16'b11000101_01000111 : OUT <= 2;  //197 / 71 = 2
    16'b11000101_01001000 : OUT <= 2;  //197 / 72 = 2
    16'b11000101_01001001 : OUT <= 2;  //197 / 73 = 2
    16'b11000101_01001010 : OUT <= 2;  //197 / 74 = 2
    16'b11000101_01001011 : OUT <= 2;  //197 / 75 = 2
    16'b11000101_01001100 : OUT <= 2;  //197 / 76 = 2
    16'b11000101_01001101 : OUT <= 2;  //197 / 77 = 2
    16'b11000101_01001110 : OUT <= 2;  //197 / 78 = 2
    16'b11000101_01001111 : OUT <= 2;  //197 / 79 = 2
    16'b11000101_01010000 : OUT <= 2;  //197 / 80 = 2
    16'b11000101_01010001 : OUT <= 2;  //197 / 81 = 2
    16'b11000101_01010010 : OUT <= 2;  //197 / 82 = 2
    16'b11000101_01010011 : OUT <= 2;  //197 / 83 = 2
    16'b11000101_01010100 : OUT <= 2;  //197 / 84 = 2
    16'b11000101_01010101 : OUT <= 2;  //197 / 85 = 2
    16'b11000101_01010110 : OUT <= 2;  //197 / 86 = 2
    16'b11000101_01010111 : OUT <= 2;  //197 / 87 = 2
    16'b11000101_01011000 : OUT <= 2;  //197 / 88 = 2
    16'b11000101_01011001 : OUT <= 2;  //197 / 89 = 2
    16'b11000101_01011010 : OUT <= 2;  //197 / 90 = 2
    16'b11000101_01011011 : OUT <= 2;  //197 / 91 = 2
    16'b11000101_01011100 : OUT <= 2;  //197 / 92 = 2
    16'b11000101_01011101 : OUT <= 2;  //197 / 93 = 2
    16'b11000101_01011110 : OUT <= 2;  //197 / 94 = 2
    16'b11000101_01011111 : OUT <= 2;  //197 / 95 = 2
    16'b11000101_01100000 : OUT <= 2;  //197 / 96 = 2
    16'b11000101_01100001 : OUT <= 2;  //197 / 97 = 2
    16'b11000101_01100010 : OUT <= 2;  //197 / 98 = 2
    16'b11000101_01100011 : OUT <= 1;  //197 / 99 = 1
    16'b11000101_01100100 : OUT <= 1;  //197 / 100 = 1
    16'b11000101_01100101 : OUT <= 1;  //197 / 101 = 1
    16'b11000101_01100110 : OUT <= 1;  //197 / 102 = 1
    16'b11000101_01100111 : OUT <= 1;  //197 / 103 = 1
    16'b11000101_01101000 : OUT <= 1;  //197 / 104 = 1
    16'b11000101_01101001 : OUT <= 1;  //197 / 105 = 1
    16'b11000101_01101010 : OUT <= 1;  //197 / 106 = 1
    16'b11000101_01101011 : OUT <= 1;  //197 / 107 = 1
    16'b11000101_01101100 : OUT <= 1;  //197 / 108 = 1
    16'b11000101_01101101 : OUT <= 1;  //197 / 109 = 1
    16'b11000101_01101110 : OUT <= 1;  //197 / 110 = 1
    16'b11000101_01101111 : OUT <= 1;  //197 / 111 = 1
    16'b11000101_01110000 : OUT <= 1;  //197 / 112 = 1
    16'b11000101_01110001 : OUT <= 1;  //197 / 113 = 1
    16'b11000101_01110010 : OUT <= 1;  //197 / 114 = 1
    16'b11000101_01110011 : OUT <= 1;  //197 / 115 = 1
    16'b11000101_01110100 : OUT <= 1;  //197 / 116 = 1
    16'b11000101_01110101 : OUT <= 1;  //197 / 117 = 1
    16'b11000101_01110110 : OUT <= 1;  //197 / 118 = 1
    16'b11000101_01110111 : OUT <= 1;  //197 / 119 = 1
    16'b11000101_01111000 : OUT <= 1;  //197 / 120 = 1
    16'b11000101_01111001 : OUT <= 1;  //197 / 121 = 1
    16'b11000101_01111010 : OUT <= 1;  //197 / 122 = 1
    16'b11000101_01111011 : OUT <= 1;  //197 / 123 = 1
    16'b11000101_01111100 : OUT <= 1;  //197 / 124 = 1
    16'b11000101_01111101 : OUT <= 1;  //197 / 125 = 1
    16'b11000101_01111110 : OUT <= 1;  //197 / 126 = 1
    16'b11000101_01111111 : OUT <= 1;  //197 / 127 = 1
    16'b11000101_10000000 : OUT <= 1;  //197 / 128 = 1
    16'b11000101_10000001 : OUT <= 1;  //197 / 129 = 1
    16'b11000101_10000010 : OUT <= 1;  //197 / 130 = 1
    16'b11000101_10000011 : OUT <= 1;  //197 / 131 = 1
    16'b11000101_10000100 : OUT <= 1;  //197 / 132 = 1
    16'b11000101_10000101 : OUT <= 1;  //197 / 133 = 1
    16'b11000101_10000110 : OUT <= 1;  //197 / 134 = 1
    16'b11000101_10000111 : OUT <= 1;  //197 / 135 = 1
    16'b11000101_10001000 : OUT <= 1;  //197 / 136 = 1
    16'b11000101_10001001 : OUT <= 1;  //197 / 137 = 1
    16'b11000101_10001010 : OUT <= 1;  //197 / 138 = 1
    16'b11000101_10001011 : OUT <= 1;  //197 / 139 = 1
    16'b11000101_10001100 : OUT <= 1;  //197 / 140 = 1
    16'b11000101_10001101 : OUT <= 1;  //197 / 141 = 1
    16'b11000101_10001110 : OUT <= 1;  //197 / 142 = 1
    16'b11000101_10001111 : OUT <= 1;  //197 / 143 = 1
    16'b11000101_10010000 : OUT <= 1;  //197 / 144 = 1
    16'b11000101_10010001 : OUT <= 1;  //197 / 145 = 1
    16'b11000101_10010010 : OUT <= 1;  //197 / 146 = 1
    16'b11000101_10010011 : OUT <= 1;  //197 / 147 = 1
    16'b11000101_10010100 : OUT <= 1;  //197 / 148 = 1
    16'b11000101_10010101 : OUT <= 1;  //197 / 149 = 1
    16'b11000101_10010110 : OUT <= 1;  //197 / 150 = 1
    16'b11000101_10010111 : OUT <= 1;  //197 / 151 = 1
    16'b11000101_10011000 : OUT <= 1;  //197 / 152 = 1
    16'b11000101_10011001 : OUT <= 1;  //197 / 153 = 1
    16'b11000101_10011010 : OUT <= 1;  //197 / 154 = 1
    16'b11000101_10011011 : OUT <= 1;  //197 / 155 = 1
    16'b11000101_10011100 : OUT <= 1;  //197 / 156 = 1
    16'b11000101_10011101 : OUT <= 1;  //197 / 157 = 1
    16'b11000101_10011110 : OUT <= 1;  //197 / 158 = 1
    16'b11000101_10011111 : OUT <= 1;  //197 / 159 = 1
    16'b11000101_10100000 : OUT <= 1;  //197 / 160 = 1
    16'b11000101_10100001 : OUT <= 1;  //197 / 161 = 1
    16'b11000101_10100010 : OUT <= 1;  //197 / 162 = 1
    16'b11000101_10100011 : OUT <= 1;  //197 / 163 = 1
    16'b11000101_10100100 : OUT <= 1;  //197 / 164 = 1
    16'b11000101_10100101 : OUT <= 1;  //197 / 165 = 1
    16'b11000101_10100110 : OUT <= 1;  //197 / 166 = 1
    16'b11000101_10100111 : OUT <= 1;  //197 / 167 = 1
    16'b11000101_10101000 : OUT <= 1;  //197 / 168 = 1
    16'b11000101_10101001 : OUT <= 1;  //197 / 169 = 1
    16'b11000101_10101010 : OUT <= 1;  //197 / 170 = 1
    16'b11000101_10101011 : OUT <= 1;  //197 / 171 = 1
    16'b11000101_10101100 : OUT <= 1;  //197 / 172 = 1
    16'b11000101_10101101 : OUT <= 1;  //197 / 173 = 1
    16'b11000101_10101110 : OUT <= 1;  //197 / 174 = 1
    16'b11000101_10101111 : OUT <= 1;  //197 / 175 = 1
    16'b11000101_10110000 : OUT <= 1;  //197 / 176 = 1
    16'b11000101_10110001 : OUT <= 1;  //197 / 177 = 1
    16'b11000101_10110010 : OUT <= 1;  //197 / 178 = 1
    16'b11000101_10110011 : OUT <= 1;  //197 / 179 = 1
    16'b11000101_10110100 : OUT <= 1;  //197 / 180 = 1
    16'b11000101_10110101 : OUT <= 1;  //197 / 181 = 1
    16'b11000101_10110110 : OUT <= 1;  //197 / 182 = 1
    16'b11000101_10110111 : OUT <= 1;  //197 / 183 = 1
    16'b11000101_10111000 : OUT <= 1;  //197 / 184 = 1
    16'b11000101_10111001 : OUT <= 1;  //197 / 185 = 1
    16'b11000101_10111010 : OUT <= 1;  //197 / 186 = 1
    16'b11000101_10111011 : OUT <= 1;  //197 / 187 = 1
    16'b11000101_10111100 : OUT <= 1;  //197 / 188 = 1
    16'b11000101_10111101 : OUT <= 1;  //197 / 189 = 1
    16'b11000101_10111110 : OUT <= 1;  //197 / 190 = 1
    16'b11000101_10111111 : OUT <= 1;  //197 / 191 = 1
    16'b11000101_11000000 : OUT <= 1;  //197 / 192 = 1
    16'b11000101_11000001 : OUT <= 1;  //197 / 193 = 1
    16'b11000101_11000010 : OUT <= 1;  //197 / 194 = 1
    16'b11000101_11000011 : OUT <= 1;  //197 / 195 = 1
    16'b11000101_11000100 : OUT <= 1;  //197 / 196 = 1
    16'b11000101_11000101 : OUT <= 1;  //197 / 197 = 1
    16'b11000101_11000110 : OUT <= 0;  //197 / 198 = 0
    16'b11000101_11000111 : OUT <= 0;  //197 / 199 = 0
    16'b11000101_11001000 : OUT <= 0;  //197 / 200 = 0
    16'b11000101_11001001 : OUT <= 0;  //197 / 201 = 0
    16'b11000101_11001010 : OUT <= 0;  //197 / 202 = 0
    16'b11000101_11001011 : OUT <= 0;  //197 / 203 = 0
    16'b11000101_11001100 : OUT <= 0;  //197 / 204 = 0
    16'b11000101_11001101 : OUT <= 0;  //197 / 205 = 0
    16'b11000101_11001110 : OUT <= 0;  //197 / 206 = 0
    16'b11000101_11001111 : OUT <= 0;  //197 / 207 = 0
    16'b11000101_11010000 : OUT <= 0;  //197 / 208 = 0
    16'b11000101_11010001 : OUT <= 0;  //197 / 209 = 0
    16'b11000101_11010010 : OUT <= 0;  //197 / 210 = 0
    16'b11000101_11010011 : OUT <= 0;  //197 / 211 = 0
    16'b11000101_11010100 : OUT <= 0;  //197 / 212 = 0
    16'b11000101_11010101 : OUT <= 0;  //197 / 213 = 0
    16'b11000101_11010110 : OUT <= 0;  //197 / 214 = 0
    16'b11000101_11010111 : OUT <= 0;  //197 / 215 = 0
    16'b11000101_11011000 : OUT <= 0;  //197 / 216 = 0
    16'b11000101_11011001 : OUT <= 0;  //197 / 217 = 0
    16'b11000101_11011010 : OUT <= 0;  //197 / 218 = 0
    16'b11000101_11011011 : OUT <= 0;  //197 / 219 = 0
    16'b11000101_11011100 : OUT <= 0;  //197 / 220 = 0
    16'b11000101_11011101 : OUT <= 0;  //197 / 221 = 0
    16'b11000101_11011110 : OUT <= 0;  //197 / 222 = 0
    16'b11000101_11011111 : OUT <= 0;  //197 / 223 = 0
    16'b11000101_11100000 : OUT <= 0;  //197 / 224 = 0
    16'b11000101_11100001 : OUT <= 0;  //197 / 225 = 0
    16'b11000101_11100010 : OUT <= 0;  //197 / 226 = 0
    16'b11000101_11100011 : OUT <= 0;  //197 / 227 = 0
    16'b11000101_11100100 : OUT <= 0;  //197 / 228 = 0
    16'b11000101_11100101 : OUT <= 0;  //197 / 229 = 0
    16'b11000101_11100110 : OUT <= 0;  //197 / 230 = 0
    16'b11000101_11100111 : OUT <= 0;  //197 / 231 = 0
    16'b11000101_11101000 : OUT <= 0;  //197 / 232 = 0
    16'b11000101_11101001 : OUT <= 0;  //197 / 233 = 0
    16'b11000101_11101010 : OUT <= 0;  //197 / 234 = 0
    16'b11000101_11101011 : OUT <= 0;  //197 / 235 = 0
    16'b11000101_11101100 : OUT <= 0;  //197 / 236 = 0
    16'b11000101_11101101 : OUT <= 0;  //197 / 237 = 0
    16'b11000101_11101110 : OUT <= 0;  //197 / 238 = 0
    16'b11000101_11101111 : OUT <= 0;  //197 / 239 = 0
    16'b11000101_11110000 : OUT <= 0;  //197 / 240 = 0
    16'b11000101_11110001 : OUT <= 0;  //197 / 241 = 0
    16'b11000101_11110010 : OUT <= 0;  //197 / 242 = 0
    16'b11000101_11110011 : OUT <= 0;  //197 / 243 = 0
    16'b11000101_11110100 : OUT <= 0;  //197 / 244 = 0
    16'b11000101_11110101 : OUT <= 0;  //197 / 245 = 0
    16'b11000101_11110110 : OUT <= 0;  //197 / 246 = 0
    16'b11000101_11110111 : OUT <= 0;  //197 / 247 = 0
    16'b11000101_11111000 : OUT <= 0;  //197 / 248 = 0
    16'b11000101_11111001 : OUT <= 0;  //197 / 249 = 0
    16'b11000101_11111010 : OUT <= 0;  //197 / 250 = 0
    16'b11000101_11111011 : OUT <= 0;  //197 / 251 = 0
    16'b11000101_11111100 : OUT <= 0;  //197 / 252 = 0
    16'b11000101_11111101 : OUT <= 0;  //197 / 253 = 0
    16'b11000101_11111110 : OUT <= 0;  //197 / 254 = 0
    16'b11000101_11111111 : OUT <= 0;  //197 / 255 = 0
    16'b11000110_00000000 : OUT <= 0;  //198 / 0 = 0
    16'b11000110_00000001 : OUT <= 198;  //198 / 1 = 198
    16'b11000110_00000010 : OUT <= 99;  //198 / 2 = 99
    16'b11000110_00000011 : OUT <= 66;  //198 / 3 = 66
    16'b11000110_00000100 : OUT <= 49;  //198 / 4 = 49
    16'b11000110_00000101 : OUT <= 39;  //198 / 5 = 39
    16'b11000110_00000110 : OUT <= 33;  //198 / 6 = 33
    16'b11000110_00000111 : OUT <= 28;  //198 / 7 = 28
    16'b11000110_00001000 : OUT <= 24;  //198 / 8 = 24
    16'b11000110_00001001 : OUT <= 22;  //198 / 9 = 22
    16'b11000110_00001010 : OUT <= 19;  //198 / 10 = 19
    16'b11000110_00001011 : OUT <= 18;  //198 / 11 = 18
    16'b11000110_00001100 : OUT <= 16;  //198 / 12 = 16
    16'b11000110_00001101 : OUT <= 15;  //198 / 13 = 15
    16'b11000110_00001110 : OUT <= 14;  //198 / 14 = 14
    16'b11000110_00001111 : OUT <= 13;  //198 / 15 = 13
    16'b11000110_00010000 : OUT <= 12;  //198 / 16 = 12
    16'b11000110_00010001 : OUT <= 11;  //198 / 17 = 11
    16'b11000110_00010010 : OUT <= 11;  //198 / 18 = 11
    16'b11000110_00010011 : OUT <= 10;  //198 / 19 = 10
    16'b11000110_00010100 : OUT <= 9;  //198 / 20 = 9
    16'b11000110_00010101 : OUT <= 9;  //198 / 21 = 9
    16'b11000110_00010110 : OUT <= 9;  //198 / 22 = 9
    16'b11000110_00010111 : OUT <= 8;  //198 / 23 = 8
    16'b11000110_00011000 : OUT <= 8;  //198 / 24 = 8
    16'b11000110_00011001 : OUT <= 7;  //198 / 25 = 7
    16'b11000110_00011010 : OUT <= 7;  //198 / 26 = 7
    16'b11000110_00011011 : OUT <= 7;  //198 / 27 = 7
    16'b11000110_00011100 : OUT <= 7;  //198 / 28 = 7
    16'b11000110_00011101 : OUT <= 6;  //198 / 29 = 6
    16'b11000110_00011110 : OUT <= 6;  //198 / 30 = 6
    16'b11000110_00011111 : OUT <= 6;  //198 / 31 = 6
    16'b11000110_00100000 : OUT <= 6;  //198 / 32 = 6
    16'b11000110_00100001 : OUT <= 6;  //198 / 33 = 6
    16'b11000110_00100010 : OUT <= 5;  //198 / 34 = 5
    16'b11000110_00100011 : OUT <= 5;  //198 / 35 = 5
    16'b11000110_00100100 : OUT <= 5;  //198 / 36 = 5
    16'b11000110_00100101 : OUT <= 5;  //198 / 37 = 5
    16'b11000110_00100110 : OUT <= 5;  //198 / 38 = 5
    16'b11000110_00100111 : OUT <= 5;  //198 / 39 = 5
    16'b11000110_00101000 : OUT <= 4;  //198 / 40 = 4
    16'b11000110_00101001 : OUT <= 4;  //198 / 41 = 4
    16'b11000110_00101010 : OUT <= 4;  //198 / 42 = 4
    16'b11000110_00101011 : OUT <= 4;  //198 / 43 = 4
    16'b11000110_00101100 : OUT <= 4;  //198 / 44 = 4
    16'b11000110_00101101 : OUT <= 4;  //198 / 45 = 4
    16'b11000110_00101110 : OUT <= 4;  //198 / 46 = 4
    16'b11000110_00101111 : OUT <= 4;  //198 / 47 = 4
    16'b11000110_00110000 : OUT <= 4;  //198 / 48 = 4
    16'b11000110_00110001 : OUT <= 4;  //198 / 49 = 4
    16'b11000110_00110010 : OUT <= 3;  //198 / 50 = 3
    16'b11000110_00110011 : OUT <= 3;  //198 / 51 = 3
    16'b11000110_00110100 : OUT <= 3;  //198 / 52 = 3
    16'b11000110_00110101 : OUT <= 3;  //198 / 53 = 3
    16'b11000110_00110110 : OUT <= 3;  //198 / 54 = 3
    16'b11000110_00110111 : OUT <= 3;  //198 / 55 = 3
    16'b11000110_00111000 : OUT <= 3;  //198 / 56 = 3
    16'b11000110_00111001 : OUT <= 3;  //198 / 57 = 3
    16'b11000110_00111010 : OUT <= 3;  //198 / 58 = 3
    16'b11000110_00111011 : OUT <= 3;  //198 / 59 = 3
    16'b11000110_00111100 : OUT <= 3;  //198 / 60 = 3
    16'b11000110_00111101 : OUT <= 3;  //198 / 61 = 3
    16'b11000110_00111110 : OUT <= 3;  //198 / 62 = 3
    16'b11000110_00111111 : OUT <= 3;  //198 / 63 = 3
    16'b11000110_01000000 : OUT <= 3;  //198 / 64 = 3
    16'b11000110_01000001 : OUT <= 3;  //198 / 65 = 3
    16'b11000110_01000010 : OUT <= 3;  //198 / 66 = 3
    16'b11000110_01000011 : OUT <= 2;  //198 / 67 = 2
    16'b11000110_01000100 : OUT <= 2;  //198 / 68 = 2
    16'b11000110_01000101 : OUT <= 2;  //198 / 69 = 2
    16'b11000110_01000110 : OUT <= 2;  //198 / 70 = 2
    16'b11000110_01000111 : OUT <= 2;  //198 / 71 = 2
    16'b11000110_01001000 : OUT <= 2;  //198 / 72 = 2
    16'b11000110_01001001 : OUT <= 2;  //198 / 73 = 2
    16'b11000110_01001010 : OUT <= 2;  //198 / 74 = 2
    16'b11000110_01001011 : OUT <= 2;  //198 / 75 = 2
    16'b11000110_01001100 : OUT <= 2;  //198 / 76 = 2
    16'b11000110_01001101 : OUT <= 2;  //198 / 77 = 2
    16'b11000110_01001110 : OUT <= 2;  //198 / 78 = 2
    16'b11000110_01001111 : OUT <= 2;  //198 / 79 = 2
    16'b11000110_01010000 : OUT <= 2;  //198 / 80 = 2
    16'b11000110_01010001 : OUT <= 2;  //198 / 81 = 2
    16'b11000110_01010010 : OUT <= 2;  //198 / 82 = 2
    16'b11000110_01010011 : OUT <= 2;  //198 / 83 = 2
    16'b11000110_01010100 : OUT <= 2;  //198 / 84 = 2
    16'b11000110_01010101 : OUT <= 2;  //198 / 85 = 2
    16'b11000110_01010110 : OUT <= 2;  //198 / 86 = 2
    16'b11000110_01010111 : OUT <= 2;  //198 / 87 = 2
    16'b11000110_01011000 : OUT <= 2;  //198 / 88 = 2
    16'b11000110_01011001 : OUT <= 2;  //198 / 89 = 2
    16'b11000110_01011010 : OUT <= 2;  //198 / 90 = 2
    16'b11000110_01011011 : OUT <= 2;  //198 / 91 = 2
    16'b11000110_01011100 : OUT <= 2;  //198 / 92 = 2
    16'b11000110_01011101 : OUT <= 2;  //198 / 93 = 2
    16'b11000110_01011110 : OUT <= 2;  //198 / 94 = 2
    16'b11000110_01011111 : OUT <= 2;  //198 / 95 = 2
    16'b11000110_01100000 : OUT <= 2;  //198 / 96 = 2
    16'b11000110_01100001 : OUT <= 2;  //198 / 97 = 2
    16'b11000110_01100010 : OUT <= 2;  //198 / 98 = 2
    16'b11000110_01100011 : OUT <= 2;  //198 / 99 = 2
    16'b11000110_01100100 : OUT <= 1;  //198 / 100 = 1
    16'b11000110_01100101 : OUT <= 1;  //198 / 101 = 1
    16'b11000110_01100110 : OUT <= 1;  //198 / 102 = 1
    16'b11000110_01100111 : OUT <= 1;  //198 / 103 = 1
    16'b11000110_01101000 : OUT <= 1;  //198 / 104 = 1
    16'b11000110_01101001 : OUT <= 1;  //198 / 105 = 1
    16'b11000110_01101010 : OUT <= 1;  //198 / 106 = 1
    16'b11000110_01101011 : OUT <= 1;  //198 / 107 = 1
    16'b11000110_01101100 : OUT <= 1;  //198 / 108 = 1
    16'b11000110_01101101 : OUT <= 1;  //198 / 109 = 1
    16'b11000110_01101110 : OUT <= 1;  //198 / 110 = 1
    16'b11000110_01101111 : OUT <= 1;  //198 / 111 = 1
    16'b11000110_01110000 : OUT <= 1;  //198 / 112 = 1
    16'b11000110_01110001 : OUT <= 1;  //198 / 113 = 1
    16'b11000110_01110010 : OUT <= 1;  //198 / 114 = 1
    16'b11000110_01110011 : OUT <= 1;  //198 / 115 = 1
    16'b11000110_01110100 : OUT <= 1;  //198 / 116 = 1
    16'b11000110_01110101 : OUT <= 1;  //198 / 117 = 1
    16'b11000110_01110110 : OUT <= 1;  //198 / 118 = 1
    16'b11000110_01110111 : OUT <= 1;  //198 / 119 = 1
    16'b11000110_01111000 : OUT <= 1;  //198 / 120 = 1
    16'b11000110_01111001 : OUT <= 1;  //198 / 121 = 1
    16'b11000110_01111010 : OUT <= 1;  //198 / 122 = 1
    16'b11000110_01111011 : OUT <= 1;  //198 / 123 = 1
    16'b11000110_01111100 : OUT <= 1;  //198 / 124 = 1
    16'b11000110_01111101 : OUT <= 1;  //198 / 125 = 1
    16'b11000110_01111110 : OUT <= 1;  //198 / 126 = 1
    16'b11000110_01111111 : OUT <= 1;  //198 / 127 = 1
    16'b11000110_10000000 : OUT <= 1;  //198 / 128 = 1
    16'b11000110_10000001 : OUT <= 1;  //198 / 129 = 1
    16'b11000110_10000010 : OUT <= 1;  //198 / 130 = 1
    16'b11000110_10000011 : OUT <= 1;  //198 / 131 = 1
    16'b11000110_10000100 : OUT <= 1;  //198 / 132 = 1
    16'b11000110_10000101 : OUT <= 1;  //198 / 133 = 1
    16'b11000110_10000110 : OUT <= 1;  //198 / 134 = 1
    16'b11000110_10000111 : OUT <= 1;  //198 / 135 = 1
    16'b11000110_10001000 : OUT <= 1;  //198 / 136 = 1
    16'b11000110_10001001 : OUT <= 1;  //198 / 137 = 1
    16'b11000110_10001010 : OUT <= 1;  //198 / 138 = 1
    16'b11000110_10001011 : OUT <= 1;  //198 / 139 = 1
    16'b11000110_10001100 : OUT <= 1;  //198 / 140 = 1
    16'b11000110_10001101 : OUT <= 1;  //198 / 141 = 1
    16'b11000110_10001110 : OUT <= 1;  //198 / 142 = 1
    16'b11000110_10001111 : OUT <= 1;  //198 / 143 = 1
    16'b11000110_10010000 : OUT <= 1;  //198 / 144 = 1
    16'b11000110_10010001 : OUT <= 1;  //198 / 145 = 1
    16'b11000110_10010010 : OUT <= 1;  //198 / 146 = 1
    16'b11000110_10010011 : OUT <= 1;  //198 / 147 = 1
    16'b11000110_10010100 : OUT <= 1;  //198 / 148 = 1
    16'b11000110_10010101 : OUT <= 1;  //198 / 149 = 1
    16'b11000110_10010110 : OUT <= 1;  //198 / 150 = 1
    16'b11000110_10010111 : OUT <= 1;  //198 / 151 = 1
    16'b11000110_10011000 : OUT <= 1;  //198 / 152 = 1
    16'b11000110_10011001 : OUT <= 1;  //198 / 153 = 1
    16'b11000110_10011010 : OUT <= 1;  //198 / 154 = 1
    16'b11000110_10011011 : OUT <= 1;  //198 / 155 = 1
    16'b11000110_10011100 : OUT <= 1;  //198 / 156 = 1
    16'b11000110_10011101 : OUT <= 1;  //198 / 157 = 1
    16'b11000110_10011110 : OUT <= 1;  //198 / 158 = 1
    16'b11000110_10011111 : OUT <= 1;  //198 / 159 = 1
    16'b11000110_10100000 : OUT <= 1;  //198 / 160 = 1
    16'b11000110_10100001 : OUT <= 1;  //198 / 161 = 1
    16'b11000110_10100010 : OUT <= 1;  //198 / 162 = 1
    16'b11000110_10100011 : OUT <= 1;  //198 / 163 = 1
    16'b11000110_10100100 : OUT <= 1;  //198 / 164 = 1
    16'b11000110_10100101 : OUT <= 1;  //198 / 165 = 1
    16'b11000110_10100110 : OUT <= 1;  //198 / 166 = 1
    16'b11000110_10100111 : OUT <= 1;  //198 / 167 = 1
    16'b11000110_10101000 : OUT <= 1;  //198 / 168 = 1
    16'b11000110_10101001 : OUT <= 1;  //198 / 169 = 1
    16'b11000110_10101010 : OUT <= 1;  //198 / 170 = 1
    16'b11000110_10101011 : OUT <= 1;  //198 / 171 = 1
    16'b11000110_10101100 : OUT <= 1;  //198 / 172 = 1
    16'b11000110_10101101 : OUT <= 1;  //198 / 173 = 1
    16'b11000110_10101110 : OUT <= 1;  //198 / 174 = 1
    16'b11000110_10101111 : OUT <= 1;  //198 / 175 = 1
    16'b11000110_10110000 : OUT <= 1;  //198 / 176 = 1
    16'b11000110_10110001 : OUT <= 1;  //198 / 177 = 1
    16'b11000110_10110010 : OUT <= 1;  //198 / 178 = 1
    16'b11000110_10110011 : OUT <= 1;  //198 / 179 = 1
    16'b11000110_10110100 : OUT <= 1;  //198 / 180 = 1
    16'b11000110_10110101 : OUT <= 1;  //198 / 181 = 1
    16'b11000110_10110110 : OUT <= 1;  //198 / 182 = 1
    16'b11000110_10110111 : OUT <= 1;  //198 / 183 = 1
    16'b11000110_10111000 : OUT <= 1;  //198 / 184 = 1
    16'b11000110_10111001 : OUT <= 1;  //198 / 185 = 1
    16'b11000110_10111010 : OUT <= 1;  //198 / 186 = 1
    16'b11000110_10111011 : OUT <= 1;  //198 / 187 = 1
    16'b11000110_10111100 : OUT <= 1;  //198 / 188 = 1
    16'b11000110_10111101 : OUT <= 1;  //198 / 189 = 1
    16'b11000110_10111110 : OUT <= 1;  //198 / 190 = 1
    16'b11000110_10111111 : OUT <= 1;  //198 / 191 = 1
    16'b11000110_11000000 : OUT <= 1;  //198 / 192 = 1
    16'b11000110_11000001 : OUT <= 1;  //198 / 193 = 1
    16'b11000110_11000010 : OUT <= 1;  //198 / 194 = 1
    16'b11000110_11000011 : OUT <= 1;  //198 / 195 = 1
    16'b11000110_11000100 : OUT <= 1;  //198 / 196 = 1
    16'b11000110_11000101 : OUT <= 1;  //198 / 197 = 1
    16'b11000110_11000110 : OUT <= 1;  //198 / 198 = 1
    16'b11000110_11000111 : OUT <= 0;  //198 / 199 = 0
    16'b11000110_11001000 : OUT <= 0;  //198 / 200 = 0
    16'b11000110_11001001 : OUT <= 0;  //198 / 201 = 0
    16'b11000110_11001010 : OUT <= 0;  //198 / 202 = 0
    16'b11000110_11001011 : OUT <= 0;  //198 / 203 = 0
    16'b11000110_11001100 : OUT <= 0;  //198 / 204 = 0
    16'b11000110_11001101 : OUT <= 0;  //198 / 205 = 0
    16'b11000110_11001110 : OUT <= 0;  //198 / 206 = 0
    16'b11000110_11001111 : OUT <= 0;  //198 / 207 = 0
    16'b11000110_11010000 : OUT <= 0;  //198 / 208 = 0
    16'b11000110_11010001 : OUT <= 0;  //198 / 209 = 0
    16'b11000110_11010010 : OUT <= 0;  //198 / 210 = 0
    16'b11000110_11010011 : OUT <= 0;  //198 / 211 = 0
    16'b11000110_11010100 : OUT <= 0;  //198 / 212 = 0
    16'b11000110_11010101 : OUT <= 0;  //198 / 213 = 0
    16'b11000110_11010110 : OUT <= 0;  //198 / 214 = 0
    16'b11000110_11010111 : OUT <= 0;  //198 / 215 = 0
    16'b11000110_11011000 : OUT <= 0;  //198 / 216 = 0
    16'b11000110_11011001 : OUT <= 0;  //198 / 217 = 0
    16'b11000110_11011010 : OUT <= 0;  //198 / 218 = 0
    16'b11000110_11011011 : OUT <= 0;  //198 / 219 = 0
    16'b11000110_11011100 : OUT <= 0;  //198 / 220 = 0
    16'b11000110_11011101 : OUT <= 0;  //198 / 221 = 0
    16'b11000110_11011110 : OUT <= 0;  //198 / 222 = 0
    16'b11000110_11011111 : OUT <= 0;  //198 / 223 = 0
    16'b11000110_11100000 : OUT <= 0;  //198 / 224 = 0
    16'b11000110_11100001 : OUT <= 0;  //198 / 225 = 0
    16'b11000110_11100010 : OUT <= 0;  //198 / 226 = 0
    16'b11000110_11100011 : OUT <= 0;  //198 / 227 = 0
    16'b11000110_11100100 : OUT <= 0;  //198 / 228 = 0
    16'b11000110_11100101 : OUT <= 0;  //198 / 229 = 0
    16'b11000110_11100110 : OUT <= 0;  //198 / 230 = 0
    16'b11000110_11100111 : OUT <= 0;  //198 / 231 = 0
    16'b11000110_11101000 : OUT <= 0;  //198 / 232 = 0
    16'b11000110_11101001 : OUT <= 0;  //198 / 233 = 0
    16'b11000110_11101010 : OUT <= 0;  //198 / 234 = 0
    16'b11000110_11101011 : OUT <= 0;  //198 / 235 = 0
    16'b11000110_11101100 : OUT <= 0;  //198 / 236 = 0
    16'b11000110_11101101 : OUT <= 0;  //198 / 237 = 0
    16'b11000110_11101110 : OUT <= 0;  //198 / 238 = 0
    16'b11000110_11101111 : OUT <= 0;  //198 / 239 = 0
    16'b11000110_11110000 : OUT <= 0;  //198 / 240 = 0
    16'b11000110_11110001 : OUT <= 0;  //198 / 241 = 0
    16'b11000110_11110010 : OUT <= 0;  //198 / 242 = 0
    16'b11000110_11110011 : OUT <= 0;  //198 / 243 = 0
    16'b11000110_11110100 : OUT <= 0;  //198 / 244 = 0
    16'b11000110_11110101 : OUT <= 0;  //198 / 245 = 0
    16'b11000110_11110110 : OUT <= 0;  //198 / 246 = 0
    16'b11000110_11110111 : OUT <= 0;  //198 / 247 = 0
    16'b11000110_11111000 : OUT <= 0;  //198 / 248 = 0
    16'b11000110_11111001 : OUT <= 0;  //198 / 249 = 0
    16'b11000110_11111010 : OUT <= 0;  //198 / 250 = 0
    16'b11000110_11111011 : OUT <= 0;  //198 / 251 = 0
    16'b11000110_11111100 : OUT <= 0;  //198 / 252 = 0
    16'b11000110_11111101 : OUT <= 0;  //198 / 253 = 0
    16'b11000110_11111110 : OUT <= 0;  //198 / 254 = 0
    16'b11000110_11111111 : OUT <= 0;  //198 / 255 = 0
    16'b11000111_00000000 : OUT <= 0;  //199 / 0 = 0
    16'b11000111_00000001 : OUT <= 199;  //199 / 1 = 199
    16'b11000111_00000010 : OUT <= 99;  //199 / 2 = 99
    16'b11000111_00000011 : OUT <= 66;  //199 / 3 = 66
    16'b11000111_00000100 : OUT <= 49;  //199 / 4 = 49
    16'b11000111_00000101 : OUT <= 39;  //199 / 5 = 39
    16'b11000111_00000110 : OUT <= 33;  //199 / 6 = 33
    16'b11000111_00000111 : OUT <= 28;  //199 / 7 = 28
    16'b11000111_00001000 : OUT <= 24;  //199 / 8 = 24
    16'b11000111_00001001 : OUT <= 22;  //199 / 9 = 22
    16'b11000111_00001010 : OUT <= 19;  //199 / 10 = 19
    16'b11000111_00001011 : OUT <= 18;  //199 / 11 = 18
    16'b11000111_00001100 : OUT <= 16;  //199 / 12 = 16
    16'b11000111_00001101 : OUT <= 15;  //199 / 13 = 15
    16'b11000111_00001110 : OUT <= 14;  //199 / 14 = 14
    16'b11000111_00001111 : OUT <= 13;  //199 / 15 = 13
    16'b11000111_00010000 : OUT <= 12;  //199 / 16 = 12
    16'b11000111_00010001 : OUT <= 11;  //199 / 17 = 11
    16'b11000111_00010010 : OUT <= 11;  //199 / 18 = 11
    16'b11000111_00010011 : OUT <= 10;  //199 / 19 = 10
    16'b11000111_00010100 : OUT <= 9;  //199 / 20 = 9
    16'b11000111_00010101 : OUT <= 9;  //199 / 21 = 9
    16'b11000111_00010110 : OUT <= 9;  //199 / 22 = 9
    16'b11000111_00010111 : OUT <= 8;  //199 / 23 = 8
    16'b11000111_00011000 : OUT <= 8;  //199 / 24 = 8
    16'b11000111_00011001 : OUT <= 7;  //199 / 25 = 7
    16'b11000111_00011010 : OUT <= 7;  //199 / 26 = 7
    16'b11000111_00011011 : OUT <= 7;  //199 / 27 = 7
    16'b11000111_00011100 : OUT <= 7;  //199 / 28 = 7
    16'b11000111_00011101 : OUT <= 6;  //199 / 29 = 6
    16'b11000111_00011110 : OUT <= 6;  //199 / 30 = 6
    16'b11000111_00011111 : OUT <= 6;  //199 / 31 = 6
    16'b11000111_00100000 : OUT <= 6;  //199 / 32 = 6
    16'b11000111_00100001 : OUT <= 6;  //199 / 33 = 6
    16'b11000111_00100010 : OUT <= 5;  //199 / 34 = 5
    16'b11000111_00100011 : OUT <= 5;  //199 / 35 = 5
    16'b11000111_00100100 : OUT <= 5;  //199 / 36 = 5
    16'b11000111_00100101 : OUT <= 5;  //199 / 37 = 5
    16'b11000111_00100110 : OUT <= 5;  //199 / 38 = 5
    16'b11000111_00100111 : OUT <= 5;  //199 / 39 = 5
    16'b11000111_00101000 : OUT <= 4;  //199 / 40 = 4
    16'b11000111_00101001 : OUT <= 4;  //199 / 41 = 4
    16'b11000111_00101010 : OUT <= 4;  //199 / 42 = 4
    16'b11000111_00101011 : OUT <= 4;  //199 / 43 = 4
    16'b11000111_00101100 : OUT <= 4;  //199 / 44 = 4
    16'b11000111_00101101 : OUT <= 4;  //199 / 45 = 4
    16'b11000111_00101110 : OUT <= 4;  //199 / 46 = 4
    16'b11000111_00101111 : OUT <= 4;  //199 / 47 = 4
    16'b11000111_00110000 : OUT <= 4;  //199 / 48 = 4
    16'b11000111_00110001 : OUT <= 4;  //199 / 49 = 4
    16'b11000111_00110010 : OUT <= 3;  //199 / 50 = 3
    16'b11000111_00110011 : OUT <= 3;  //199 / 51 = 3
    16'b11000111_00110100 : OUT <= 3;  //199 / 52 = 3
    16'b11000111_00110101 : OUT <= 3;  //199 / 53 = 3
    16'b11000111_00110110 : OUT <= 3;  //199 / 54 = 3
    16'b11000111_00110111 : OUT <= 3;  //199 / 55 = 3
    16'b11000111_00111000 : OUT <= 3;  //199 / 56 = 3
    16'b11000111_00111001 : OUT <= 3;  //199 / 57 = 3
    16'b11000111_00111010 : OUT <= 3;  //199 / 58 = 3
    16'b11000111_00111011 : OUT <= 3;  //199 / 59 = 3
    16'b11000111_00111100 : OUT <= 3;  //199 / 60 = 3
    16'b11000111_00111101 : OUT <= 3;  //199 / 61 = 3
    16'b11000111_00111110 : OUT <= 3;  //199 / 62 = 3
    16'b11000111_00111111 : OUT <= 3;  //199 / 63 = 3
    16'b11000111_01000000 : OUT <= 3;  //199 / 64 = 3
    16'b11000111_01000001 : OUT <= 3;  //199 / 65 = 3
    16'b11000111_01000010 : OUT <= 3;  //199 / 66 = 3
    16'b11000111_01000011 : OUT <= 2;  //199 / 67 = 2
    16'b11000111_01000100 : OUT <= 2;  //199 / 68 = 2
    16'b11000111_01000101 : OUT <= 2;  //199 / 69 = 2
    16'b11000111_01000110 : OUT <= 2;  //199 / 70 = 2
    16'b11000111_01000111 : OUT <= 2;  //199 / 71 = 2
    16'b11000111_01001000 : OUT <= 2;  //199 / 72 = 2
    16'b11000111_01001001 : OUT <= 2;  //199 / 73 = 2
    16'b11000111_01001010 : OUT <= 2;  //199 / 74 = 2
    16'b11000111_01001011 : OUT <= 2;  //199 / 75 = 2
    16'b11000111_01001100 : OUT <= 2;  //199 / 76 = 2
    16'b11000111_01001101 : OUT <= 2;  //199 / 77 = 2
    16'b11000111_01001110 : OUT <= 2;  //199 / 78 = 2
    16'b11000111_01001111 : OUT <= 2;  //199 / 79 = 2
    16'b11000111_01010000 : OUT <= 2;  //199 / 80 = 2
    16'b11000111_01010001 : OUT <= 2;  //199 / 81 = 2
    16'b11000111_01010010 : OUT <= 2;  //199 / 82 = 2
    16'b11000111_01010011 : OUT <= 2;  //199 / 83 = 2
    16'b11000111_01010100 : OUT <= 2;  //199 / 84 = 2
    16'b11000111_01010101 : OUT <= 2;  //199 / 85 = 2
    16'b11000111_01010110 : OUT <= 2;  //199 / 86 = 2
    16'b11000111_01010111 : OUT <= 2;  //199 / 87 = 2
    16'b11000111_01011000 : OUT <= 2;  //199 / 88 = 2
    16'b11000111_01011001 : OUT <= 2;  //199 / 89 = 2
    16'b11000111_01011010 : OUT <= 2;  //199 / 90 = 2
    16'b11000111_01011011 : OUT <= 2;  //199 / 91 = 2
    16'b11000111_01011100 : OUT <= 2;  //199 / 92 = 2
    16'b11000111_01011101 : OUT <= 2;  //199 / 93 = 2
    16'b11000111_01011110 : OUT <= 2;  //199 / 94 = 2
    16'b11000111_01011111 : OUT <= 2;  //199 / 95 = 2
    16'b11000111_01100000 : OUT <= 2;  //199 / 96 = 2
    16'b11000111_01100001 : OUT <= 2;  //199 / 97 = 2
    16'b11000111_01100010 : OUT <= 2;  //199 / 98 = 2
    16'b11000111_01100011 : OUT <= 2;  //199 / 99 = 2
    16'b11000111_01100100 : OUT <= 1;  //199 / 100 = 1
    16'b11000111_01100101 : OUT <= 1;  //199 / 101 = 1
    16'b11000111_01100110 : OUT <= 1;  //199 / 102 = 1
    16'b11000111_01100111 : OUT <= 1;  //199 / 103 = 1
    16'b11000111_01101000 : OUT <= 1;  //199 / 104 = 1
    16'b11000111_01101001 : OUT <= 1;  //199 / 105 = 1
    16'b11000111_01101010 : OUT <= 1;  //199 / 106 = 1
    16'b11000111_01101011 : OUT <= 1;  //199 / 107 = 1
    16'b11000111_01101100 : OUT <= 1;  //199 / 108 = 1
    16'b11000111_01101101 : OUT <= 1;  //199 / 109 = 1
    16'b11000111_01101110 : OUT <= 1;  //199 / 110 = 1
    16'b11000111_01101111 : OUT <= 1;  //199 / 111 = 1
    16'b11000111_01110000 : OUT <= 1;  //199 / 112 = 1
    16'b11000111_01110001 : OUT <= 1;  //199 / 113 = 1
    16'b11000111_01110010 : OUT <= 1;  //199 / 114 = 1
    16'b11000111_01110011 : OUT <= 1;  //199 / 115 = 1
    16'b11000111_01110100 : OUT <= 1;  //199 / 116 = 1
    16'b11000111_01110101 : OUT <= 1;  //199 / 117 = 1
    16'b11000111_01110110 : OUT <= 1;  //199 / 118 = 1
    16'b11000111_01110111 : OUT <= 1;  //199 / 119 = 1
    16'b11000111_01111000 : OUT <= 1;  //199 / 120 = 1
    16'b11000111_01111001 : OUT <= 1;  //199 / 121 = 1
    16'b11000111_01111010 : OUT <= 1;  //199 / 122 = 1
    16'b11000111_01111011 : OUT <= 1;  //199 / 123 = 1
    16'b11000111_01111100 : OUT <= 1;  //199 / 124 = 1
    16'b11000111_01111101 : OUT <= 1;  //199 / 125 = 1
    16'b11000111_01111110 : OUT <= 1;  //199 / 126 = 1
    16'b11000111_01111111 : OUT <= 1;  //199 / 127 = 1
    16'b11000111_10000000 : OUT <= 1;  //199 / 128 = 1
    16'b11000111_10000001 : OUT <= 1;  //199 / 129 = 1
    16'b11000111_10000010 : OUT <= 1;  //199 / 130 = 1
    16'b11000111_10000011 : OUT <= 1;  //199 / 131 = 1
    16'b11000111_10000100 : OUT <= 1;  //199 / 132 = 1
    16'b11000111_10000101 : OUT <= 1;  //199 / 133 = 1
    16'b11000111_10000110 : OUT <= 1;  //199 / 134 = 1
    16'b11000111_10000111 : OUT <= 1;  //199 / 135 = 1
    16'b11000111_10001000 : OUT <= 1;  //199 / 136 = 1
    16'b11000111_10001001 : OUT <= 1;  //199 / 137 = 1
    16'b11000111_10001010 : OUT <= 1;  //199 / 138 = 1
    16'b11000111_10001011 : OUT <= 1;  //199 / 139 = 1
    16'b11000111_10001100 : OUT <= 1;  //199 / 140 = 1
    16'b11000111_10001101 : OUT <= 1;  //199 / 141 = 1
    16'b11000111_10001110 : OUT <= 1;  //199 / 142 = 1
    16'b11000111_10001111 : OUT <= 1;  //199 / 143 = 1
    16'b11000111_10010000 : OUT <= 1;  //199 / 144 = 1
    16'b11000111_10010001 : OUT <= 1;  //199 / 145 = 1
    16'b11000111_10010010 : OUT <= 1;  //199 / 146 = 1
    16'b11000111_10010011 : OUT <= 1;  //199 / 147 = 1
    16'b11000111_10010100 : OUT <= 1;  //199 / 148 = 1
    16'b11000111_10010101 : OUT <= 1;  //199 / 149 = 1
    16'b11000111_10010110 : OUT <= 1;  //199 / 150 = 1
    16'b11000111_10010111 : OUT <= 1;  //199 / 151 = 1
    16'b11000111_10011000 : OUT <= 1;  //199 / 152 = 1
    16'b11000111_10011001 : OUT <= 1;  //199 / 153 = 1
    16'b11000111_10011010 : OUT <= 1;  //199 / 154 = 1
    16'b11000111_10011011 : OUT <= 1;  //199 / 155 = 1
    16'b11000111_10011100 : OUT <= 1;  //199 / 156 = 1
    16'b11000111_10011101 : OUT <= 1;  //199 / 157 = 1
    16'b11000111_10011110 : OUT <= 1;  //199 / 158 = 1
    16'b11000111_10011111 : OUT <= 1;  //199 / 159 = 1
    16'b11000111_10100000 : OUT <= 1;  //199 / 160 = 1
    16'b11000111_10100001 : OUT <= 1;  //199 / 161 = 1
    16'b11000111_10100010 : OUT <= 1;  //199 / 162 = 1
    16'b11000111_10100011 : OUT <= 1;  //199 / 163 = 1
    16'b11000111_10100100 : OUT <= 1;  //199 / 164 = 1
    16'b11000111_10100101 : OUT <= 1;  //199 / 165 = 1
    16'b11000111_10100110 : OUT <= 1;  //199 / 166 = 1
    16'b11000111_10100111 : OUT <= 1;  //199 / 167 = 1
    16'b11000111_10101000 : OUT <= 1;  //199 / 168 = 1
    16'b11000111_10101001 : OUT <= 1;  //199 / 169 = 1
    16'b11000111_10101010 : OUT <= 1;  //199 / 170 = 1
    16'b11000111_10101011 : OUT <= 1;  //199 / 171 = 1
    16'b11000111_10101100 : OUT <= 1;  //199 / 172 = 1
    16'b11000111_10101101 : OUT <= 1;  //199 / 173 = 1
    16'b11000111_10101110 : OUT <= 1;  //199 / 174 = 1
    16'b11000111_10101111 : OUT <= 1;  //199 / 175 = 1
    16'b11000111_10110000 : OUT <= 1;  //199 / 176 = 1
    16'b11000111_10110001 : OUT <= 1;  //199 / 177 = 1
    16'b11000111_10110010 : OUT <= 1;  //199 / 178 = 1
    16'b11000111_10110011 : OUT <= 1;  //199 / 179 = 1
    16'b11000111_10110100 : OUT <= 1;  //199 / 180 = 1
    16'b11000111_10110101 : OUT <= 1;  //199 / 181 = 1
    16'b11000111_10110110 : OUT <= 1;  //199 / 182 = 1
    16'b11000111_10110111 : OUT <= 1;  //199 / 183 = 1
    16'b11000111_10111000 : OUT <= 1;  //199 / 184 = 1
    16'b11000111_10111001 : OUT <= 1;  //199 / 185 = 1
    16'b11000111_10111010 : OUT <= 1;  //199 / 186 = 1
    16'b11000111_10111011 : OUT <= 1;  //199 / 187 = 1
    16'b11000111_10111100 : OUT <= 1;  //199 / 188 = 1
    16'b11000111_10111101 : OUT <= 1;  //199 / 189 = 1
    16'b11000111_10111110 : OUT <= 1;  //199 / 190 = 1
    16'b11000111_10111111 : OUT <= 1;  //199 / 191 = 1
    16'b11000111_11000000 : OUT <= 1;  //199 / 192 = 1
    16'b11000111_11000001 : OUT <= 1;  //199 / 193 = 1
    16'b11000111_11000010 : OUT <= 1;  //199 / 194 = 1
    16'b11000111_11000011 : OUT <= 1;  //199 / 195 = 1
    16'b11000111_11000100 : OUT <= 1;  //199 / 196 = 1
    16'b11000111_11000101 : OUT <= 1;  //199 / 197 = 1
    16'b11000111_11000110 : OUT <= 1;  //199 / 198 = 1
    16'b11000111_11000111 : OUT <= 1;  //199 / 199 = 1
    16'b11000111_11001000 : OUT <= 0;  //199 / 200 = 0
    16'b11000111_11001001 : OUT <= 0;  //199 / 201 = 0
    16'b11000111_11001010 : OUT <= 0;  //199 / 202 = 0
    16'b11000111_11001011 : OUT <= 0;  //199 / 203 = 0
    16'b11000111_11001100 : OUT <= 0;  //199 / 204 = 0
    16'b11000111_11001101 : OUT <= 0;  //199 / 205 = 0
    16'b11000111_11001110 : OUT <= 0;  //199 / 206 = 0
    16'b11000111_11001111 : OUT <= 0;  //199 / 207 = 0
    16'b11000111_11010000 : OUT <= 0;  //199 / 208 = 0
    16'b11000111_11010001 : OUT <= 0;  //199 / 209 = 0
    16'b11000111_11010010 : OUT <= 0;  //199 / 210 = 0
    16'b11000111_11010011 : OUT <= 0;  //199 / 211 = 0
    16'b11000111_11010100 : OUT <= 0;  //199 / 212 = 0
    16'b11000111_11010101 : OUT <= 0;  //199 / 213 = 0
    16'b11000111_11010110 : OUT <= 0;  //199 / 214 = 0
    16'b11000111_11010111 : OUT <= 0;  //199 / 215 = 0
    16'b11000111_11011000 : OUT <= 0;  //199 / 216 = 0
    16'b11000111_11011001 : OUT <= 0;  //199 / 217 = 0
    16'b11000111_11011010 : OUT <= 0;  //199 / 218 = 0
    16'b11000111_11011011 : OUT <= 0;  //199 / 219 = 0
    16'b11000111_11011100 : OUT <= 0;  //199 / 220 = 0
    16'b11000111_11011101 : OUT <= 0;  //199 / 221 = 0
    16'b11000111_11011110 : OUT <= 0;  //199 / 222 = 0
    16'b11000111_11011111 : OUT <= 0;  //199 / 223 = 0
    16'b11000111_11100000 : OUT <= 0;  //199 / 224 = 0
    16'b11000111_11100001 : OUT <= 0;  //199 / 225 = 0
    16'b11000111_11100010 : OUT <= 0;  //199 / 226 = 0
    16'b11000111_11100011 : OUT <= 0;  //199 / 227 = 0
    16'b11000111_11100100 : OUT <= 0;  //199 / 228 = 0
    16'b11000111_11100101 : OUT <= 0;  //199 / 229 = 0
    16'b11000111_11100110 : OUT <= 0;  //199 / 230 = 0
    16'b11000111_11100111 : OUT <= 0;  //199 / 231 = 0
    16'b11000111_11101000 : OUT <= 0;  //199 / 232 = 0
    16'b11000111_11101001 : OUT <= 0;  //199 / 233 = 0
    16'b11000111_11101010 : OUT <= 0;  //199 / 234 = 0
    16'b11000111_11101011 : OUT <= 0;  //199 / 235 = 0
    16'b11000111_11101100 : OUT <= 0;  //199 / 236 = 0
    16'b11000111_11101101 : OUT <= 0;  //199 / 237 = 0
    16'b11000111_11101110 : OUT <= 0;  //199 / 238 = 0
    16'b11000111_11101111 : OUT <= 0;  //199 / 239 = 0
    16'b11000111_11110000 : OUT <= 0;  //199 / 240 = 0
    16'b11000111_11110001 : OUT <= 0;  //199 / 241 = 0
    16'b11000111_11110010 : OUT <= 0;  //199 / 242 = 0
    16'b11000111_11110011 : OUT <= 0;  //199 / 243 = 0
    16'b11000111_11110100 : OUT <= 0;  //199 / 244 = 0
    16'b11000111_11110101 : OUT <= 0;  //199 / 245 = 0
    16'b11000111_11110110 : OUT <= 0;  //199 / 246 = 0
    16'b11000111_11110111 : OUT <= 0;  //199 / 247 = 0
    16'b11000111_11111000 : OUT <= 0;  //199 / 248 = 0
    16'b11000111_11111001 : OUT <= 0;  //199 / 249 = 0
    16'b11000111_11111010 : OUT <= 0;  //199 / 250 = 0
    16'b11000111_11111011 : OUT <= 0;  //199 / 251 = 0
    16'b11000111_11111100 : OUT <= 0;  //199 / 252 = 0
    16'b11000111_11111101 : OUT <= 0;  //199 / 253 = 0
    16'b11000111_11111110 : OUT <= 0;  //199 / 254 = 0
    16'b11000111_11111111 : OUT <= 0;  //199 / 255 = 0
    16'b11001000_00000000 : OUT <= 0;  //200 / 0 = 0
    16'b11001000_00000001 : OUT <= 200;  //200 / 1 = 200
    16'b11001000_00000010 : OUT <= 100;  //200 / 2 = 100
    16'b11001000_00000011 : OUT <= 66;  //200 / 3 = 66
    16'b11001000_00000100 : OUT <= 50;  //200 / 4 = 50
    16'b11001000_00000101 : OUT <= 40;  //200 / 5 = 40
    16'b11001000_00000110 : OUT <= 33;  //200 / 6 = 33
    16'b11001000_00000111 : OUT <= 28;  //200 / 7 = 28
    16'b11001000_00001000 : OUT <= 25;  //200 / 8 = 25
    16'b11001000_00001001 : OUT <= 22;  //200 / 9 = 22
    16'b11001000_00001010 : OUT <= 20;  //200 / 10 = 20
    16'b11001000_00001011 : OUT <= 18;  //200 / 11 = 18
    16'b11001000_00001100 : OUT <= 16;  //200 / 12 = 16
    16'b11001000_00001101 : OUT <= 15;  //200 / 13 = 15
    16'b11001000_00001110 : OUT <= 14;  //200 / 14 = 14
    16'b11001000_00001111 : OUT <= 13;  //200 / 15 = 13
    16'b11001000_00010000 : OUT <= 12;  //200 / 16 = 12
    16'b11001000_00010001 : OUT <= 11;  //200 / 17 = 11
    16'b11001000_00010010 : OUT <= 11;  //200 / 18 = 11
    16'b11001000_00010011 : OUT <= 10;  //200 / 19 = 10
    16'b11001000_00010100 : OUT <= 10;  //200 / 20 = 10
    16'b11001000_00010101 : OUT <= 9;  //200 / 21 = 9
    16'b11001000_00010110 : OUT <= 9;  //200 / 22 = 9
    16'b11001000_00010111 : OUT <= 8;  //200 / 23 = 8
    16'b11001000_00011000 : OUT <= 8;  //200 / 24 = 8
    16'b11001000_00011001 : OUT <= 8;  //200 / 25 = 8
    16'b11001000_00011010 : OUT <= 7;  //200 / 26 = 7
    16'b11001000_00011011 : OUT <= 7;  //200 / 27 = 7
    16'b11001000_00011100 : OUT <= 7;  //200 / 28 = 7
    16'b11001000_00011101 : OUT <= 6;  //200 / 29 = 6
    16'b11001000_00011110 : OUT <= 6;  //200 / 30 = 6
    16'b11001000_00011111 : OUT <= 6;  //200 / 31 = 6
    16'b11001000_00100000 : OUT <= 6;  //200 / 32 = 6
    16'b11001000_00100001 : OUT <= 6;  //200 / 33 = 6
    16'b11001000_00100010 : OUT <= 5;  //200 / 34 = 5
    16'b11001000_00100011 : OUT <= 5;  //200 / 35 = 5
    16'b11001000_00100100 : OUT <= 5;  //200 / 36 = 5
    16'b11001000_00100101 : OUT <= 5;  //200 / 37 = 5
    16'b11001000_00100110 : OUT <= 5;  //200 / 38 = 5
    16'b11001000_00100111 : OUT <= 5;  //200 / 39 = 5
    16'b11001000_00101000 : OUT <= 5;  //200 / 40 = 5
    16'b11001000_00101001 : OUT <= 4;  //200 / 41 = 4
    16'b11001000_00101010 : OUT <= 4;  //200 / 42 = 4
    16'b11001000_00101011 : OUT <= 4;  //200 / 43 = 4
    16'b11001000_00101100 : OUT <= 4;  //200 / 44 = 4
    16'b11001000_00101101 : OUT <= 4;  //200 / 45 = 4
    16'b11001000_00101110 : OUT <= 4;  //200 / 46 = 4
    16'b11001000_00101111 : OUT <= 4;  //200 / 47 = 4
    16'b11001000_00110000 : OUT <= 4;  //200 / 48 = 4
    16'b11001000_00110001 : OUT <= 4;  //200 / 49 = 4
    16'b11001000_00110010 : OUT <= 4;  //200 / 50 = 4
    16'b11001000_00110011 : OUT <= 3;  //200 / 51 = 3
    16'b11001000_00110100 : OUT <= 3;  //200 / 52 = 3
    16'b11001000_00110101 : OUT <= 3;  //200 / 53 = 3
    16'b11001000_00110110 : OUT <= 3;  //200 / 54 = 3
    16'b11001000_00110111 : OUT <= 3;  //200 / 55 = 3
    16'b11001000_00111000 : OUT <= 3;  //200 / 56 = 3
    16'b11001000_00111001 : OUT <= 3;  //200 / 57 = 3
    16'b11001000_00111010 : OUT <= 3;  //200 / 58 = 3
    16'b11001000_00111011 : OUT <= 3;  //200 / 59 = 3
    16'b11001000_00111100 : OUT <= 3;  //200 / 60 = 3
    16'b11001000_00111101 : OUT <= 3;  //200 / 61 = 3
    16'b11001000_00111110 : OUT <= 3;  //200 / 62 = 3
    16'b11001000_00111111 : OUT <= 3;  //200 / 63 = 3
    16'b11001000_01000000 : OUT <= 3;  //200 / 64 = 3
    16'b11001000_01000001 : OUT <= 3;  //200 / 65 = 3
    16'b11001000_01000010 : OUT <= 3;  //200 / 66 = 3
    16'b11001000_01000011 : OUT <= 2;  //200 / 67 = 2
    16'b11001000_01000100 : OUT <= 2;  //200 / 68 = 2
    16'b11001000_01000101 : OUT <= 2;  //200 / 69 = 2
    16'b11001000_01000110 : OUT <= 2;  //200 / 70 = 2
    16'b11001000_01000111 : OUT <= 2;  //200 / 71 = 2
    16'b11001000_01001000 : OUT <= 2;  //200 / 72 = 2
    16'b11001000_01001001 : OUT <= 2;  //200 / 73 = 2
    16'b11001000_01001010 : OUT <= 2;  //200 / 74 = 2
    16'b11001000_01001011 : OUT <= 2;  //200 / 75 = 2
    16'b11001000_01001100 : OUT <= 2;  //200 / 76 = 2
    16'b11001000_01001101 : OUT <= 2;  //200 / 77 = 2
    16'b11001000_01001110 : OUT <= 2;  //200 / 78 = 2
    16'b11001000_01001111 : OUT <= 2;  //200 / 79 = 2
    16'b11001000_01010000 : OUT <= 2;  //200 / 80 = 2
    16'b11001000_01010001 : OUT <= 2;  //200 / 81 = 2
    16'b11001000_01010010 : OUT <= 2;  //200 / 82 = 2
    16'b11001000_01010011 : OUT <= 2;  //200 / 83 = 2
    16'b11001000_01010100 : OUT <= 2;  //200 / 84 = 2
    16'b11001000_01010101 : OUT <= 2;  //200 / 85 = 2
    16'b11001000_01010110 : OUT <= 2;  //200 / 86 = 2
    16'b11001000_01010111 : OUT <= 2;  //200 / 87 = 2
    16'b11001000_01011000 : OUT <= 2;  //200 / 88 = 2
    16'b11001000_01011001 : OUT <= 2;  //200 / 89 = 2
    16'b11001000_01011010 : OUT <= 2;  //200 / 90 = 2
    16'b11001000_01011011 : OUT <= 2;  //200 / 91 = 2
    16'b11001000_01011100 : OUT <= 2;  //200 / 92 = 2
    16'b11001000_01011101 : OUT <= 2;  //200 / 93 = 2
    16'b11001000_01011110 : OUT <= 2;  //200 / 94 = 2
    16'b11001000_01011111 : OUT <= 2;  //200 / 95 = 2
    16'b11001000_01100000 : OUT <= 2;  //200 / 96 = 2
    16'b11001000_01100001 : OUT <= 2;  //200 / 97 = 2
    16'b11001000_01100010 : OUT <= 2;  //200 / 98 = 2
    16'b11001000_01100011 : OUT <= 2;  //200 / 99 = 2
    16'b11001000_01100100 : OUT <= 2;  //200 / 100 = 2
    16'b11001000_01100101 : OUT <= 1;  //200 / 101 = 1
    16'b11001000_01100110 : OUT <= 1;  //200 / 102 = 1
    16'b11001000_01100111 : OUT <= 1;  //200 / 103 = 1
    16'b11001000_01101000 : OUT <= 1;  //200 / 104 = 1
    16'b11001000_01101001 : OUT <= 1;  //200 / 105 = 1
    16'b11001000_01101010 : OUT <= 1;  //200 / 106 = 1
    16'b11001000_01101011 : OUT <= 1;  //200 / 107 = 1
    16'b11001000_01101100 : OUT <= 1;  //200 / 108 = 1
    16'b11001000_01101101 : OUT <= 1;  //200 / 109 = 1
    16'b11001000_01101110 : OUT <= 1;  //200 / 110 = 1
    16'b11001000_01101111 : OUT <= 1;  //200 / 111 = 1
    16'b11001000_01110000 : OUT <= 1;  //200 / 112 = 1
    16'b11001000_01110001 : OUT <= 1;  //200 / 113 = 1
    16'b11001000_01110010 : OUT <= 1;  //200 / 114 = 1
    16'b11001000_01110011 : OUT <= 1;  //200 / 115 = 1
    16'b11001000_01110100 : OUT <= 1;  //200 / 116 = 1
    16'b11001000_01110101 : OUT <= 1;  //200 / 117 = 1
    16'b11001000_01110110 : OUT <= 1;  //200 / 118 = 1
    16'b11001000_01110111 : OUT <= 1;  //200 / 119 = 1
    16'b11001000_01111000 : OUT <= 1;  //200 / 120 = 1
    16'b11001000_01111001 : OUT <= 1;  //200 / 121 = 1
    16'b11001000_01111010 : OUT <= 1;  //200 / 122 = 1
    16'b11001000_01111011 : OUT <= 1;  //200 / 123 = 1
    16'b11001000_01111100 : OUT <= 1;  //200 / 124 = 1
    16'b11001000_01111101 : OUT <= 1;  //200 / 125 = 1
    16'b11001000_01111110 : OUT <= 1;  //200 / 126 = 1
    16'b11001000_01111111 : OUT <= 1;  //200 / 127 = 1
    16'b11001000_10000000 : OUT <= 1;  //200 / 128 = 1
    16'b11001000_10000001 : OUT <= 1;  //200 / 129 = 1
    16'b11001000_10000010 : OUT <= 1;  //200 / 130 = 1
    16'b11001000_10000011 : OUT <= 1;  //200 / 131 = 1
    16'b11001000_10000100 : OUT <= 1;  //200 / 132 = 1
    16'b11001000_10000101 : OUT <= 1;  //200 / 133 = 1
    16'b11001000_10000110 : OUT <= 1;  //200 / 134 = 1
    16'b11001000_10000111 : OUT <= 1;  //200 / 135 = 1
    16'b11001000_10001000 : OUT <= 1;  //200 / 136 = 1
    16'b11001000_10001001 : OUT <= 1;  //200 / 137 = 1
    16'b11001000_10001010 : OUT <= 1;  //200 / 138 = 1
    16'b11001000_10001011 : OUT <= 1;  //200 / 139 = 1
    16'b11001000_10001100 : OUT <= 1;  //200 / 140 = 1
    16'b11001000_10001101 : OUT <= 1;  //200 / 141 = 1
    16'b11001000_10001110 : OUT <= 1;  //200 / 142 = 1
    16'b11001000_10001111 : OUT <= 1;  //200 / 143 = 1
    16'b11001000_10010000 : OUT <= 1;  //200 / 144 = 1
    16'b11001000_10010001 : OUT <= 1;  //200 / 145 = 1
    16'b11001000_10010010 : OUT <= 1;  //200 / 146 = 1
    16'b11001000_10010011 : OUT <= 1;  //200 / 147 = 1
    16'b11001000_10010100 : OUT <= 1;  //200 / 148 = 1
    16'b11001000_10010101 : OUT <= 1;  //200 / 149 = 1
    16'b11001000_10010110 : OUT <= 1;  //200 / 150 = 1
    16'b11001000_10010111 : OUT <= 1;  //200 / 151 = 1
    16'b11001000_10011000 : OUT <= 1;  //200 / 152 = 1
    16'b11001000_10011001 : OUT <= 1;  //200 / 153 = 1
    16'b11001000_10011010 : OUT <= 1;  //200 / 154 = 1
    16'b11001000_10011011 : OUT <= 1;  //200 / 155 = 1
    16'b11001000_10011100 : OUT <= 1;  //200 / 156 = 1
    16'b11001000_10011101 : OUT <= 1;  //200 / 157 = 1
    16'b11001000_10011110 : OUT <= 1;  //200 / 158 = 1
    16'b11001000_10011111 : OUT <= 1;  //200 / 159 = 1
    16'b11001000_10100000 : OUT <= 1;  //200 / 160 = 1
    16'b11001000_10100001 : OUT <= 1;  //200 / 161 = 1
    16'b11001000_10100010 : OUT <= 1;  //200 / 162 = 1
    16'b11001000_10100011 : OUT <= 1;  //200 / 163 = 1
    16'b11001000_10100100 : OUT <= 1;  //200 / 164 = 1
    16'b11001000_10100101 : OUT <= 1;  //200 / 165 = 1
    16'b11001000_10100110 : OUT <= 1;  //200 / 166 = 1
    16'b11001000_10100111 : OUT <= 1;  //200 / 167 = 1
    16'b11001000_10101000 : OUT <= 1;  //200 / 168 = 1
    16'b11001000_10101001 : OUT <= 1;  //200 / 169 = 1
    16'b11001000_10101010 : OUT <= 1;  //200 / 170 = 1
    16'b11001000_10101011 : OUT <= 1;  //200 / 171 = 1
    16'b11001000_10101100 : OUT <= 1;  //200 / 172 = 1
    16'b11001000_10101101 : OUT <= 1;  //200 / 173 = 1
    16'b11001000_10101110 : OUT <= 1;  //200 / 174 = 1
    16'b11001000_10101111 : OUT <= 1;  //200 / 175 = 1
    16'b11001000_10110000 : OUT <= 1;  //200 / 176 = 1
    16'b11001000_10110001 : OUT <= 1;  //200 / 177 = 1
    16'b11001000_10110010 : OUT <= 1;  //200 / 178 = 1
    16'b11001000_10110011 : OUT <= 1;  //200 / 179 = 1
    16'b11001000_10110100 : OUT <= 1;  //200 / 180 = 1
    16'b11001000_10110101 : OUT <= 1;  //200 / 181 = 1
    16'b11001000_10110110 : OUT <= 1;  //200 / 182 = 1
    16'b11001000_10110111 : OUT <= 1;  //200 / 183 = 1
    16'b11001000_10111000 : OUT <= 1;  //200 / 184 = 1
    16'b11001000_10111001 : OUT <= 1;  //200 / 185 = 1
    16'b11001000_10111010 : OUT <= 1;  //200 / 186 = 1
    16'b11001000_10111011 : OUT <= 1;  //200 / 187 = 1
    16'b11001000_10111100 : OUT <= 1;  //200 / 188 = 1
    16'b11001000_10111101 : OUT <= 1;  //200 / 189 = 1
    16'b11001000_10111110 : OUT <= 1;  //200 / 190 = 1
    16'b11001000_10111111 : OUT <= 1;  //200 / 191 = 1
    16'b11001000_11000000 : OUT <= 1;  //200 / 192 = 1
    16'b11001000_11000001 : OUT <= 1;  //200 / 193 = 1
    16'b11001000_11000010 : OUT <= 1;  //200 / 194 = 1
    16'b11001000_11000011 : OUT <= 1;  //200 / 195 = 1
    16'b11001000_11000100 : OUT <= 1;  //200 / 196 = 1
    16'b11001000_11000101 : OUT <= 1;  //200 / 197 = 1
    16'b11001000_11000110 : OUT <= 1;  //200 / 198 = 1
    16'b11001000_11000111 : OUT <= 1;  //200 / 199 = 1
    16'b11001000_11001000 : OUT <= 1;  //200 / 200 = 1
    16'b11001000_11001001 : OUT <= 0;  //200 / 201 = 0
    16'b11001000_11001010 : OUT <= 0;  //200 / 202 = 0
    16'b11001000_11001011 : OUT <= 0;  //200 / 203 = 0
    16'b11001000_11001100 : OUT <= 0;  //200 / 204 = 0
    16'b11001000_11001101 : OUT <= 0;  //200 / 205 = 0
    16'b11001000_11001110 : OUT <= 0;  //200 / 206 = 0
    16'b11001000_11001111 : OUT <= 0;  //200 / 207 = 0
    16'b11001000_11010000 : OUT <= 0;  //200 / 208 = 0
    16'b11001000_11010001 : OUT <= 0;  //200 / 209 = 0
    16'b11001000_11010010 : OUT <= 0;  //200 / 210 = 0
    16'b11001000_11010011 : OUT <= 0;  //200 / 211 = 0
    16'b11001000_11010100 : OUT <= 0;  //200 / 212 = 0
    16'b11001000_11010101 : OUT <= 0;  //200 / 213 = 0
    16'b11001000_11010110 : OUT <= 0;  //200 / 214 = 0
    16'b11001000_11010111 : OUT <= 0;  //200 / 215 = 0
    16'b11001000_11011000 : OUT <= 0;  //200 / 216 = 0
    16'b11001000_11011001 : OUT <= 0;  //200 / 217 = 0
    16'b11001000_11011010 : OUT <= 0;  //200 / 218 = 0
    16'b11001000_11011011 : OUT <= 0;  //200 / 219 = 0
    16'b11001000_11011100 : OUT <= 0;  //200 / 220 = 0
    16'b11001000_11011101 : OUT <= 0;  //200 / 221 = 0
    16'b11001000_11011110 : OUT <= 0;  //200 / 222 = 0
    16'b11001000_11011111 : OUT <= 0;  //200 / 223 = 0
    16'b11001000_11100000 : OUT <= 0;  //200 / 224 = 0
    16'b11001000_11100001 : OUT <= 0;  //200 / 225 = 0
    16'b11001000_11100010 : OUT <= 0;  //200 / 226 = 0
    16'b11001000_11100011 : OUT <= 0;  //200 / 227 = 0
    16'b11001000_11100100 : OUT <= 0;  //200 / 228 = 0
    16'b11001000_11100101 : OUT <= 0;  //200 / 229 = 0
    16'b11001000_11100110 : OUT <= 0;  //200 / 230 = 0
    16'b11001000_11100111 : OUT <= 0;  //200 / 231 = 0
    16'b11001000_11101000 : OUT <= 0;  //200 / 232 = 0
    16'b11001000_11101001 : OUT <= 0;  //200 / 233 = 0
    16'b11001000_11101010 : OUT <= 0;  //200 / 234 = 0
    16'b11001000_11101011 : OUT <= 0;  //200 / 235 = 0
    16'b11001000_11101100 : OUT <= 0;  //200 / 236 = 0
    16'b11001000_11101101 : OUT <= 0;  //200 / 237 = 0
    16'b11001000_11101110 : OUT <= 0;  //200 / 238 = 0
    16'b11001000_11101111 : OUT <= 0;  //200 / 239 = 0
    16'b11001000_11110000 : OUT <= 0;  //200 / 240 = 0
    16'b11001000_11110001 : OUT <= 0;  //200 / 241 = 0
    16'b11001000_11110010 : OUT <= 0;  //200 / 242 = 0
    16'b11001000_11110011 : OUT <= 0;  //200 / 243 = 0
    16'b11001000_11110100 : OUT <= 0;  //200 / 244 = 0
    16'b11001000_11110101 : OUT <= 0;  //200 / 245 = 0
    16'b11001000_11110110 : OUT <= 0;  //200 / 246 = 0
    16'b11001000_11110111 : OUT <= 0;  //200 / 247 = 0
    16'b11001000_11111000 : OUT <= 0;  //200 / 248 = 0
    16'b11001000_11111001 : OUT <= 0;  //200 / 249 = 0
    16'b11001000_11111010 : OUT <= 0;  //200 / 250 = 0
    16'b11001000_11111011 : OUT <= 0;  //200 / 251 = 0
    16'b11001000_11111100 : OUT <= 0;  //200 / 252 = 0
    16'b11001000_11111101 : OUT <= 0;  //200 / 253 = 0
    16'b11001000_11111110 : OUT <= 0;  //200 / 254 = 0
    16'b11001000_11111111 : OUT <= 0;  //200 / 255 = 0
    16'b11001001_00000000 : OUT <= 0;  //201 / 0 = 0
    16'b11001001_00000001 : OUT <= 201;  //201 / 1 = 201
    16'b11001001_00000010 : OUT <= 100;  //201 / 2 = 100
    16'b11001001_00000011 : OUT <= 67;  //201 / 3 = 67
    16'b11001001_00000100 : OUT <= 50;  //201 / 4 = 50
    16'b11001001_00000101 : OUT <= 40;  //201 / 5 = 40
    16'b11001001_00000110 : OUT <= 33;  //201 / 6 = 33
    16'b11001001_00000111 : OUT <= 28;  //201 / 7 = 28
    16'b11001001_00001000 : OUT <= 25;  //201 / 8 = 25
    16'b11001001_00001001 : OUT <= 22;  //201 / 9 = 22
    16'b11001001_00001010 : OUT <= 20;  //201 / 10 = 20
    16'b11001001_00001011 : OUT <= 18;  //201 / 11 = 18
    16'b11001001_00001100 : OUT <= 16;  //201 / 12 = 16
    16'b11001001_00001101 : OUT <= 15;  //201 / 13 = 15
    16'b11001001_00001110 : OUT <= 14;  //201 / 14 = 14
    16'b11001001_00001111 : OUT <= 13;  //201 / 15 = 13
    16'b11001001_00010000 : OUT <= 12;  //201 / 16 = 12
    16'b11001001_00010001 : OUT <= 11;  //201 / 17 = 11
    16'b11001001_00010010 : OUT <= 11;  //201 / 18 = 11
    16'b11001001_00010011 : OUT <= 10;  //201 / 19 = 10
    16'b11001001_00010100 : OUT <= 10;  //201 / 20 = 10
    16'b11001001_00010101 : OUT <= 9;  //201 / 21 = 9
    16'b11001001_00010110 : OUT <= 9;  //201 / 22 = 9
    16'b11001001_00010111 : OUT <= 8;  //201 / 23 = 8
    16'b11001001_00011000 : OUT <= 8;  //201 / 24 = 8
    16'b11001001_00011001 : OUT <= 8;  //201 / 25 = 8
    16'b11001001_00011010 : OUT <= 7;  //201 / 26 = 7
    16'b11001001_00011011 : OUT <= 7;  //201 / 27 = 7
    16'b11001001_00011100 : OUT <= 7;  //201 / 28 = 7
    16'b11001001_00011101 : OUT <= 6;  //201 / 29 = 6
    16'b11001001_00011110 : OUT <= 6;  //201 / 30 = 6
    16'b11001001_00011111 : OUT <= 6;  //201 / 31 = 6
    16'b11001001_00100000 : OUT <= 6;  //201 / 32 = 6
    16'b11001001_00100001 : OUT <= 6;  //201 / 33 = 6
    16'b11001001_00100010 : OUT <= 5;  //201 / 34 = 5
    16'b11001001_00100011 : OUT <= 5;  //201 / 35 = 5
    16'b11001001_00100100 : OUT <= 5;  //201 / 36 = 5
    16'b11001001_00100101 : OUT <= 5;  //201 / 37 = 5
    16'b11001001_00100110 : OUT <= 5;  //201 / 38 = 5
    16'b11001001_00100111 : OUT <= 5;  //201 / 39 = 5
    16'b11001001_00101000 : OUT <= 5;  //201 / 40 = 5
    16'b11001001_00101001 : OUT <= 4;  //201 / 41 = 4
    16'b11001001_00101010 : OUT <= 4;  //201 / 42 = 4
    16'b11001001_00101011 : OUT <= 4;  //201 / 43 = 4
    16'b11001001_00101100 : OUT <= 4;  //201 / 44 = 4
    16'b11001001_00101101 : OUT <= 4;  //201 / 45 = 4
    16'b11001001_00101110 : OUT <= 4;  //201 / 46 = 4
    16'b11001001_00101111 : OUT <= 4;  //201 / 47 = 4
    16'b11001001_00110000 : OUT <= 4;  //201 / 48 = 4
    16'b11001001_00110001 : OUT <= 4;  //201 / 49 = 4
    16'b11001001_00110010 : OUT <= 4;  //201 / 50 = 4
    16'b11001001_00110011 : OUT <= 3;  //201 / 51 = 3
    16'b11001001_00110100 : OUT <= 3;  //201 / 52 = 3
    16'b11001001_00110101 : OUT <= 3;  //201 / 53 = 3
    16'b11001001_00110110 : OUT <= 3;  //201 / 54 = 3
    16'b11001001_00110111 : OUT <= 3;  //201 / 55 = 3
    16'b11001001_00111000 : OUT <= 3;  //201 / 56 = 3
    16'b11001001_00111001 : OUT <= 3;  //201 / 57 = 3
    16'b11001001_00111010 : OUT <= 3;  //201 / 58 = 3
    16'b11001001_00111011 : OUT <= 3;  //201 / 59 = 3
    16'b11001001_00111100 : OUT <= 3;  //201 / 60 = 3
    16'b11001001_00111101 : OUT <= 3;  //201 / 61 = 3
    16'b11001001_00111110 : OUT <= 3;  //201 / 62 = 3
    16'b11001001_00111111 : OUT <= 3;  //201 / 63 = 3
    16'b11001001_01000000 : OUT <= 3;  //201 / 64 = 3
    16'b11001001_01000001 : OUT <= 3;  //201 / 65 = 3
    16'b11001001_01000010 : OUT <= 3;  //201 / 66 = 3
    16'b11001001_01000011 : OUT <= 3;  //201 / 67 = 3
    16'b11001001_01000100 : OUT <= 2;  //201 / 68 = 2
    16'b11001001_01000101 : OUT <= 2;  //201 / 69 = 2
    16'b11001001_01000110 : OUT <= 2;  //201 / 70 = 2
    16'b11001001_01000111 : OUT <= 2;  //201 / 71 = 2
    16'b11001001_01001000 : OUT <= 2;  //201 / 72 = 2
    16'b11001001_01001001 : OUT <= 2;  //201 / 73 = 2
    16'b11001001_01001010 : OUT <= 2;  //201 / 74 = 2
    16'b11001001_01001011 : OUT <= 2;  //201 / 75 = 2
    16'b11001001_01001100 : OUT <= 2;  //201 / 76 = 2
    16'b11001001_01001101 : OUT <= 2;  //201 / 77 = 2
    16'b11001001_01001110 : OUT <= 2;  //201 / 78 = 2
    16'b11001001_01001111 : OUT <= 2;  //201 / 79 = 2
    16'b11001001_01010000 : OUT <= 2;  //201 / 80 = 2
    16'b11001001_01010001 : OUT <= 2;  //201 / 81 = 2
    16'b11001001_01010010 : OUT <= 2;  //201 / 82 = 2
    16'b11001001_01010011 : OUT <= 2;  //201 / 83 = 2
    16'b11001001_01010100 : OUT <= 2;  //201 / 84 = 2
    16'b11001001_01010101 : OUT <= 2;  //201 / 85 = 2
    16'b11001001_01010110 : OUT <= 2;  //201 / 86 = 2
    16'b11001001_01010111 : OUT <= 2;  //201 / 87 = 2
    16'b11001001_01011000 : OUT <= 2;  //201 / 88 = 2
    16'b11001001_01011001 : OUT <= 2;  //201 / 89 = 2
    16'b11001001_01011010 : OUT <= 2;  //201 / 90 = 2
    16'b11001001_01011011 : OUT <= 2;  //201 / 91 = 2
    16'b11001001_01011100 : OUT <= 2;  //201 / 92 = 2
    16'b11001001_01011101 : OUT <= 2;  //201 / 93 = 2
    16'b11001001_01011110 : OUT <= 2;  //201 / 94 = 2
    16'b11001001_01011111 : OUT <= 2;  //201 / 95 = 2
    16'b11001001_01100000 : OUT <= 2;  //201 / 96 = 2
    16'b11001001_01100001 : OUT <= 2;  //201 / 97 = 2
    16'b11001001_01100010 : OUT <= 2;  //201 / 98 = 2
    16'b11001001_01100011 : OUT <= 2;  //201 / 99 = 2
    16'b11001001_01100100 : OUT <= 2;  //201 / 100 = 2
    16'b11001001_01100101 : OUT <= 1;  //201 / 101 = 1
    16'b11001001_01100110 : OUT <= 1;  //201 / 102 = 1
    16'b11001001_01100111 : OUT <= 1;  //201 / 103 = 1
    16'b11001001_01101000 : OUT <= 1;  //201 / 104 = 1
    16'b11001001_01101001 : OUT <= 1;  //201 / 105 = 1
    16'b11001001_01101010 : OUT <= 1;  //201 / 106 = 1
    16'b11001001_01101011 : OUT <= 1;  //201 / 107 = 1
    16'b11001001_01101100 : OUT <= 1;  //201 / 108 = 1
    16'b11001001_01101101 : OUT <= 1;  //201 / 109 = 1
    16'b11001001_01101110 : OUT <= 1;  //201 / 110 = 1
    16'b11001001_01101111 : OUT <= 1;  //201 / 111 = 1
    16'b11001001_01110000 : OUT <= 1;  //201 / 112 = 1
    16'b11001001_01110001 : OUT <= 1;  //201 / 113 = 1
    16'b11001001_01110010 : OUT <= 1;  //201 / 114 = 1
    16'b11001001_01110011 : OUT <= 1;  //201 / 115 = 1
    16'b11001001_01110100 : OUT <= 1;  //201 / 116 = 1
    16'b11001001_01110101 : OUT <= 1;  //201 / 117 = 1
    16'b11001001_01110110 : OUT <= 1;  //201 / 118 = 1
    16'b11001001_01110111 : OUT <= 1;  //201 / 119 = 1
    16'b11001001_01111000 : OUT <= 1;  //201 / 120 = 1
    16'b11001001_01111001 : OUT <= 1;  //201 / 121 = 1
    16'b11001001_01111010 : OUT <= 1;  //201 / 122 = 1
    16'b11001001_01111011 : OUT <= 1;  //201 / 123 = 1
    16'b11001001_01111100 : OUT <= 1;  //201 / 124 = 1
    16'b11001001_01111101 : OUT <= 1;  //201 / 125 = 1
    16'b11001001_01111110 : OUT <= 1;  //201 / 126 = 1
    16'b11001001_01111111 : OUT <= 1;  //201 / 127 = 1
    16'b11001001_10000000 : OUT <= 1;  //201 / 128 = 1
    16'b11001001_10000001 : OUT <= 1;  //201 / 129 = 1
    16'b11001001_10000010 : OUT <= 1;  //201 / 130 = 1
    16'b11001001_10000011 : OUT <= 1;  //201 / 131 = 1
    16'b11001001_10000100 : OUT <= 1;  //201 / 132 = 1
    16'b11001001_10000101 : OUT <= 1;  //201 / 133 = 1
    16'b11001001_10000110 : OUT <= 1;  //201 / 134 = 1
    16'b11001001_10000111 : OUT <= 1;  //201 / 135 = 1
    16'b11001001_10001000 : OUT <= 1;  //201 / 136 = 1
    16'b11001001_10001001 : OUT <= 1;  //201 / 137 = 1
    16'b11001001_10001010 : OUT <= 1;  //201 / 138 = 1
    16'b11001001_10001011 : OUT <= 1;  //201 / 139 = 1
    16'b11001001_10001100 : OUT <= 1;  //201 / 140 = 1
    16'b11001001_10001101 : OUT <= 1;  //201 / 141 = 1
    16'b11001001_10001110 : OUT <= 1;  //201 / 142 = 1
    16'b11001001_10001111 : OUT <= 1;  //201 / 143 = 1
    16'b11001001_10010000 : OUT <= 1;  //201 / 144 = 1
    16'b11001001_10010001 : OUT <= 1;  //201 / 145 = 1
    16'b11001001_10010010 : OUT <= 1;  //201 / 146 = 1
    16'b11001001_10010011 : OUT <= 1;  //201 / 147 = 1
    16'b11001001_10010100 : OUT <= 1;  //201 / 148 = 1
    16'b11001001_10010101 : OUT <= 1;  //201 / 149 = 1
    16'b11001001_10010110 : OUT <= 1;  //201 / 150 = 1
    16'b11001001_10010111 : OUT <= 1;  //201 / 151 = 1
    16'b11001001_10011000 : OUT <= 1;  //201 / 152 = 1
    16'b11001001_10011001 : OUT <= 1;  //201 / 153 = 1
    16'b11001001_10011010 : OUT <= 1;  //201 / 154 = 1
    16'b11001001_10011011 : OUT <= 1;  //201 / 155 = 1
    16'b11001001_10011100 : OUT <= 1;  //201 / 156 = 1
    16'b11001001_10011101 : OUT <= 1;  //201 / 157 = 1
    16'b11001001_10011110 : OUT <= 1;  //201 / 158 = 1
    16'b11001001_10011111 : OUT <= 1;  //201 / 159 = 1
    16'b11001001_10100000 : OUT <= 1;  //201 / 160 = 1
    16'b11001001_10100001 : OUT <= 1;  //201 / 161 = 1
    16'b11001001_10100010 : OUT <= 1;  //201 / 162 = 1
    16'b11001001_10100011 : OUT <= 1;  //201 / 163 = 1
    16'b11001001_10100100 : OUT <= 1;  //201 / 164 = 1
    16'b11001001_10100101 : OUT <= 1;  //201 / 165 = 1
    16'b11001001_10100110 : OUT <= 1;  //201 / 166 = 1
    16'b11001001_10100111 : OUT <= 1;  //201 / 167 = 1
    16'b11001001_10101000 : OUT <= 1;  //201 / 168 = 1
    16'b11001001_10101001 : OUT <= 1;  //201 / 169 = 1
    16'b11001001_10101010 : OUT <= 1;  //201 / 170 = 1
    16'b11001001_10101011 : OUT <= 1;  //201 / 171 = 1
    16'b11001001_10101100 : OUT <= 1;  //201 / 172 = 1
    16'b11001001_10101101 : OUT <= 1;  //201 / 173 = 1
    16'b11001001_10101110 : OUT <= 1;  //201 / 174 = 1
    16'b11001001_10101111 : OUT <= 1;  //201 / 175 = 1
    16'b11001001_10110000 : OUT <= 1;  //201 / 176 = 1
    16'b11001001_10110001 : OUT <= 1;  //201 / 177 = 1
    16'b11001001_10110010 : OUT <= 1;  //201 / 178 = 1
    16'b11001001_10110011 : OUT <= 1;  //201 / 179 = 1
    16'b11001001_10110100 : OUT <= 1;  //201 / 180 = 1
    16'b11001001_10110101 : OUT <= 1;  //201 / 181 = 1
    16'b11001001_10110110 : OUT <= 1;  //201 / 182 = 1
    16'b11001001_10110111 : OUT <= 1;  //201 / 183 = 1
    16'b11001001_10111000 : OUT <= 1;  //201 / 184 = 1
    16'b11001001_10111001 : OUT <= 1;  //201 / 185 = 1
    16'b11001001_10111010 : OUT <= 1;  //201 / 186 = 1
    16'b11001001_10111011 : OUT <= 1;  //201 / 187 = 1
    16'b11001001_10111100 : OUT <= 1;  //201 / 188 = 1
    16'b11001001_10111101 : OUT <= 1;  //201 / 189 = 1
    16'b11001001_10111110 : OUT <= 1;  //201 / 190 = 1
    16'b11001001_10111111 : OUT <= 1;  //201 / 191 = 1
    16'b11001001_11000000 : OUT <= 1;  //201 / 192 = 1
    16'b11001001_11000001 : OUT <= 1;  //201 / 193 = 1
    16'b11001001_11000010 : OUT <= 1;  //201 / 194 = 1
    16'b11001001_11000011 : OUT <= 1;  //201 / 195 = 1
    16'b11001001_11000100 : OUT <= 1;  //201 / 196 = 1
    16'b11001001_11000101 : OUT <= 1;  //201 / 197 = 1
    16'b11001001_11000110 : OUT <= 1;  //201 / 198 = 1
    16'b11001001_11000111 : OUT <= 1;  //201 / 199 = 1
    16'b11001001_11001000 : OUT <= 1;  //201 / 200 = 1
    16'b11001001_11001001 : OUT <= 1;  //201 / 201 = 1
    16'b11001001_11001010 : OUT <= 0;  //201 / 202 = 0
    16'b11001001_11001011 : OUT <= 0;  //201 / 203 = 0
    16'b11001001_11001100 : OUT <= 0;  //201 / 204 = 0
    16'b11001001_11001101 : OUT <= 0;  //201 / 205 = 0
    16'b11001001_11001110 : OUT <= 0;  //201 / 206 = 0
    16'b11001001_11001111 : OUT <= 0;  //201 / 207 = 0
    16'b11001001_11010000 : OUT <= 0;  //201 / 208 = 0
    16'b11001001_11010001 : OUT <= 0;  //201 / 209 = 0
    16'b11001001_11010010 : OUT <= 0;  //201 / 210 = 0
    16'b11001001_11010011 : OUT <= 0;  //201 / 211 = 0
    16'b11001001_11010100 : OUT <= 0;  //201 / 212 = 0
    16'b11001001_11010101 : OUT <= 0;  //201 / 213 = 0
    16'b11001001_11010110 : OUT <= 0;  //201 / 214 = 0
    16'b11001001_11010111 : OUT <= 0;  //201 / 215 = 0
    16'b11001001_11011000 : OUT <= 0;  //201 / 216 = 0
    16'b11001001_11011001 : OUT <= 0;  //201 / 217 = 0
    16'b11001001_11011010 : OUT <= 0;  //201 / 218 = 0
    16'b11001001_11011011 : OUT <= 0;  //201 / 219 = 0
    16'b11001001_11011100 : OUT <= 0;  //201 / 220 = 0
    16'b11001001_11011101 : OUT <= 0;  //201 / 221 = 0
    16'b11001001_11011110 : OUT <= 0;  //201 / 222 = 0
    16'b11001001_11011111 : OUT <= 0;  //201 / 223 = 0
    16'b11001001_11100000 : OUT <= 0;  //201 / 224 = 0
    16'b11001001_11100001 : OUT <= 0;  //201 / 225 = 0
    16'b11001001_11100010 : OUT <= 0;  //201 / 226 = 0
    16'b11001001_11100011 : OUT <= 0;  //201 / 227 = 0
    16'b11001001_11100100 : OUT <= 0;  //201 / 228 = 0
    16'b11001001_11100101 : OUT <= 0;  //201 / 229 = 0
    16'b11001001_11100110 : OUT <= 0;  //201 / 230 = 0
    16'b11001001_11100111 : OUT <= 0;  //201 / 231 = 0
    16'b11001001_11101000 : OUT <= 0;  //201 / 232 = 0
    16'b11001001_11101001 : OUT <= 0;  //201 / 233 = 0
    16'b11001001_11101010 : OUT <= 0;  //201 / 234 = 0
    16'b11001001_11101011 : OUT <= 0;  //201 / 235 = 0
    16'b11001001_11101100 : OUT <= 0;  //201 / 236 = 0
    16'b11001001_11101101 : OUT <= 0;  //201 / 237 = 0
    16'b11001001_11101110 : OUT <= 0;  //201 / 238 = 0
    16'b11001001_11101111 : OUT <= 0;  //201 / 239 = 0
    16'b11001001_11110000 : OUT <= 0;  //201 / 240 = 0
    16'b11001001_11110001 : OUT <= 0;  //201 / 241 = 0
    16'b11001001_11110010 : OUT <= 0;  //201 / 242 = 0
    16'b11001001_11110011 : OUT <= 0;  //201 / 243 = 0
    16'b11001001_11110100 : OUT <= 0;  //201 / 244 = 0
    16'b11001001_11110101 : OUT <= 0;  //201 / 245 = 0
    16'b11001001_11110110 : OUT <= 0;  //201 / 246 = 0
    16'b11001001_11110111 : OUT <= 0;  //201 / 247 = 0
    16'b11001001_11111000 : OUT <= 0;  //201 / 248 = 0
    16'b11001001_11111001 : OUT <= 0;  //201 / 249 = 0
    16'b11001001_11111010 : OUT <= 0;  //201 / 250 = 0
    16'b11001001_11111011 : OUT <= 0;  //201 / 251 = 0
    16'b11001001_11111100 : OUT <= 0;  //201 / 252 = 0
    16'b11001001_11111101 : OUT <= 0;  //201 / 253 = 0
    16'b11001001_11111110 : OUT <= 0;  //201 / 254 = 0
    16'b11001001_11111111 : OUT <= 0;  //201 / 255 = 0
    16'b11001010_00000000 : OUT <= 0;  //202 / 0 = 0
    16'b11001010_00000001 : OUT <= 202;  //202 / 1 = 202
    16'b11001010_00000010 : OUT <= 101;  //202 / 2 = 101
    16'b11001010_00000011 : OUT <= 67;  //202 / 3 = 67
    16'b11001010_00000100 : OUT <= 50;  //202 / 4 = 50
    16'b11001010_00000101 : OUT <= 40;  //202 / 5 = 40
    16'b11001010_00000110 : OUT <= 33;  //202 / 6 = 33
    16'b11001010_00000111 : OUT <= 28;  //202 / 7 = 28
    16'b11001010_00001000 : OUT <= 25;  //202 / 8 = 25
    16'b11001010_00001001 : OUT <= 22;  //202 / 9 = 22
    16'b11001010_00001010 : OUT <= 20;  //202 / 10 = 20
    16'b11001010_00001011 : OUT <= 18;  //202 / 11 = 18
    16'b11001010_00001100 : OUT <= 16;  //202 / 12 = 16
    16'b11001010_00001101 : OUT <= 15;  //202 / 13 = 15
    16'b11001010_00001110 : OUT <= 14;  //202 / 14 = 14
    16'b11001010_00001111 : OUT <= 13;  //202 / 15 = 13
    16'b11001010_00010000 : OUT <= 12;  //202 / 16 = 12
    16'b11001010_00010001 : OUT <= 11;  //202 / 17 = 11
    16'b11001010_00010010 : OUT <= 11;  //202 / 18 = 11
    16'b11001010_00010011 : OUT <= 10;  //202 / 19 = 10
    16'b11001010_00010100 : OUT <= 10;  //202 / 20 = 10
    16'b11001010_00010101 : OUT <= 9;  //202 / 21 = 9
    16'b11001010_00010110 : OUT <= 9;  //202 / 22 = 9
    16'b11001010_00010111 : OUT <= 8;  //202 / 23 = 8
    16'b11001010_00011000 : OUT <= 8;  //202 / 24 = 8
    16'b11001010_00011001 : OUT <= 8;  //202 / 25 = 8
    16'b11001010_00011010 : OUT <= 7;  //202 / 26 = 7
    16'b11001010_00011011 : OUT <= 7;  //202 / 27 = 7
    16'b11001010_00011100 : OUT <= 7;  //202 / 28 = 7
    16'b11001010_00011101 : OUT <= 6;  //202 / 29 = 6
    16'b11001010_00011110 : OUT <= 6;  //202 / 30 = 6
    16'b11001010_00011111 : OUT <= 6;  //202 / 31 = 6
    16'b11001010_00100000 : OUT <= 6;  //202 / 32 = 6
    16'b11001010_00100001 : OUT <= 6;  //202 / 33 = 6
    16'b11001010_00100010 : OUT <= 5;  //202 / 34 = 5
    16'b11001010_00100011 : OUT <= 5;  //202 / 35 = 5
    16'b11001010_00100100 : OUT <= 5;  //202 / 36 = 5
    16'b11001010_00100101 : OUT <= 5;  //202 / 37 = 5
    16'b11001010_00100110 : OUT <= 5;  //202 / 38 = 5
    16'b11001010_00100111 : OUT <= 5;  //202 / 39 = 5
    16'b11001010_00101000 : OUT <= 5;  //202 / 40 = 5
    16'b11001010_00101001 : OUT <= 4;  //202 / 41 = 4
    16'b11001010_00101010 : OUT <= 4;  //202 / 42 = 4
    16'b11001010_00101011 : OUT <= 4;  //202 / 43 = 4
    16'b11001010_00101100 : OUT <= 4;  //202 / 44 = 4
    16'b11001010_00101101 : OUT <= 4;  //202 / 45 = 4
    16'b11001010_00101110 : OUT <= 4;  //202 / 46 = 4
    16'b11001010_00101111 : OUT <= 4;  //202 / 47 = 4
    16'b11001010_00110000 : OUT <= 4;  //202 / 48 = 4
    16'b11001010_00110001 : OUT <= 4;  //202 / 49 = 4
    16'b11001010_00110010 : OUT <= 4;  //202 / 50 = 4
    16'b11001010_00110011 : OUT <= 3;  //202 / 51 = 3
    16'b11001010_00110100 : OUT <= 3;  //202 / 52 = 3
    16'b11001010_00110101 : OUT <= 3;  //202 / 53 = 3
    16'b11001010_00110110 : OUT <= 3;  //202 / 54 = 3
    16'b11001010_00110111 : OUT <= 3;  //202 / 55 = 3
    16'b11001010_00111000 : OUT <= 3;  //202 / 56 = 3
    16'b11001010_00111001 : OUT <= 3;  //202 / 57 = 3
    16'b11001010_00111010 : OUT <= 3;  //202 / 58 = 3
    16'b11001010_00111011 : OUT <= 3;  //202 / 59 = 3
    16'b11001010_00111100 : OUT <= 3;  //202 / 60 = 3
    16'b11001010_00111101 : OUT <= 3;  //202 / 61 = 3
    16'b11001010_00111110 : OUT <= 3;  //202 / 62 = 3
    16'b11001010_00111111 : OUT <= 3;  //202 / 63 = 3
    16'b11001010_01000000 : OUT <= 3;  //202 / 64 = 3
    16'b11001010_01000001 : OUT <= 3;  //202 / 65 = 3
    16'b11001010_01000010 : OUT <= 3;  //202 / 66 = 3
    16'b11001010_01000011 : OUT <= 3;  //202 / 67 = 3
    16'b11001010_01000100 : OUT <= 2;  //202 / 68 = 2
    16'b11001010_01000101 : OUT <= 2;  //202 / 69 = 2
    16'b11001010_01000110 : OUT <= 2;  //202 / 70 = 2
    16'b11001010_01000111 : OUT <= 2;  //202 / 71 = 2
    16'b11001010_01001000 : OUT <= 2;  //202 / 72 = 2
    16'b11001010_01001001 : OUT <= 2;  //202 / 73 = 2
    16'b11001010_01001010 : OUT <= 2;  //202 / 74 = 2
    16'b11001010_01001011 : OUT <= 2;  //202 / 75 = 2
    16'b11001010_01001100 : OUT <= 2;  //202 / 76 = 2
    16'b11001010_01001101 : OUT <= 2;  //202 / 77 = 2
    16'b11001010_01001110 : OUT <= 2;  //202 / 78 = 2
    16'b11001010_01001111 : OUT <= 2;  //202 / 79 = 2
    16'b11001010_01010000 : OUT <= 2;  //202 / 80 = 2
    16'b11001010_01010001 : OUT <= 2;  //202 / 81 = 2
    16'b11001010_01010010 : OUT <= 2;  //202 / 82 = 2
    16'b11001010_01010011 : OUT <= 2;  //202 / 83 = 2
    16'b11001010_01010100 : OUT <= 2;  //202 / 84 = 2
    16'b11001010_01010101 : OUT <= 2;  //202 / 85 = 2
    16'b11001010_01010110 : OUT <= 2;  //202 / 86 = 2
    16'b11001010_01010111 : OUT <= 2;  //202 / 87 = 2
    16'b11001010_01011000 : OUT <= 2;  //202 / 88 = 2
    16'b11001010_01011001 : OUT <= 2;  //202 / 89 = 2
    16'b11001010_01011010 : OUT <= 2;  //202 / 90 = 2
    16'b11001010_01011011 : OUT <= 2;  //202 / 91 = 2
    16'b11001010_01011100 : OUT <= 2;  //202 / 92 = 2
    16'b11001010_01011101 : OUT <= 2;  //202 / 93 = 2
    16'b11001010_01011110 : OUT <= 2;  //202 / 94 = 2
    16'b11001010_01011111 : OUT <= 2;  //202 / 95 = 2
    16'b11001010_01100000 : OUT <= 2;  //202 / 96 = 2
    16'b11001010_01100001 : OUT <= 2;  //202 / 97 = 2
    16'b11001010_01100010 : OUT <= 2;  //202 / 98 = 2
    16'b11001010_01100011 : OUT <= 2;  //202 / 99 = 2
    16'b11001010_01100100 : OUT <= 2;  //202 / 100 = 2
    16'b11001010_01100101 : OUT <= 2;  //202 / 101 = 2
    16'b11001010_01100110 : OUT <= 1;  //202 / 102 = 1
    16'b11001010_01100111 : OUT <= 1;  //202 / 103 = 1
    16'b11001010_01101000 : OUT <= 1;  //202 / 104 = 1
    16'b11001010_01101001 : OUT <= 1;  //202 / 105 = 1
    16'b11001010_01101010 : OUT <= 1;  //202 / 106 = 1
    16'b11001010_01101011 : OUT <= 1;  //202 / 107 = 1
    16'b11001010_01101100 : OUT <= 1;  //202 / 108 = 1
    16'b11001010_01101101 : OUT <= 1;  //202 / 109 = 1
    16'b11001010_01101110 : OUT <= 1;  //202 / 110 = 1
    16'b11001010_01101111 : OUT <= 1;  //202 / 111 = 1
    16'b11001010_01110000 : OUT <= 1;  //202 / 112 = 1
    16'b11001010_01110001 : OUT <= 1;  //202 / 113 = 1
    16'b11001010_01110010 : OUT <= 1;  //202 / 114 = 1
    16'b11001010_01110011 : OUT <= 1;  //202 / 115 = 1
    16'b11001010_01110100 : OUT <= 1;  //202 / 116 = 1
    16'b11001010_01110101 : OUT <= 1;  //202 / 117 = 1
    16'b11001010_01110110 : OUT <= 1;  //202 / 118 = 1
    16'b11001010_01110111 : OUT <= 1;  //202 / 119 = 1
    16'b11001010_01111000 : OUT <= 1;  //202 / 120 = 1
    16'b11001010_01111001 : OUT <= 1;  //202 / 121 = 1
    16'b11001010_01111010 : OUT <= 1;  //202 / 122 = 1
    16'b11001010_01111011 : OUT <= 1;  //202 / 123 = 1
    16'b11001010_01111100 : OUT <= 1;  //202 / 124 = 1
    16'b11001010_01111101 : OUT <= 1;  //202 / 125 = 1
    16'b11001010_01111110 : OUT <= 1;  //202 / 126 = 1
    16'b11001010_01111111 : OUT <= 1;  //202 / 127 = 1
    16'b11001010_10000000 : OUT <= 1;  //202 / 128 = 1
    16'b11001010_10000001 : OUT <= 1;  //202 / 129 = 1
    16'b11001010_10000010 : OUT <= 1;  //202 / 130 = 1
    16'b11001010_10000011 : OUT <= 1;  //202 / 131 = 1
    16'b11001010_10000100 : OUT <= 1;  //202 / 132 = 1
    16'b11001010_10000101 : OUT <= 1;  //202 / 133 = 1
    16'b11001010_10000110 : OUT <= 1;  //202 / 134 = 1
    16'b11001010_10000111 : OUT <= 1;  //202 / 135 = 1
    16'b11001010_10001000 : OUT <= 1;  //202 / 136 = 1
    16'b11001010_10001001 : OUT <= 1;  //202 / 137 = 1
    16'b11001010_10001010 : OUT <= 1;  //202 / 138 = 1
    16'b11001010_10001011 : OUT <= 1;  //202 / 139 = 1
    16'b11001010_10001100 : OUT <= 1;  //202 / 140 = 1
    16'b11001010_10001101 : OUT <= 1;  //202 / 141 = 1
    16'b11001010_10001110 : OUT <= 1;  //202 / 142 = 1
    16'b11001010_10001111 : OUT <= 1;  //202 / 143 = 1
    16'b11001010_10010000 : OUT <= 1;  //202 / 144 = 1
    16'b11001010_10010001 : OUT <= 1;  //202 / 145 = 1
    16'b11001010_10010010 : OUT <= 1;  //202 / 146 = 1
    16'b11001010_10010011 : OUT <= 1;  //202 / 147 = 1
    16'b11001010_10010100 : OUT <= 1;  //202 / 148 = 1
    16'b11001010_10010101 : OUT <= 1;  //202 / 149 = 1
    16'b11001010_10010110 : OUT <= 1;  //202 / 150 = 1
    16'b11001010_10010111 : OUT <= 1;  //202 / 151 = 1
    16'b11001010_10011000 : OUT <= 1;  //202 / 152 = 1
    16'b11001010_10011001 : OUT <= 1;  //202 / 153 = 1
    16'b11001010_10011010 : OUT <= 1;  //202 / 154 = 1
    16'b11001010_10011011 : OUT <= 1;  //202 / 155 = 1
    16'b11001010_10011100 : OUT <= 1;  //202 / 156 = 1
    16'b11001010_10011101 : OUT <= 1;  //202 / 157 = 1
    16'b11001010_10011110 : OUT <= 1;  //202 / 158 = 1
    16'b11001010_10011111 : OUT <= 1;  //202 / 159 = 1
    16'b11001010_10100000 : OUT <= 1;  //202 / 160 = 1
    16'b11001010_10100001 : OUT <= 1;  //202 / 161 = 1
    16'b11001010_10100010 : OUT <= 1;  //202 / 162 = 1
    16'b11001010_10100011 : OUT <= 1;  //202 / 163 = 1
    16'b11001010_10100100 : OUT <= 1;  //202 / 164 = 1
    16'b11001010_10100101 : OUT <= 1;  //202 / 165 = 1
    16'b11001010_10100110 : OUT <= 1;  //202 / 166 = 1
    16'b11001010_10100111 : OUT <= 1;  //202 / 167 = 1
    16'b11001010_10101000 : OUT <= 1;  //202 / 168 = 1
    16'b11001010_10101001 : OUT <= 1;  //202 / 169 = 1
    16'b11001010_10101010 : OUT <= 1;  //202 / 170 = 1
    16'b11001010_10101011 : OUT <= 1;  //202 / 171 = 1
    16'b11001010_10101100 : OUT <= 1;  //202 / 172 = 1
    16'b11001010_10101101 : OUT <= 1;  //202 / 173 = 1
    16'b11001010_10101110 : OUT <= 1;  //202 / 174 = 1
    16'b11001010_10101111 : OUT <= 1;  //202 / 175 = 1
    16'b11001010_10110000 : OUT <= 1;  //202 / 176 = 1
    16'b11001010_10110001 : OUT <= 1;  //202 / 177 = 1
    16'b11001010_10110010 : OUT <= 1;  //202 / 178 = 1
    16'b11001010_10110011 : OUT <= 1;  //202 / 179 = 1
    16'b11001010_10110100 : OUT <= 1;  //202 / 180 = 1
    16'b11001010_10110101 : OUT <= 1;  //202 / 181 = 1
    16'b11001010_10110110 : OUT <= 1;  //202 / 182 = 1
    16'b11001010_10110111 : OUT <= 1;  //202 / 183 = 1
    16'b11001010_10111000 : OUT <= 1;  //202 / 184 = 1
    16'b11001010_10111001 : OUT <= 1;  //202 / 185 = 1
    16'b11001010_10111010 : OUT <= 1;  //202 / 186 = 1
    16'b11001010_10111011 : OUT <= 1;  //202 / 187 = 1
    16'b11001010_10111100 : OUT <= 1;  //202 / 188 = 1
    16'b11001010_10111101 : OUT <= 1;  //202 / 189 = 1
    16'b11001010_10111110 : OUT <= 1;  //202 / 190 = 1
    16'b11001010_10111111 : OUT <= 1;  //202 / 191 = 1
    16'b11001010_11000000 : OUT <= 1;  //202 / 192 = 1
    16'b11001010_11000001 : OUT <= 1;  //202 / 193 = 1
    16'b11001010_11000010 : OUT <= 1;  //202 / 194 = 1
    16'b11001010_11000011 : OUT <= 1;  //202 / 195 = 1
    16'b11001010_11000100 : OUT <= 1;  //202 / 196 = 1
    16'b11001010_11000101 : OUT <= 1;  //202 / 197 = 1
    16'b11001010_11000110 : OUT <= 1;  //202 / 198 = 1
    16'b11001010_11000111 : OUT <= 1;  //202 / 199 = 1
    16'b11001010_11001000 : OUT <= 1;  //202 / 200 = 1
    16'b11001010_11001001 : OUT <= 1;  //202 / 201 = 1
    16'b11001010_11001010 : OUT <= 1;  //202 / 202 = 1
    16'b11001010_11001011 : OUT <= 0;  //202 / 203 = 0
    16'b11001010_11001100 : OUT <= 0;  //202 / 204 = 0
    16'b11001010_11001101 : OUT <= 0;  //202 / 205 = 0
    16'b11001010_11001110 : OUT <= 0;  //202 / 206 = 0
    16'b11001010_11001111 : OUT <= 0;  //202 / 207 = 0
    16'b11001010_11010000 : OUT <= 0;  //202 / 208 = 0
    16'b11001010_11010001 : OUT <= 0;  //202 / 209 = 0
    16'b11001010_11010010 : OUT <= 0;  //202 / 210 = 0
    16'b11001010_11010011 : OUT <= 0;  //202 / 211 = 0
    16'b11001010_11010100 : OUT <= 0;  //202 / 212 = 0
    16'b11001010_11010101 : OUT <= 0;  //202 / 213 = 0
    16'b11001010_11010110 : OUT <= 0;  //202 / 214 = 0
    16'b11001010_11010111 : OUT <= 0;  //202 / 215 = 0
    16'b11001010_11011000 : OUT <= 0;  //202 / 216 = 0
    16'b11001010_11011001 : OUT <= 0;  //202 / 217 = 0
    16'b11001010_11011010 : OUT <= 0;  //202 / 218 = 0
    16'b11001010_11011011 : OUT <= 0;  //202 / 219 = 0
    16'b11001010_11011100 : OUT <= 0;  //202 / 220 = 0
    16'b11001010_11011101 : OUT <= 0;  //202 / 221 = 0
    16'b11001010_11011110 : OUT <= 0;  //202 / 222 = 0
    16'b11001010_11011111 : OUT <= 0;  //202 / 223 = 0
    16'b11001010_11100000 : OUT <= 0;  //202 / 224 = 0
    16'b11001010_11100001 : OUT <= 0;  //202 / 225 = 0
    16'b11001010_11100010 : OUT <= 0;  //202 / 226 = 0
    16'b11001010_11100011 : OUT <= 0;  //202 / 227 = 0
    16'b11001010_11100100 : OUT <= 0;  //202 / 228 = 0
    16'b11001010_11100101 : OUT <= 0;  //202 / 229 = 0
    16'b11001010_11100110 : OUT <= 0;  //202 / 230 = 0
    16'b11001010_11100111 : OUT <= 0;  //202 / 231 = 0
    16'b11001010_11101000 : OUT <= 0;  //202 / 232 = 0
    16'b11001010_11101001 : OUT <= 0;  //202 / 233 = 0
    16'b11001010_11101010 : OUT <= 0;  //202 / 234 = 0
    16'b11001010_11101011 : OUT <= 0;  //202 / 235 = 0
    16'b11001010_11101100 : OUT <= 0;  //202 / 236 = 0
    16'b11001010_11101101 : OUT <= 0;  //202 / 237 = 0
    16'b11001010_11101110 : OUT <= 0;  //202 / 238 = 0
    16'b11001010_11101111 : OUT <= 0;  //202 / 239 = 0
    16'b11001010_11110000 : OUT <= 0;  //202 / 240 = 0
    16'b11001010_11110001 : OUT <= 0;  //202 / 241 = 0
    16'b11001010_11110010 : OUT <= 0;  //202 / 242 = 0
    16'b11001010_11110011 : OUT <= 0;  //202 / 243 = 0
    16'b11001010_11110100 : OUT <= 0;  //202 / 244 = 0
    16'b11001010_11110101 : OUT <= 0;  //202 / 245 = 0
    16'b11001010_11110110 : OUT <= 0;  //202 / 246 = 0
    16'b11001010_11110111 : OUT <= 0;  //202 / 247 = 0
    16'b11001010_11111000 : OUT <= 0;  //202 / 248 = 0
    16'b11001010_11111001 : OUT <= 0;  //202 / 249 = 0
    16'b11001010_11111010 : OUT <= 0;  //202 / 250 = 0
    16'b11001010_11111011 : OUT <= 0;  //202 / 251 = 0
    16'b11001010_11111100 : OUT <= 0;  //202 / 252 = 0
    16'b11001010_11111101 : OUT <= 0;  //202 / 253 = 0
    16'b11001010_11111110 : OUT <= 0;  //202 / 254 = 0
    16'b11001010_11111111 : OUT <= 0;  //202 / 255 = 0
    16'b11001011_00000000 : OUT <= 0;  //203 / 0 = 0
    16'b11001011_00000001 : OUT <= 203;  //203 / 1 = 203
    16'b11001011_00000010 : OUT <= 101;  //203 / 2 = 101
    16'b11001011_00000011 : OUT <= 67;  //203 / 3 = 67
    16'b11001011_00000100 : OUT <= 50;  //203 / 4 = 50
    16'b11001011_00000101 : OUT <= 40;  //203 / 5 = 40
    16'b11001011_00000110 : OUT <= 33;  //203 / 6 = 33
    16'b11001011_00000111 : OUT <= 29;  //203 / 7 = 29
    16'b11001011_00001000 : OUT <= 25;  //203 / 8 = 25
    16'b11001011_00001001 : OUT <= 22;  //203 / 9 = 22
    16'b11001011_00001010 : OUT <= 20;  //203 / 10 = 20
    16'b11001011_00001011 : OUT <= 18;  //203 / 11 = 18
    16'b11001011_00001100 : OUT <= 16;  //203 / 12 = 16
    16'b11001011_00001101 : OUT <= 15;  //203 / 13 = 15
    16'b11001011_00001110 : OUT <= 14;  //203 / 14 = 14
    16'b11001011_00001111 : OUT <= 13;  //203 / 15 = 13
    16'b11001011_00010000 : OUT <= 12;  //203 / 16 = 12
    16'b11001011_00010001 : OUT <= 11;  //203 / 17 = 11
    16'b11001011_00010010 : OUT <= 11;  //203 / 18 = 11
    16'b11001011_00010011 : OUT <= 10;  //203 / 19 = 10
    16'b11001011_00010100 : OUT <= 10;  //203 / 20 = 10
    16'b11001011_00010101 : OUT <= 9;  //203 / 21 = 9
    16'b11001011_00010110 : OUT <= 9;  //203 / 22 = 9
    16'b11001011_00010111 : OUT <= 8;  //203 / 23 = 8
    16'b11001011_00011000 : OUT <= 8;  //203 / 24 = 8
    16'b11001011_00011001 : OUT <= 8;  //203 / 25 = 8
    16'b11001011_00011010 : OUT <= 7;  //203 / 26 = 7
    16'b11001011_00011011 : OUT <= 7;  //203 / 27 = 7
    16'b11001011_00011100 : OUT <= 7;  //203 / 28 = 7
    16'b11001011_00011101 : OUT <= 7;  //203 / 29 = 7
    16'b11001011_00011110 : OUT <= 6;  //203 / 30 = 6
    16'b11001011_00011111 : OUT <= 6;  //203 / 31 = 6
    16'b11001011_00100000 : OUT <= 6;  //203 / 32 = 6
    16'b11001011_00100001 : OUT <= 6;  //203 / 33 = 6
    16'b11001011_00100010 : OUT <= 5;  //203 / 34 = 5
    16'b11001011_00100011 : OUT <= 5;  //203 / 35 = 5
    16'b11001011_00100100 : OUT <= 5;  //203 / 36 = 5
    16'b11001011_00100101 : OUT <= 5;  //203 / 37 = 5
    16'b11001011_00100110 : OUT <= 5;  //203 / 38 = 5
    16'b11001011_00100111 : OUT <= 5;  //203 / 39 = 5
    16'b11001011_00101000 : OUT <= 5;  //203 / 40 = 5
    16'b11001011_00101001 : OUT <= 4;  //203 / 41 = 4
    16'b11001011_00101010 : OUT <= 4;  //203 / 42 = 4
    16'b11001011_00101011 : OUT <= 4;  //203 / 43 = 4
    16'b11001011_00101100 : OUT <= 4;  //203 / 44 = 4
    16'b11001011_00101101 : OUT <= 4;  //203 / 45 = 4
    16'b11001011_00101110 : OUT <= 4;  //203 / 46 = 4
    16'b11001011_00101111 : OUT <= 4;  //203 / 47 = 4
    16'b11001011_00110000 : OUT <= 4;  //203 / 48 = 4
    16'b11001011_00110001 : OUT <= 4;  //203 / 49 = 4
    16'b11001011_00110010 : OUT <= 4;  //203 / 50 = 4
    16'b11001011_00110011 : OUT <= 3;  //203 / 51 = 3
    16'b11001011_00110100 : OUT <= 3;  //203 / 52 = 3
    16'b11001011_00110101 : OUT <= 3;  //203 / 53 = 3
    16'b11001011_00110110 : OUT <= 3;  //203 / 54 = 3
    16'b11001011_00110111 : OUT <= 3;  //203 / 55 = 3
    16'b11001011_00111000 : OUT <= 3;  //203 / 56 = 3
    16'b11001011_00111001 : OUT <= 3;  //203 / 57 = 3
    16'b11001011_00111010 : OUT <= 3;  //203 / 58 = 3
    16'b11001011_00111011 : OUT <= 3;  //203 / 59 = 3
    16'b11001011_00111100 : OUT <= 3;  //203 / 60 = 3
    16'b11001011_00111101 : OUT <= 3;  //203 / 61 = 3
    16'b11001011_00111110 : OUT <= 3;  //203 / 62 = 3
    16'b11001011_00111111 : OUT <= 3;  //203 / 63 = 3
    16'b11001011_01000000 : OUT <= 3;  //203 / 64 = 3
    16'b11001011_01000001 : OUT <= 3;  //203 / 65 = 3
    16'b11001011_01000010 : OUT <= 3;  //203 / 66 = 3
    16'b11001011_01000011 : OUT <= 3;  //203 / 67 = 3
    16'b11001011_01000100 : OUT <= 2;  //203 / 68 = 2
    16'b11001011_01000101 : OUT <= 2;  //203 / 69 = 2
    16'b11001011_01000110 : OUT <= 2;  //203 / 70 = 2
    16'b11001011_01000111 : OUT <= 2;  //203 / 71 = 2
    16'b11001011_01001000 : OUT <= 2;  //203 / 72 = 2
    16'b11001011_01001001 : OUT <= 2;  //203 / 73 = 2
    16'b11001011_01001010 : OUT <= 2;  //203 / 74 = 2
    16'b11001011_01001011 : OUT <= 2;  //203 / 75 = 2
    16'b11001011_01001100 : OUT <= 2;  //203 / 76 = 2
    16'b11001011_01001101 : OUT <= 2;  //203 / 77 = 2
    16'b11001011_01001110 : OUT <= 2;  //203 / 78 = 2
    16'b11001011_01001111 : OUT <= 2;  //203 / 79 = 2
    16'b11001011_01010000 : OUT <= 2;  //203 / 80 = 2
    16'b11001011_01010001 : OUT <= 2;  //203 / 81 = 2
    16'b11001011_01010010 : OUT <= 2;  //203 / 82 = 2
    16'b11001011_01010011 : OUT <= 2;  //203 / 83 = 2
    16'b11001011_01010100 : OUT <= 2;  //203 / 84 = 2
    16'b11001011_01010101 : OUT <= 2;  //203 / 85 = 2
    16'b11001011_01010110 : OUT <= 2;  //203 / 86 = 2
    16'b11001011_01010111 : OUT <= 2;  //203 / 87 = 2
    16'b11001011_01011000 : OUT <= 2;  //203 / 88 = 2
    16'b11001011_01011001 : OUT <= 2;  //203 / 89 = 2
    16'b11001011_01011010 : OUT <= 2;  //203 / 90 = 2
    16'b11001011_01011011 : OUT <= 2;  //203 / 91 = 2
    16'b11001011_01011100 : OUT <= 2;  //203 / 92 = 2
    16'b11001011_01011101 : OUT <= 2;  //203 / 93 = 2
    16'b11001011_01011110 : OUT <= 2;  //203 / 94 = 2
    16'b11001011_01011111 : OUT <= 2;  //203 / 95 = 2
    16'b11001011_01100000 : OUT <= 2;  //203 / 96 = 2
    16'b11001011_01100001 : OUT <= 2;  //203 / 97 = 2
    16'b11001011_01100010 : OUT <= 2;  //203 / 98 = 2
    16'b11001011_01100011 : OUT <= 2;  //203 / 99 = 2
    16'b11001011_01100100 : OUT <= 2;  //203 / 100 = 2
    16'b11001011_01100101 : OUT <= 2;  //203 / 101 = 2
    16'b11001011_01100110 : OUT <= 1;  //203 / 102 = 1
    16'b11001011_01100111 : OUT <= 1;  //203 / 103 = 1
    16'b11001011_01101000 : OUT <= 1;  //203 / 104 = 1
    16'b11001011_01101001 : OUT <= 1;  //203 / 105 = 1
    16'b11001011_01101010 : OUT <= 1;  //203 / 106 = 1
    16'b11001011_01101011 : OUT <= 1;  //203 / 107 = 1
    16'b11001011_01101100 : OUT <= 1;  //203 / 108 = 1
    16'b11001011_01101101 : OUT <= 1;  //203 / 109 = 1
    16'b11001011_01101110 : OUT <= 1;  //203 / 110 = 1
    16'b11001011_01101111 : OUT <= 1;  //203 / 111 = 1
    16'b11001011_01110000 : OUT <= 1;  //203 / 112 = 1
    16'b11001011_01110001 : OUT <= 1;  //203 / 113 = 1
    16'b11001011_01110010 : OUT <= 1;  //203 / 114 = 1
    16'b11001011_01110011 : OUT <= 1;  //203 / 115 = 1
    16'b11001011_01110100 : OUT <= 1;  //203 / 116 = 1
    16'b11001011_01110101 : OUT <= 1;  //203 / 117 = 1
    16'b11001011_01110110 : OUT <= 1;  //203 / 118 = 1
    16'b11001011_01110111 : OUT <= 1;  //203 / 119 = 1
    16'b11001011_01111000 : OUT <= 1;  //203 / 120 = 1
    16'b11001011_01111001 : OUT <= 1;  //203 / 121 = 1
    16'b11001011_01111010 : OUT <= 1;  //203 / 122 = 1
    16'b11001011_01111011 : OUT <= 1;  //203 / 123 = 1
    16'b11001011_01111100 : OUT <= 1;  //203 / 124 = 1
    16'b11001011_01111101 : OUT <= 1;  //203 / 125 = 1
    16'b11001011_01111110 : OUT <= 1;  //203 / 126 = 1
    16'b11001011_01111111 : OUT <= 1;  //203 / 127 = 1
    16'b11001011_10000000 : OUT <= 1;  //203 / 128 = 1
    16'b11001011_10000001 : OUT <= 1;  //203 / 129 = 1
    16'b11001011_10000010 : OUT <= 1;  //203 / 130 = 1
    16'b11001011_10000011 : OUT <= 1;  //203 / 131 = 1
    16'b11001011_10000100 : OUT <= 1;  //203 / 132 = 1
    16'b11001011_10000101 : OUT <= 1;  //203 / 133 = 1
    16'b11001011_10000110 : OUT <= 1;  //203 / 134 = 1
    16'b11001011_10000111 : OUT <= 1;  //203 / 135 = 1
    16'b11001011_10001000 : OUT <= 1;  //203 / 136 = 1
    16'b11001011_10001001 : OUT <= 1;  //203 / 137 = 1
    16'b11001011_10001010 : OUT <= 1;  //203 / 138 = 1
    16'b11001011_10001011 : OUT <= 1;  //203 / 139 = 1
    16'b11001011_10001100 : OUT <= 1;  //203 / 140 = 1
    16'b11001011_10001101 : OUT <= 1;  //203 / 141 = 1
    16'b11001011_10001110 : OUT <= 1;  //203 / 142 = 1
    16'b11001011_10001111 : OUT <= 1;  //203 / 143 = 1
    16'b11001011_10010000 : OUT <= 1;  //203 / 144 = 1
    16'b11001011_10010001 : OUT <= 1;  //203 / 145 = 1
    16'b11001011_10010010 : OUT <= 1;  //203 / 146 = 1
    16'b11001011_10010011 : OUT <= 1;  //203 / 147 = 1
    16'b11001011_10010100 : OUT <= 1;  //203 / 148 = 1
    16'b11001011_10010101 : OUT <= 1;  //203 / 149 = 1
    16'b11001011_10010110 : OUT <= 1;  //203 / 150 = 1
    16'b11001011_10010111 : OUT <= 1;  //203 / 151 = 1
    16'b11001011_10011000 : OUT <= 1;  //203 / 152 = 1
    16'b11001011_10011001 : OUT <= 1;  //203 / 153 = 1
    16'b11001011_10011010 : OUT <= 1;  //203 / 154 = 1
    16'b11001011_10011011 : OUT <= 1;  //203 / 155 = 1
    16'b11001011_10011100 : OUT <= 1;  //203 / 156 = 1
    16'b11001011_10011101 : OUT <= 1;  //203 / 157 = 1
    16'b11001011_10011110 : OUT <= 1;  //203 / 158 = 1
    16'b11001011_10011111 : OUT <= 1;  //203 / 159 = 1
    16'b11001011_10100000 : OUT <= 1;  //203 / 160 = 1
    16'b11001011_10100001 : OUT <= 1;  //203 / 161 = 1
    16'b11001011_10100010 : OUT <= 1;  //203 / 162 = 1
    16'b11001011_10100011 : OUT <= 1;  //203 / 163 = 1
    16'b11001011_10100100 : OUT <= 1;  //203 / 164 = 1
    16'b11001011_10100101 : OUT <= 1;  //203 / 165 = 1
    16'b11001011_10100110 : OUT <= 1;  //203 / 166 = 1
    16'b11001011_10100111 : OUT <= 1;  //203 / 167 = 1
    16'b11001011_10101000 : OUT <= 1;  //203 / 168 = 1
    16'b11001011_10101001 : OUT <= 1;  //203 / 169 = 1
    16'b11001011_10101010 : OUT <= 1;  //203 / 170 = 1
    16'b11001011_10101011 : OUT <= 1;  //203 / 171 = 1
    16'b11001011_10101100 : OUT <= 1;  //203 / 172 = 1
    16'b11001011_10101101 : OUT <= 1;  //203 / 173 = 1
    16'b11001011_10101110 : OUT <= 1;  //203 / 174 = 1
    16'b11001011_10101111 : OUT <= 1;  //203 / 175 = 1
    16'b11001011_10110000 : OUT <= 1;  //203 / 176 = 1
    16'b11001011_10110001 : OUT <= 1;  //203 / 177 = 1
    16'b11001011_10110010 : OUT <= 1;  //203 / 178 = 1
    16'b11001011_10110011 : OUT <= 1;  //203 / 179 = 1
    16'b11001011_10110100 : OUT <= 1;  //203 / 180 = 1
    16'b11001011_10110101 : OUT <= 1;  //203 / 181 = 1
    16'b11001011_10110110 : OUT <= 1;  //203 / 182 = 1
    16'b11001011_10110111 : OUT <= 1;  //203 / 183 = 1
    16'b11001011_10111000 : OUT <= 1;  //203 / 184 = 1
    16'b11001011_10111001 : OUT <= 1;  //203 / 185 = 1
    16'b11001011_10111010 : OUT <= 1;  //203 / 186 = 1
    16'b11001011_10111011 : OUT <= 1;  //203 / 187 = 1
    16'b11001011_10111100 : OUT <= 1;  //203 / 188 = 1
    16'b11001011_10111101 : OUT <= 1;  //203 / 189 = 1
    16'b11001011_10111110 : OUT <= 1;  //203 / 190 = 1
    16'b11001011_10111111 : OUT <= 1;  //203 / 191 = 1
    16'b11001011_11000000 : OUT <= 1;  //203 / 192 = 1
    16'b11001011_11000001 : OUT <= 1;  //203 / 193 = 1
    16'b11001011_11000010 : OUT <= 1;  //203 / 194 = 1
    16'b11001011_11000011 : OUT <= 1;  //203 / 195 = 1
    16'b11001011_11000100 : OUT <= 1;  //203 / 196 = 1
    16'b11001011_11000101 : OUT <= 1;  //203 / 197 = 1
    16'b11001011_11000110 : OUT <= 1;  //203 / 198 = 1
    16'b11001011_11000111 : OUT <= 1;  //203 / 199 = 1
    16'b11001011_11001000 : OUT <= 1;  //203 / 200 = 1
    16'b11001011_11001001 : OUT <= 1;  //203 / 201 = 1
    16'b11001011_11001010 : OUT <= 1;  //203 / 202 = 1
    16'b11001011_11001011 : OUT <= 1;  //203 / 203 = 1
    16'b11001011_11001100 : OUT <= 0;  //203 / 204 = 0
    16'b11001011_11001101 : OUT <= 0;  //203 / 205 = 0
    16'b11001011_11001110 : OUT <= 0;  //203 / 206 = 0
    16'b11001011_11001111 : OUT <= 0;  //203 / 207 = 0
    16'b11001011_11010000 : OUT <= 0;  //203 / 208 = 0
    16'b11001011_11010001 : OUT <= 0;  //203 / 209 = 0
    16'b11001011_11010010 : OUT <= 0;  //203 / 210 = 0
    16'b11001011_11010011 : OUT <= 0;  //203 / 211 = 0
    16'b11001011_11010100 : OUT <= 0;  //203 / 212 = 0
    16'b11001011_11010101 : OUT <= 0;  //203 / 213 = 0
    16'b11001011_11010110 : OUT <= 0;  //203 / 214 = 0
    16'b11001011_11010111 : OUT <= 0;  //203 / 215 = 0
    16'b11001011_11011000 : OUT <= 0;  //203 / 216 = 0
    16'b11001011_11011001 : OUT <= 0;  //203 / 217 = 0
    16'b11001011_11011010 : OUT <= 0;  //203 / 218 = 0
    16'b11001011_11011011 : OUT <= 0;  //203 / 219 = 0
    16'b11001011_11011100 : OUT <= 0;  //203 / 220 = 0
    16'b11001011_11011101 : OUT <= 0;  //203 / 221 = 0
    16'b11001011_11011110 : OUT <= 0;  //203 / 222 = 0
    16'b11001011_11011111 : OUT <= 0;  //203 / 223 = 0
    16'b11001011_11100000 : OUT <= 0;  //203 / 224 = 0
    16'b11001011_11100001 : OUT <= 0;  //203 / 225 = 0
    16'b11001011_11100010 : OUT <= 0;  //203 / 226 = 0
    16'b11001011_11100011 : OUT <= 0;  //203 / 227 = 0
    16'b11001011_11100100 : OUT <= 0;  //203 / 228 = 0
    16'b11001011_11100101 : OUT <= 0;  //203 / 229 = 0
    16'b11001011_11100110 : OUT <= 0;  //203 / 230 = 0
    16'b11001011_11100111 : OUT <= 0;  //203 / 231 = 0
    16'b11001011_11101000 : OUT <= 0;  //203 / 232 = 0
    16'b11001011_11101001 : OUT <= 0;  //203 / 233 = 0
    16'b11001011_11101010 : OUT <= 0;  //203 / 234 = 0
    16'b11001011_11101011 : OUT <= 0;  //203 / 235 = 0
    16'b11001011_11101100 : OUT <= 0;  //203 / 236 = 0
    16'b11001011_11101101 : OUT <= 0;  //203 / 237 = 0
    16'b11001011_11101110 : OUT <= 0;  //203 / 238 = 0
    16'b11001011_11101111 : OUT <= 0;  //203 / 239 = 0
    16'b11001011_11110000 : OUT <= 0;  //203 / 240 = 0
    16'b11001011_11110001 : OUT <= 0;  //203 / 241 = 0
    16'b11001011_11110010 : OUT <= 0;  //203 / 242 = 0
    16'b11001011_11110011 : OUT <= 0;  //203 / 243 = 0
    16'b11001011_11110100 : OUT <= 0;  //203 / 244 = 0
    16'b11001011_11110101 : OUT <= 0;  //203 / 245 = 0
    16'b11001011_11110110 : OUT <= 0;  //203 / 246 = 0
    16'b11001011_11110111 : OUT <= 0;  //203 / 247 = 0
    16'b11001011_11111000 : OUT <= 0;  //203 / 248 = 0
    16'b11001011_11111001 : OUT <= 0;  //203 / 249 = 0
    16'b11001011_11111010 : OUT <= 0;  //203 / 250 = 0
    16'b11001011_11111011 : OUT <= 0;  //203 / 251 = 0
    16'b11001011_11111100 : OUT <= 0;  //203 / 252 = 0
    16'b11001011_11111101 : OUT <= 0;  //203 / 253 = 0
    16'b11001011_11111110 : OUT <= 0;  //203 / 254 = 0
    16'b11001011_11111111 : OUT <= 0;  //203 / 255 = 0
    16'b11001100_00000000 : OUT <= 0;  //204 / 0 = 0
    16'b11001100_00000001 : OUT <= 204;  //204 / 1 = 204
    16'b11001100_00000010 : OUT <= 102;  //204 / 2 = 102
    16'b11001100_00000011 : OUT <= 68;  //204 / 3 = 68
    16'b11001100_00000100 : OUT <= 51;  //204 / 4 = 51
    16'b11001100_00000101 : OUT <= 40;  //204 / 5 = 40
    16'b11001100_00000110 : OUT <= 34;  //204 / 6 = 34
    16'b11001100_00000111 : OUT <= 29;  //204 / 7 = 29
    16'b11001100_00001000 : OUT <= 25;  //204 / 8 = 25
    16'b11001100_00001001 : OUT <= 22;  //204 / 9 = 22
    16'b11001100_00001010 : OUT <= 20;  //204 / 10 = 20
    16'b11001100_00001011 : OUT <= 18;  //204 / 11 = 18
    16'b11001100_00001100 : OUT <= 17;  //204 / 12 = 17
    16'b11001100_00001101 : OUT <= 15;  //204 / 13 = 15
    16'b11001100_00001110 : OUT <= 14;  //204 / 14 = 14
    16'b11001100_00001111 : OUT <= 13;  //204 / 15 = 13
    16'b11001100_00010000 : OUT <= 12;  //204 / 16 = 12
    16'b11001100_00010001 : OUT <= 12;  //204 / 17 = 12
    16'b11001100_00010010 : OUT <= 11;  //204 / 18 = 11
    16'b11001100_00010011 : OUT <= 10;  //204 / 19 = 10
    16'b11001100_00010100 : OUT <= 10;  //204 / 20 = 10
    16'b11001100_00010101 : OUT <= 9;  //204 / 21 = 9
    16'b11001100_00010110 : OUT <= 9;  //204 / 22 = 9
    16'b11001100_00010111 : OUT <= 8;  //204 / 23 = 8
    16'b11001100_00011000 : OUT <= 8;  //204 / 24 = 8
    16'b11001100_00011001 : OUT <= 8;  //204 / 25 = 8
    16'b11001100_00011010 : OUT <= 7;  //204 / 26 = 7
    16'b11001100_00011011 : OUT <= 7;  //204 / 27 = 7
    16'b11001100_00011100 : OUT <= 7;  //204 / 28 = 7
    16'b11001100_00011101 : OUT <= 7;  //204 / 29 = 7
    16'b11001100_00011110 : OUT <= 6;  //204 / 30 = 6
    16'b11001100_00011111 : OUT <= 6;  //204 / 31 = 6
    16'b11001100_00100000 : OUT <= 6;  //204 / 32 = 6
    16'b11001100_00100001 : OUT <= 6;  //204 / 33 = 6
    16'b11001100_00100010 : OUT <= 6;  //204 / 34 = 6
    16'b11001100_00100011 : OUT <= 5;  //204 / 35 = 5
    16'b11001100_00100100 : OUT <= 5;  //204 / 36 = 5
    16'b11001100_00100101 : OUT <= 5;  //204 / 37 = 5
    16'b11001100_00100110 : OUT <= 5;  //204 / 38 = 5
    16'b11001100_00100111 : OUT <= 5;  //204 / 39 = 5
    16'b11001100_00101000 : OUT <= 5;  //204 / 40 = 5
    16'b11001100_00101001 : OUT <= 4;  //204 / 41 = 4
    16'b11001100_00101010 : OUT <= 4;  //204 / 42 = 4
    16'b11001100_00101011 : OUT <= 4;  //204 / 43 = 4
    16'b11001100_00101100 : OUT <= 4;  //204 / 44 = 4
    16'b11001100_00101101 : OUT <= 4;  //204 / 45 = 4
    16'b11001100_00101110 : OUT <= 4;  //204 / 46 = 4
    16'b11001100_00101111 : OUT <= 4;  //204 / 47 = 4
    16'b11001100_00110000 : OUT <= 4;  //204 / 48 = 4
    16'b11001100_00110001 : OUT <= 4;  //204 / 49 = 4
    16'b11001100_00110010 : OUT <= 4;  //204 / 50 = 4
    16'b11001100_00110011 : OUT <= 4;  //204 / 51 = 4
    16'b11001100_00110100 : OUT <= 3;  //204 / 52 = 3
    16'b11001100_00110101 : OUT <= 3;  //204 / 53 = 3
    16'b11001100_00110110 : OUT <= 3;  //204 / 54 = 3
    16'b11001100_00110111 : OUT <= 3;  //204 / 55 = 3
    16'b11001100_00111000 : OUT <= 3;  //204 / 56 = 3
    16'b11001100_00111001 : OUT <= 3;  //204 / 57 = 3
    16'b11001100_00111010 : OUT <= 3;  //204 / 58 = 3
    16'b11001100_00111011 : OUT <= 3;  //204 / 59 = 3
    16'b11001100_00111100 : OUT <= 3;  //204 / 60 = 3
    16'b11001100_00111101 : OUT <= 3;  //204 / 61 = 3
    16'b11001100_00111110 : OUT <= 3;  //204 / 62 = 3
    16'b11001100_00111111 : OUT <= 3;  //204 / 63 = 3
    16'b11001100_01000000 : OUT <= 3;  //204 / 64 = 3
    16'b11001100_01000001 : OUT <= 3;  //204 / 65 = 3
    16'b11001100_01000010 : OUT <= 3;  //204 / 66 = 3
    16'b11001100_01000011 : OUT <= 3;  //204 / 67 = 3
    16'b11001100_01000100 : OUT <= 3;  //204 / 68 = 3
    16'b11001100_01000101 : OUT <= 2;  //204 / 69 = 2
    16'b11001100_01000110 : OUT <= 2;  //204 / 70 = 2
    16'b11001100_01000111 : OUT <= 2;  //204 / 71 = 2
    16'b11001100_01001000 : OUT <= 2;  //204 / 72 = 2
    16'b11001100_01001001 : OUT <= 2;  //204 / 73 = 2
    16'b11001100_01001010 : OUT <= 2;  //204 / 74 = 2
    16'b11001100_01001011 : OUT <= 2;  //204 / 75 = 2
    16'b11001100_01001100 : OUT <= 2;  //204 / 76 = 2
    16'b11001100_01001101 : OUT <= 2;  //204 / 77 = 2
    16'b11001100_01001110 : OUT <= 2;  //204 / 78 = 2
    16'b11001100_01001111 : OUT <= 2;  //204 / 79 = 2
    16'b11001100_01010000 : OUT <= 2;  //204 / 80 = 2
    16'b11001100_01010001 : OUT <= 2;  //204 / 81 = 2
    16'b11001100_01010010 : OUT <= 2;  //204 / 82 = 2
    16'b11001100_01010011 : OUT <= 2;  //204 / 83 = 2
    16'b11001100_01010100 : OUT <= 2;  //204 / 84 = 2
    16'b11001100_01010101 : OUT <= 2;  //204 / 85 = 2
    16'b11001100_01010110 : OUT <= 2;  //204 / 86 = 2
    16'b11001100_01010111 : OUT <= 2;  //204 / 87 = 2
    16'b11001100_01011000 : OUT <= 2;  //204 / 88 = 2
    16'b11001100_01011001 : OUT <= 2;  //204 / 89 = 2
    16'b11001100_01011010 : OUT <= 2;  //204 / 90 = 2
    16'b11001100_01011011 : OUT <= 2;  //204 / 91 = 2
    16'b11001100_01011100 : OUT <= 2;  //204 / 92 = 2
    16'b11001100_01011101 : OUT <= 2;  //204 / 93 = 2
    16'b11001100_01011110 : OUT <= 2;  //204 / 94 = 2
    16'b11001100_01011111 : OUT <= 2;  //204 / 95 = 2
    16'b11001100_01100000 : OUT <= 2;  //204 / 96 = 2
    16'b11001100_01100001 : OUT <= 2;  //204 / 97 = 2
    16'b11001100_01100010 : OUT <= 2;  //204 / 98 = 2
    16'b11001100_01100011 : OUT <= 2;  //204 / 99 = 2
    16'b11001100_01100100 : OUT <= 2;  //204 / 100 = 2
    16'b11001100_01100101 : OUT <= 2;  //204 / 101 = 2
    16'b11001100_01100110 : OUT <= 2;  //204 / 102 = 2
    16'b11001100_01100111 : OUT <= 1;  //204 / 103 = 1
    16'b11001100_01101000 : OUT <= 1;  //204 / 104 = 1
    16'b11001100_01101001 : OUT <= 1;  //204 / 105 = 1
    16'b11001100_01101010 : OUT <= 1;  //204 / 106 = 1
    16'b11001100_01101011 : OUT <= 1;  //204 / 107 = 1
    16'b11001100_01101100 : OUT <= 1;  //204 / 108 = 1
    16'b11001100_01101101 : OUT <= 1;  //204 / 109 = 1
    16'b11001100_01101110 : OUT <= 1;  //204 / 110 = 1
    16'b11001100_01101111 : OUT <= 1;  //204 / 111 = 1
    16'b11001100_01110000 : OUT <= 1;  //204 / 112 = 1
    16'b11001100_01110001 : OUT <= 1;  //204 / 113 = 1
    16'b11001100_01110010 : OUT <= 1;  //204 / 114 = 1
    16'b11001100_01110011 : OUT <= 1;  //204 / 115 = 1
    16'b11001100_01110100 : OUT <= 1;  //204 / 116 = 1
    16'b11001100_01110101 : OUT <= 1;  //204 / 117 = 1
    16'b11001100_01110110 : OUT <= 1;  //204 / 118 = 1
    16'b11001100_01110111 : OUT <= 1;  //204 / 119 = 1
    16'b11001100_01111000 : OUT <= 1;  //204 / 120 = 1
    16'b11001100_01111001 : OUT <= 1;  //204 / 121 = 1
    16'b11001100_01111010 : OUT <= 1;  //204 / 122 = 1
    16'b11001100_01111011 : OUT <= 1;  //204 / 123 = 1
    16'b11001100_01111100 : OUT <= 1;  //204 / 124 = 1
    16'b11001100_01111101 : OUT <= 1;  //204 / 125 = 1
    16'b11001100_01111110 : OUT <= 1;  //204 / 126 = 1
    16'b11001100_01111111 : OUT <= 1;  //204 / 127 = 1
    16'b11001100_10000000 : OUT <= 1;  //204 / 128 = 1
    16'b11001100_10000001 : OUT <= 1;  //204 / 129 = 1
    16'b11001100_10000010 : OUT <= 1;  //204 / 130 = 1
    16'b11001100_10000011 : OUT <= 1;  //204 / 131 = 1
    16'b11001100_10000100 : OUT <= 1;  //204 / 132 = 1
    16'b11001100_10000101 : OUT <= 1;  //204 / 133 = 1
    16'b11001100_10000110 : OUT <= 1;  //204 / 134 = 1
    16'b11001100_10000111 : OUT <= 1;  //204 / 135 = 1
    16'b11001100_10001000 : OUT <= 1;  //204 / 136 = 1
    16'b11001100_10001001 : OUT <= 1;  //204 / 137 = 1
    16'b11001100_10001010 : OUT <= 1;  //204 / 138 = 1
    16'b11001100_10001011 : OUT <= 1;  //204 / 139 = 1
    16'b11001100_10001100 : OUT <= 1;  //204 / 140 = 1
    16'b11001100_10001101 : OUT <= 1;  //204 / 141 = 1
    16'b11001100_10001110 : OUT <= 1;  //204 / 142 = 1
    16'b11001100_10001111 : OUT <= 1;  //204 / 143 = 1
    16'b11001100_10010000 : OUT <= 1;  //204 / 144 = 1
    16'b11001100_10010001 : OUT <= 1;  //204 / 145 = 1
    16'b11001100_10010010 : OUT <= 1;  //204 / 146 = 1
    16'b11001100_10010011 : OUT <= 1;  //204 / 147 = 1
    16'b11001100_10010100 : OUT <= 1;  //204 / 148 = 1
    16'b11001100_10010101 : OUT <= 1;  //204 / 149 = 1
    16'b11001100_10010110 : OUT <= 1;  //204 / 150 = 1
    16'b11001100_10010111 : OUT <= 1;  //204 / 151 = 1
    16'b11001100_10011000 : OUT <= 1;  //204 / 152 = 1
    16'b11001100_10011001 : OUT <= 1;  //204 / 153 = 1
    16'b11001100_10011010 : OUT <= 1;  //204 / 154 = 1
    16'b11001100_10011011 : OUT <= 1;  //204 / 155 = 1
    16'b11001100_10011100 : OUT <= 1;  //204 / 156 = 1
    16'b11001100_10011101 : OUT <= 1;  //204 / 157 = 1
    16'b11001100_10011110 : OUT <= 1;  //204 / 158 = 1
    16'b11001100_10011111 : OUT <= 1;  //204 / 159 = 1
    16'b11001100_10100000 : OUT <= 1;  //204 / 160 = 1
    16'b11001100_10100001 : OUT <= 1;  //204 / 161 = 1
    16'b11001100_10100010 : OUT <= 1;  //204 / 162 = 1
    16'b11001100_10100011 : OUT <= 1;  //204 / 163 = 1
    16'b11001100_10100100 : OUT <= 1;  //204 / 164 = 1
    16'b11001100_10100101 : OUT <= 1;  //204 / 165 = 1
    16'b11001100_10100110 : OUT <= 1;  //204 / 166 = 1
    16'b11001100_10100111 : OUT <= 1;  //204 / 167 = 1
    16'b11001100_10101000 : OUT <= 1;  //204 / 168 = 1
    16'b11001100_10101001 : OUT <= 1;  //204 / 169 = 1
    16'b11001100_10101010 : OUT <= 1;  //204 / 170 = 1
    16'b11001100_10101011 : OUT <= 1;  //204 / 171 = 1
    16'b11001100_10101100 : OUT <= 1;  //204 / 172 = 1
    16'b11001100_10101101 : OUT <= 1;  //204 / 173 = 1
    16'b11001100_10101110 : OUT <= 1;  //204 / 174 = 1
    16'b11001100_10101111 : OUT <= 1;  //204 / 175 = 1
    16'b11001100_10110000 : OUT <= 1;  //204 / 176 = 1
    16'b11001100_10110001 : OUT <= 1;  //204 / 177 = 1
    16'b11001100_10110010 : OUT <= 1;  //204 / 178 = 1
    16'b11001100_10110011 : OUT <= 1;  //204 / 179 = 1
    16'b11001100_10110100 : OUT <= 1;  //204 / 180 = 1
    16'b11001100_10110101 : OUT <= 1;  //204 / 181 = 1
    16'b11001100_10110110 : OUT <= 1;  //204 / 182 = 1
    16'b11001100_10110111 : OUT <= 1;  //204 / 183 = 1
    16'b11001100_10111000 : OUT <= 1;  //204 / 184 = 1
    16'b11001100_10111001 : OUT <= 1;  //204 / 185 = 1
    16'b11001100_10111010 : OUT <= 1;  //204 / 186 = 1
    16'b11001100_10111011 : OUT <= 1;  //204 / 187 = 1
    16'b11001100_10111100 : OUT <= 1;  //204 / 188 = 1
    16'b11001100_10111101 : OUT <= 1;  //204 / 189 = 1
    16'b11001100_10111110 : OUT <= 1;  //204 / 190 = 1
    16'b11001100_10111111 : OUT <= 1;  //204 / 191 = 1
    16'b11001100_11000000 : OUT <= 1;  //204 / 192 = 1
    16'b11001100_11000001 : OUT <= 1;  //204 / 193 = 1
    16'b11001100_11000010 : OUT <= 1;  //204 / 194 = 1
    16'b11001100_11000011 : OUT <= 1;  //204 / 195 = 1
    16'b11001100_11000100 : OUT <= 1;  //204 / 196 = 1
    16'b11001100_11000101 : OUT <= 1;  //204 / 197 = 1
    16'b11001100_11000110 : OUT <= 1;  //204 / 198 = 1
    16'b11001100_11000111 : OUT <= 1;  //204 / 199 = 1
    16'b11001100_11001000 : OUT <= 1;  //204 / 200 = 1
    16'b11001100_11001001 : OUT <= 1;  //204 / 201 = 1
    16'b11001100_11001010 : OUT <= 1;  //204 / 202 = 1
    16'b11001100_11001011 : OUT <= 1;  //204 / 203 = 1
    16'b11001100_11001100 : OUT <= 1;  //204 / 204 = 1
    16'b11001100_11001101 : OUT <= 0;  //204 / 205 = 0
    16'b11001100_11001110 : OUT <= 0;  //204 / 206 = 0
    16'b11001100_11001111 : OUT <= 0;  //204 / 207 = 0
    16'b11001100_11010000 : OUT <= 0;  //204 / 208 = 0
    16'b11001100_11010001 : OUT <= 0;  //204 / 209 = 0
    16'b11001100_11010010 : OUT <= 0;  //204 / 210 = 0
    16'b11001100_11010011 : OUT <= 0;  //204 / 211 = 0
    16'b11001100_11010100 : OUT <= 0;  //204 / 212 = 0
    16'b11001100_11010101 : OUT <= 0;  //204 / 213 = 0
    16'b11001100_11010110 : OUT <= 0;  //204 / 214 = 0
    16'b11001100_11010111 : OUT <= 0;  //204 / 215 = 0
    16'b11001100_11011000 : OUT <= 0;  //204 / 216 = 0
    16'b11001100_11011001 : OUT <= 0;  //204 / 217 = 0
    16'b11001100_11011010 : OUT <= 0;  //204 / 218 = 0
    16'b11001100_11011011 : OUT <= 0;  //204 / 219 = 0
    16'b11001100_11011100 : OUT <= 0;  //204 / 220 = 0
    16'b11001100_11011101 : OUT <= 0;  //204 / 221 = 0
    16'b11001100_11011110 : OUT <= 0;  //204 / 222 = 0
    16'b11001100_11011111 : OUT <= 0;  //204 / 223 = 0
    16'b11001100_11100000 : OUT <= 0;  //204 / 224 = 0
    16'b11001100_11100001 : OUT <= 0;  //204 / 225 = 0
    16'b11001100_11100010 : OUT <= 0;  //204 / 226 = 0
    16'b11001100_11100011 : OUT <= 0;  //204 / 227 = 0
    16'b11001100_11100100 : OUT <= 0;  //204 / 228 = 0
    16'b11001100_11100101 : OUT <= 0;  //204 / 229 = 0
    16'b11001100_11100110 : OUT <= 0;  //204 / 230 = 0
    16'b11001100_11100111 : OUT <= 0;  //204 / 231 = 0
    16'b11001100_11101000 : OUT <= 0;  //204 / 232 = 0
    16'b11001100_11101001 : OUT <= 0;  //204 / 233 = 0
    16'b11001100_11101010 : OUT <= 0;  //204 / 234 = 0
    16'b11001100_11101011 : OUT <= 0;  //204 / 235 = 0
    16'b11001100_11101100 : OUT <= 0;  //204 / 236 = 0
    16'b11001100_11101101 : OUT <= 0;  //204 / 237 = 0
    16'b11001100_11101110 : OUT <= 0;  //204 / 238 = 0
    16'b11001100_11101111 : OUT <= 0;  //204 / 239 = 0
    16'b11001100_11110000 : OUT <= 0;  //204 / 240 = 0
    16'b11001100_11110001 : OUT <= 0;  //204 / 241 = 0
    16'b11001100_11110010 : OUT <= 0;  //204 / 242 = 0
    16'b11001100_11110011 : OUT <= 0;  //204 / 243 = 0
    16'b11001100_11110100 : OUT <= 0;  //204 / 244 = 0
    16'b11001100_11110101 : OUT <= 0;  //204 / 245 = 0
    16'b11001100_11110110 : OUT <= 0;  //204 / 246 = 0
    16'b11001100_11110111 : OUT <= 0;  //204 / 247 = 0
    16'b11001100_11111000 : OUT <= 0;  //204 / 248 = 0
    16'b11001100_11111001 : OUT <= 0;  //204 / 249 = 0
    16'b11001100_11111010 : OUT <= 0;  //204 / 250 = 0
    16'b11001100_11111011 : OUT <= 0;  //204 / 251 = 0
    16'b11001100_11111100 : OUT <= 0;  //204 / 252 = 0
    16'b11001100_11111101 : OUT <= 0;  //204 / 253 = 0
    16'b11001100_11111110 : OUT <= 0;  //204 / 254 = 0
    16'b11001100_11111111 : OUT <= 0;  //204 / 255 = 0
    16'b11001101_00000000 : OUT <= 0;  //205 / 0 = 0
    16'b11001101_00000001 : OUT <= 205;  //205 / 1 = 205
    16'b11001101_00000010 : OUT <= 102;  //205 / 2 = 102
    16'b11001101_00000011 : OUT <= 68;  //205 / 3 = 68
    16'b11001101_00000100 : OUT <= 51;  //205 / 4 = 51
    16'b11001101_00000101 : OUT <= 41;  //205 / 5 = 41
    16'b11001101_00000110 : OUT <= 34;  //205 / 6 = 34
    16'b11001101_00000111 : OUT <= 29;  //205 / 7 = 29
    16'b11001101_00001000 : OUT <= 25;  //205 / 8 = 25
    16'b11001101_00001001 : OUT <= 22;  //205 / 9 = 22
    16'b11001101_00001010 : OUT <= 20;  //205 / 10 = 20
    16'b11001101_00001011 : OUT <= 18;  //205 / 11 = 18
    16'b11001101_00001100 : OUT <= 17;  //205 / 12 = 17
    16'b11001101_00001101 : OUT <= 15;  //205 / 13 = 15
    16'b11001101_00001110 : OUT <= 14;  //205 / 14 = 14
    16'b11001101_00001111 : OUT <= 13;  //205 / 15 = 13
    16'b11001101_00010000 : OUT <= 12;  //205 / 16 = 12
    16'b11001101_00010001 : OUT <= 12;  //205 / 17 = 12
    16'b11001101_00010010 : OUT <= 11;  //205 / 18 = 11
    16'b11001101_00010011 : OUT <= 10;  //205 / 19 = 10
    16'b11001101_00010100 : OUT <= 10;  //205 / 20 = 10
    16'b11001101_00010101 : OUT <= 9;  //205 / 21 = 9
    16'b11001101_00010110 : OUT <= 9;  //205 / 22 = 9
    16'b11001101_00010111 : OUT <= 8;  //205 / 23 = 8
    16'b11001101_00011000 : OUT <= 8;  //205 / 24 = 8
    16'b11001101_00011001 : OUT <= 8;  //205 / 25 = 8
    16'b11001101_00011010 : OUT <= 7;  //205 / 26 = 7
    16'b11001101_00011011 : OUT <= 7;  //205 / 27 = 7
    16'b11001101_00011100 : OUT <= 7;  //205 / 28 = 7
    16'b11001101_00011101 : OUT <= 7;  //205 / 29 = 7
    16'b11001101_00011110 : OUT <= 6;  //205 / 30 = 6
    16'b11001101_00011111 : OUT <= 6;  //205 / 31 = 6
    16'b11001101_00100000 : OUT <= 6;  //205 / 32 = 6
    16'b11001101_00100001 : OUT <= 6;  //205 / 33 = 6
    16'b11001101_00100010 : OUT <= 6;  //205 / 34 = 6
    16'b11001101_00100011 : OUT <= 5;  //205 / 35 = 5
    16'b11001101_00100100 : OUT <= 5;  //205 / 36 = 5
    16'b11001101_00100101 : OUT <= 5;  //205 / 37 = 5
    16'b11001101_00100110 : OUT <= 5;  //205 / 38 = 5
    16'b11001101_00100111 : OUT <= 5;  //205 / 39 = 5
    16'b11001101_00101000 : OUT <= 5;  //205 / 40 = 5
    16'b11001101_00101001 : OUT <= 5;  //205 / 41 = 5
    16'b11001101_00101010 : OUT <= 4;  //205 / 42 = 4
    16'b11001101_00101011 : OUT <= 4;  //205 / 43 = 4
    16'b11001101_00101100 : OUT <= 4;  //205 / 44 = 4
    16'b11001101_00101101 : OUT <= 4;  //205 / 45 = 4
    16'b11001101_00101110 : OUT <= 4;  //205 / 46 = 4
    16'b11001101_00101111 : OUT <= 4;  //205 / 47 = 4
    16'b11001101_00110000 : OUT <= 4;  //205 / 48 = 4
    16'b11001101_00110001 : OUT <= 4;  //205 / 49 = 4
    16'b11001101_00110010 : OUT <= 4;  //205 / 50 = 4
    16'b11001101_00110011 : OUT <= 4;  //205 / 51 = 4
    16'b11001101_00110100 : OUT <= 3;  //205 / 52 = 3
    16'b11001101_00110101 : OUT <= 3;  //205 / 53 = 3
    16'b11001101_00110110 : OUT <= 3;  //205 / 54 = 3
    16'b11001101_00110111 : OUT <= 3;  //205 / 55 = 3
    16'b11001101_00111000 : OUT <= 3;  //205 / 56 = 3
    16'b11001101_00111001 : OUT <= 3;  //205 / 57 = 3
    16'b11001101_00111010 : OUT <= 3;  //205 / 58 = 3
    16'b11001101_00111011 : OUT <= 3;  //205 / 59 = 3
    16'b11001101_00111100 : OUT <= 3;  //205 / 60 = 3
    16'b11001101_00111101 : OUT <= 3;  //205 / 61 = 3
    16'b11001101_00111110 : OUT <= 3;  //205 / 62 = 3
    16'b11001101_00111111 : OUT <= 3;  //205 / 63 = 3
    16'b11001101_01000000 : OUT <= 3;  //205 / 64 = 3
    16'b11001101_01000001 : OUT <= 3;  //205 / 65 = 3
    16'b11001101_01000010 : OUT <= 3;  //205 / 66 = 3
    16'b11001101_01000011 : OUT <= 3;  //205 / 67 = 3
    16'b11001101_01000100 : OUT <= 3;  //205 / 68 = 3
    16'b11001101_01000101 : OUT <= 2;  //205 / 69 = 2
    16'b11001101_01000110 : OUT <= 2;  //205 / 70 = 2
    16'b11001101_01000111 : OUT <= 2;  //205 / 71 = 2
    16'b11001101_01001000 : OUT <= 2;  //205 / 72 = 2
    16'b11001101_01001001 : OUT <= 2;  //205 / 73 = 2
    16'b11001101_01001010 : OUT <= 2;  //205 / 74 = 2
    16'b11001101_01001011 : OUT <= 2;  //205 / 75 = 2
    16'b11001101_01001100 : OUT <= 2;  //205 / 76 = 2
    16'b11001101_01001101 : OUT <= 2;  //205 / 77 = 2
    16'b11001101_01001110 : OUT <= 2;  //205 / 78 = 2
    16'b11001101_01001111 : OUT <= 2;  //205 / 79 = 2
    16'b11001101_01010000 : OUT <= 2;  //205 / 80 = 2
    16'b11001101_01010001 : OUT <= 2;  //205 / 81 = 2
    16'b11001101_01010010 : OUT <= 2;  //205 / 82 = 2
    16'b11001101_01010011 : OUT <= 2;  //205 / 83 = 2
    16'b11001101_01010100 : OUT <= 2;  //205 / 84 = 2
    16'b11001101_01010101 : OUT <= 2;  //205 / 85 = 2
    16'b11001101_01010110 : OUT <= 2;  //205 / 86 = 2
    16'b11001101_01010111 : OUT <= 2;  //205 / 87 = 2
    16'b11001101_01011000 : OUT <= 2;  //205 / 88 = 2
    16'b11001101_01011001 : OUT <= 2;  //205 / 89 = 2
    16'b11001101_01011010 : OUT <= 2;  //205 / 90 = 2
    16'b11001101_01011011 : OUT <= 2;  //205 / 91 = 2
    16'b11001101_01011100 : OUT <= 2;  //205 / 92 = 2
    16'b11001101_01011101 : OUT <= 2;  //205 / 93 = 2
    16'b11001101_01011110 : OUT <= 2;  //205 / 94 = 2
    16'b11001101_01011111 : OUT <= 2;  //205 / 95 = 2
    16'b11001101_01100000 : OUT <= 2;  //205 / 96 = 2
    16'b11001101_01100001 : OUT <= 2;  //205 / 97 = 2
    16'b11001101_01100010 : OUT <= 2;  //205 / 98 = 2
    16'b11001101_01100011 : OUT <= 2;  //205 / 99 = 2
    16'b11001101_01100100 : OUT <= 2;  //205 / 100 = 2
    16'b11001101_01100101 : OUT <= 2;  //205 / 101 = 2
    16'b11001101_01100110 : OUT <= 2;  //205 / 102 = 2
    16'b11001101_01100111 : OUT <= 1;  //205 / 103 = 1
    16'b11001101_01101000 : OUT <= 1;  //205 / 104 = 1
    16'b11001101_01101001 : OUT <= 1;  //205 / 105 = 1
    16'b11001101_01101010 : OUT <= 1;  //205 / 106 = 1
    16'b11001101_01101011 : OUT <= 1;  //205 / 107 = 1
    16'b11001101_01101100 : OUT <= 1;  //205 / 108 = 1
    16'b11001101_01101101 : OUT <= 1;  //205 / 109 = 1
    16'b11001101_01101110 : OUT <= 1;  //205 / 110 = 1
    16'b11001101_01101111 : OUT <= 1;  //205 / 111 = 1
    16'b11001101_01110000 : OUT <= 1;  //205 / 112 = 1
    16'b11001101_01110001 : OUT <= 1;  //205 / 113 = 1
    16'b11001101_01110010 : OUT <= 1;  //205 / 114 = 1
    16'b11001101_01110011 : OUT <= 1;  //205 / 115 = 1
    16'b11001101_01110100 : OUT <= 1;  //205 / 116 = 1
    16'b11001101_01110101 : OUT <= 1;  //205 / 117 = 1
    16'b11001101_01110110 : OUT <= 1;  //205 / 118 = 1
    16'b11001101_01110111 : OUT <= 1;  //205 / 119 = 1
    16'b11001101_01111000 : OUT <= 1;  //205 / 120 = 1
    16'b11001101_01111001 : OUT <= 1;  //205 / 121 = 1
    16'b11001101_01111010 : OUT <= 1;  //205 / 122 = 1
    16'b11001101_01111011 : OUT <= 1;  //205 / 123 = 1
    16'b11001101_01111100 : OUT <= 1;  //205 / 124 = 1
    16'b11001101_01111101 : OUT <= 1;  //205 / 125 = 1
    16'b11001101_01111110 : OUT <= 1;  //205 / 126 = 1
    16'b11001101_01111111 : OUT <= 1;  //205 / 127 = 1
    16'b11001101_10000000 : OUT <= 1;  //205 / 128 = 1
    16'b11001101_10000001 : OUT <= 1;  //205 / 129 = 1
    16'b11001101_10000010 : OUT <= 1;  //205 / 130 = 1
    16'b11001101_10000011 : OUT <= 1;  //205 / 131 = 1
    16'b11001101_10000100 : OUT <= 1;  //205 / 132 = 1
    16'b11001101_10000101 : OUT <= 1;  //205 / 133 = 1
    16'b11001101_10000110 : OUT <= 1;  //205 / 134 = 1
    16'b11001101_10000111 : OUT <= 1;  //205 / 135 = 1
    16'b11001101_10001000 : OUT <= 1;  //205 / 136 = 1
    16'b11001101_10001001 : OUT <= 1;  //205 / 137 = 1
    16'b11001101_10001010 : OUT <= 1;  //205 / 138 = 1
    16'b11001101_10001011 : OUT <= 1;  //205 / 139 = 1
    16'b11001101_10001100 : OUT <= 1;  //205 / 140 = 1
    16'b11001101_10001101 : OUT <= 1;  //205 / 141 = 1
    16'b11001101_10001110 : OUT <= 1;  //205 / 142 = 1
    16'b11001101_10001111 : OUT <= 1;  //205 / 143 = 1
    16'b11001101_10010000 : OUT <= 1;  //205 / 144 = 1
    16'b11001101_10010001 : OUT <= 1;  //205 / 145 = 1
    16'b11001101_10010010 : OUT <= 1;  //205 / 146 = 1
    16'b11001101_10010011 : OUT <= 1;  //205 / 147 = 1
    16'b11001101_10010100 : OUT <= 1;  //205 / 148 = 1
    16'b11001101_10010101 : OUT <= 1;  //205 / 149 = 1
    16'b11001101_10010110 : OUT <= 1;  //205 / 150 = 1
    16'b11001101_10010111 : OUT <= 1;  //205 / 151 = 1
    16'b11001101_10011000 : OUT <= 1;  //205 / 152 = 1
    16'b11001101_10011001 : OUT <= 1;  //205 / 153 = 1
    16'b11001101_10011010 : OUT <= 1;  //205 / 154 = 1
    16'b11001101_10011011 : OUT <= 1;  //205 / 155 = 1
    16'b11001101_10011100 : OUT <= 1;  //205 / 156 = 1
    16'b11001101_10011101 : OUT <= 1;  //205 / 157 = 1
    16'b11001101_10011110 : OUT <= 1;  //205 / 158 = 1
    16'b11001101_10011111 : OUT <= 1;  //205 / 159 = 1
    16'b11001101_10100000 : OUT <= 1;  //205 / 160 = 1
    16'b11001101_10100001 : OUT <= 1;  //205 / 161 = 1
    16'b11001101_10100010 : OUT <= 1;  //205 / 162 = 1
    16'b11001101_10100011 : OUT <= 1;  //205 / 163 = 1
    16'b11001101_10100100 : OUT <= 1;  //205 / 164 = 1
    16'b11001101_10100101 : OUT <= 1;  //205 / 165 = 1
    16'b11001101_10100110 : OUT <= 1;  //205 / 166 = 1
    16'b11001101_10100111 : OUT <= 1;  //205 / 167 = 1
    16'b11001101_10101000 : OUT <= 1;  //205 / 168 = 1
    16'b11001101_10101001 : OUT <= 1;  //205 / 169 = 1
    16'b11001101_10101010 : OUT <= 1;  //205 / 170 = 1
    16'b11001101_10101011 : OUT <= 1;  //205 / 171 = 1
    16'b11001101_10101100 : OUT <= 1;  //205 / 172 = 1
    16'b11001101_10101101 : OUT <= 1;  //205 / 173 = 1
    16'b11001101_10101110 : OUT <= 1;  //205 / 174 = 1
    16'b11001101_10101111 : OUT <= 1;  //205 / 175 = 1
    16'b11001101_10110000 : OUT <= 1;  //205 / 176 = 1
    16'b11001101_10110001 : OUT <= 1;  //205 / 177 = 1
    16'b11001101_10110010 : OUT <= 1;  //205 / 178 = 1
    16'b11001101_10110011 : OUT <= 1;  //205 / 179 = 1
    16'b11001101_10110100 : OUT <= 1;  //205 / 180 = 1
    16'b11001101_10110101 : OUT <= 1;  //205 / 181 = 1
    16'b11001101_10110110 : OUT <= 1;  //205 / 182 = 1
    16'b11001101_10110111 : OUT <= 1;  //205 / 183 = 1
    16'b11001101_10111000 : OUT <= 1;  //205 / 184 = 1
    16'b11001101_10111001 : OUT <= 1;  //205 / 185 = 1
    16'b11001101_10111010 : OUT <= 1;  //205 / 186 = 1
    16'b11001101_10111011 : OUT <= 1;  //205 / 187 = 1
    16'b11001101_10111100 : OUT <= 1;  //205 / 188 = 1
    16'b11001101_10111101 : OUT <= 1;  //205 / 189 = 1
    16'b11001101_10111110 : OUT <= 1;  //205 / 190 = 1
    16'b11001101_10111111 : OUT <= 1;  //205 / 191 = 1
    16'b11001101_11000000 : OUT <= 1;  //205 / 192 = 1
    16'b11001101_11000001 : OUT <= 1;  //205 / 193 = 1
    16'b11001101_11000010 : OUT <= 1;  //205 / 194 = 1
    16'b11001101_11000011 : OUT <= 1;  //205 / 195 = 1
    16'b11001101_11000100 : OUT <= 1;  //205 / 196 = 1
    16'b11001101_11000101 : OUT <= 1;  //205 / 197 = 1
    16'b11001101_11000110 : OUT <= 1;  //205 / 198 = 1
    16'b11001101_11000111 : OUT <= 1;  //205 / 199 = 1
    16'b11001101_11001000 : OUT <= 1;  //205 / 200 = 1
    16'b11001101_11001001 : OUT <= 1;  //205 / 201 = 1
    16'b11001101_11001010 : OUT <= 1;  //205 / 202 = 1
    16'b11001101_11001011 : OUT <= 1;  //205 / 203 = 1
    16'b11001101_11001100 : OUT <= 1;  //205 / 204 = 1
    16'b11001101_11001101 : OUT <= 1;  //205 / 205 = 1
    16'b11001101_11001110 : OUT <= 0;  //205 / 206 = 0
    16'b11001101_11001111 : OUT <= 0;  //205 / 207 = 0
    16'b11001101_11010000 : OUT <= 0;  //205 / 208 = 0
    16'b11001101_11010001 : OUT <= 0;  //205 / 209 = 0
    16'b11001101_11010010 : OUT <= 0;  //205 / 210 = 0
    16'b11001101_11010011 : OUT <= 0;  //205 / 211 = 0
    16'b11001101_11010100 : OUT <= 0;  //205 / 212 = 0
    16'b11001101_11010101 : OUT <= 0;  //205 / 213 = 0
    16'b11001101_11010110 : OUT <= 0;  //205 / 214 = 0
    16'b11001101_11010111 : OUT <= 0;  //205 / 215 = 0
    16'b11001101_11011000 : OUT <= 0;  //205 / 216 = 0
    16'b11001101_11011001 : OUT <= 0;  //205 / 217 = 0
    16'b11001101_11011010 : OUT <= 0;  //205 / 218 = 0
    16'b11001101_11011011 : OUT <= 0;  //205 / 219 = 0
    16'b11001101_11011100 : OUT <= 0;  //205 / 220 = 0
    16'b11001101_11011101 : OUT <= 0;  //205 / 221 = 0
    16'b11001101_11011110 : OUT <= 0;  //205 / 222 = 0
    16'b11001101_11011111 : OUT <= 0;  //205 / 223 = 0
    16'b11001101_11100000 : OUT <= 0;  //205 / 224 = 0
    16'b11001101_11100001 : OUT <= 0;  //205 / 225 = 0
    16'b11001101_11100010 : OUT <= 0;  //205 / 226 = 0
    16'b11001101_11100011 : OUT <= 0;  //205 / 227 = 0
    16'b11001101_11100100 : OUT <= 0;  //205 / 228 = 0
    16'b11001101_11100101 : OUT <= 0;  //205 / 229 = 0
    16'b11001101_11100110 : OUT <= 0;  //205 / 230 = 0
    16'b11001101_11100111 : OUT <= 0;  //205 / 231 = 0
    16'b11001101_11101000 : OUT <= 0;  //205 / 232 = 0
    16'b11001101_11101001 : OUT <= 0;  //205 / 233 = 0
    16'b11001101_11101010 : OUT <= 0;  //205 / 234 = 0
    16'b11001101_11101011 : OUT <= 0;  //205 / 235 = 0
    16'b11001101_11101100 : OUT <= 0;  //205 / 236 = 0
    16'b11001101_11101101 : OUT <= 0;  //205 / 237 = 0
    16'b11001101_11101110 : OUT <= 0;  //205 / 238 = 0
    16'b11001101_11101111 : OUT <= 0;  //205 / 239 = 0
    16'b11001101_11110000 : OUT <= 0;  //205 / 240 = 0
    16'b11001101_11110001 : OUT <= 0;  //205 / 241 = 0
    16'b11001101_11110010 : OUT <= 0;  //205 / 242 = 0
    16'b11001101_11110011 : OUT <= 0;  //205 / 243 = 0
    16'b11001101_11110100 : OUT <= 0;  //205 / 244 = 0
    16'b11001101_11110101 : OUT <= 0;  //205 / 245 = 0
    16'b11001101_11110110 : OUT <= 0;  //205 / 246 = 0
    16'b11001101_11110111 : OUT <= 0;  //205 / 247 = 0
    16'b11001101_11111000 : OUT <= 0;  //205 / 248 = 0
    16'b11001101_11111001 : OUT <= 0;  //205 / 249 = 0
    16'b11001101_11111010 : OUT <= 0;  //205 / 250 = 0
    16'b11001101_11111011 : OUT <= 0;  //205 / 251 = 0
    16'b11001101_11111100 : OUT <= 0;  //205 / 252 = 0
    16'b11001101_11111101 : OUT <= 0;  //205 / 253 = 0
    16'b11001101_11111110 : OUT <= 0;  //205 / 254 = 0
    16'b11001101_11111111 : OUT <= 0;  //205 / 255 = 0
    16'b11001110_00000000 : OUT <= 0;  //206 / 0 = 0
    16'b11001110_00000001 : OUT <= 206;  //206 / 1 = 206
    16'b11001110_00000010 : OUT <= 103;  //206 / 2 = 103
    16'b11001110_00000011 : OUT <= 68;  //206 / 3 = 68
    16'b11001110_00000100 : OUT <= 51;  //206 / 4 = 51
    16'b11001110_00000101 : OUT <= 41;  //206 / 5 = 41
    16'b11001110_00000110 : OUT <= 34;  //206 / 6 = 34
    16'b11001110_00000111 : OUT <= 29;  //206 / 7 = 29
    16'b11001110_00001000 : OUT <= 25;  //206 / 8 = 25
    16'b11001110_00001001 : OUT <= 22;  //206 / 9 = 22
    16'b11001110_00001010 : OUT <= 20;  //206 / 10 = 20
    16'b11001110_00001011 : OUT <= 18;  //206 / 11 = 18
    16'b11001110_00001100 : OUT <= 17;  //206 / 12 = 17
    16'b11001110_00001101 : OUT <= 15;  //206 / 13 = 15
    16'b11001110_00001110 : OUT <= 14;  //206 / 14 = 14
    16'b11001110_00001111 : OUT <= 13;  //206 / 15 = 13
    16'b11001110_00010000 : OUT <= 12;  //206 / 16 = 12
    16'b11001110_00010001 : OUT <= 12;  //206 / 17 = 12
    16'b11001110_00010010 : OUT <= 11;  //206 / 18 = 11
    16'b11001110_00010011 : OUT <= 10;  //206 / 19 = 10
    16'b11001110_00010100 : OUT <= 10;  //206 / 20 = 10
    16'b11001110_00010101 : OUT <= 9;  //206 / 21 = 9
    16'b11001110_00010110 : OUT <= 9;  //206 / 22 = 9
    16'b11001110_00010111 : OUT <= 8;  //206 / 23 = 8
    16'b11001110_00011000 : OUT <= 8;  //206 / 24 = 8
    16'b11001110_00011001 : OUT <= 8;  //206 / 25 = 8
    16'b11001110_00011010 : OUT <= 7;  //206 / 26 = 7
    16'b11001110_00011011 : OUT <= 7;  //206 / 27 = 7
    16'b11001110_00011100 : OUT <= 7;  //206 / 28 = 7
    16'b11001110_00011101 : OUT <= 7;  //206 / 29 = 7
    16'b11001110_00011110 : OUT <= 6;  //206 / 30 = 6
    16'b11001110_00011111 : OUT <= 6;  //206 / 31 = 6
    16'b11001110_00100000 : OUT <= 6;  //206 / 32 = 6
    16'b11001110_00100001 : OUT <= 6;  //206 / 33 = 6
    16'b11001110_00100010 : OUT <= 6;  //206 / 34 = 6
    16'b11001110_00100011 : OUT <= 5;  //206 / 35 = 5
    16'b11001110_00100100 : OUT <= 5;  //206 / 36 = 5
    16'b11001110_00100101 : OUT <= 5;  //206 / 37 = 5
    16'b11001110_00100110 : OUT <= 5;  //206 / 38 = 5
    16'b11001110_00100111 : OUT <= 5;  //206 / 39 = 5
    16'b11001110_00101000 : OUT <= 5;  //206 / 40 = 5
    16'b11001110_00101001 : OUT <= 5;  //206 / 41 = 5
    16'b11001110_00101010 : OUT <= 4;  //206 / 42 = 4
    16'b11001110_00101011 : OUT <= 4;  //206 / 43 = 4
    16'b11001110_00101100 : OUT <= 4;  //206 / 44 = 4
    16'b11001110_00101101 : OUT <= 4;  //206 / 45 = 4
    16'b11001110_00101110 : OUT <= 4;  //206 / 46 = 4
    16'b11001110_00101111 : OUT <= 4;  //206 / 47 = 4
    16'b11001110_00110000 : OUT <= 4;  //206 / 48 = 4
    16'b11001110_00110001 : OUT <= 4;  //206 / 49 = 4
    16'b11001110_00110010 : OUT <= 4;  //206 / 50 = 4
    16'b11001110_00110011 : OUT <= 4;  //206 / 51 = 4
    16'b11001110_00110100 : OUT <= 3;  //206 / 52 = 3
    16'b11001110_00110101 : OUT <= 3;  //206 / 53 = 3
    16'b11001110_00110110 : OUT <= 3;  //206 / 54 = 3
    16'b11001110_00110111 : OUT <= 3;  //206 / 55 = 3
    16'b11001110_00111000 : OUT <= 3;  //206 / 56 = 3
    16'b11001110_00111001 : OUT <= 3;  //206 / 57 = 3
    16'b11001110_00111010 : OUT <= 3;  //206 / 58 = 3
    16'b11001110_00111011 : OUT <= 3;  //206 / 59 = 3
    16'b11001110_00111100 : OUT <= 3;  //206 / 60 = 3
    16'b11001110_00111101 : OUT <= 3;  //206 / 61 = 3
    16'b11001110_00111110 : OUT <= 3;  //206 / 62 = 3
    16'b11001110_00111111 : OUT <= 3;  //206 / 63 = 3
    16'b11001110_01000000 : OUT <= 3;  //206 / 64 = 3
    16'b11001110_01000001 : OUT <= 3;  //206 / 65 = 3
    16'b11001110_01000010 : OUT <= 3;  //206 / 66 = 3
    16'b11001110_01000011 : OUT <= 3;  //206 / 67 = 3
    16'b11001110_01000100 : OUT <= 3;  //206 / 68 = 3
    16'b11001110_01000101 : OUT <= 2;  //206 / 69 = 2
    16'b11001110_01000110 : OUT <= 2;  //206 / 70 = 2
    16'b11001110_01000111 : OUT <= 2;  //206 / 71 = 2
    16'b11001110_01001000 : OUT <= 2;  //206 / 72 = 2
    16'b11001110_01001001 : OUT <= 2;  //206 / 73 = 2
    16'b11001110_01001010 : OUT <= 2;  //206 / 74 = 2
    16'b11001110_01001011 : OUT <= 2;  //206 / 75 = 2
    16'b11001110_01001100 : OUT <= 2;  //206 / 76 = 2
    16'b11001110_01001101 : OUT <= 2;  //206 / 77 = 2
    16'b11001110_01001110 : OUT <= 2;  //206 / 78 = 2
    16'b11001110_01001111 : OUT <= 2;  //206 / 79 = 2
    16'b11001110_01010000 : OUT <= 2;  //206 / 80 = 2
    16'b11001110_01010001 : OUT <= 2;  //206 / 81 = 2
    16'b11001110_01010010 : OUT <= 2;  //206 / 82 = 2
    16'b11001110_01010011 : OUT <= 2;  //206 / 83 = 2
    16'b11001110_01010100 : OUT <= 2;  //206 / 84 = 2
    16'b11001110_01010101 : OUT <= 2;  //206 / 85 = 2
    16'b11001110_01010110 : OUT <= 2;  //206 / 86 = 2
    16'b11001110_01010111 : OUT <= 2;  //206 / 87 = 2
    16'b11001110_01011000 : OUT <= 2;  //206 / 88 = 2
    16'b11001110_01011001 : OUT <= 2;  //206 / 89 = 2
    16'b11001110_01011010 : OUT <= 2;  //206 / 90 = 2
    16'b11001110_01011011 : OUT <= 2;  //206 / 91 = 2
    16'b11001110_01011100 : OUT <= 2;  //206 / 92 = 2
    16'b11001110_01011101 : OUT <= 2;  //206 / 93 = 2
    16'b11001110_01011110 : OUT <= 2;  //206 / 94 = 2
    16'b11001110_01011111 : OUT <= 2;  //206 / 95 = 2
    16'b11001110_01100000 : OUT <= 2;  //206 / 96 = 2
    16'b11001110_01100001 : OUT <= 2;  //206 / 97 = 2
    16'b11001110_01100010 : OUT <= 2;  //206 / 98 = 2
    16'b11001110_01100011 : OUT <= 2;  //206 / 99 = 2
    16'b11001110_01100100 : OUT <= 2;  //206 / 100 = 2
    16'b11001110_01100101 : OUT <= 2;  //206 / 101 = 2
    16'b11001110_01100110 : OUT <= 2;  //206 / 102 = 2
    16'b11001110_01100111 : OUT <= 2;  //206 / 103 = 2
    16'b11001110_01101000 : OUT <= 1;  //206 / 104 = 1
    16'b11001110_01101001 : OUT <= 1;  //206 / 105 = 1
    16'b11001110_01101010 : OUT <= 1;  //206 / 106 = 1
    16'b11001110_01101011 : OUT <= 1;  //206 / 107 = 1
    16'b11001110_01101100 : OUT <= 1;  //206 / 108 = 1
    16'b11001110_01101101 : OUT <= 1;  //206 / 109 = 1
    16'b11001110_01101110 : OUT <= 1;  //206 / 110 = 1
    16'b11001110_01101111 : OUT <= 1;  //206 / 111 = 1
    16'b11001110_01110000 : OUT <= 1;  //206 / 112 = 1
    16'b11001110_01110001 : OUT <= 1;  //206 / 113 = 1
    16'b11001110_01110010 : OUT <= 1;  //206 / 114 = 1
    16'b11001110_01110011 : OUT <= 1;  //206 / 115 = 1
    16'b11001110_01110100 : OUT <= 1;  //206 / 116 = 1
    16'b11001110_01110101 : OUT <= 1;  //206 / 117 = 1
    16'b11001110_01110110 : OUT <= 1;  //206 / 118 = 1
    16'b11001110_01110111 : OUT <= 1;  //206 / 119 = 1
    16'b11001110_01111000 : OUT <= 1;  //206 / 120 = 1
    16'b11001110_01111001 : OUT <= 1;  //206 / 121 = 1
    16'b11001110_01111010 : OUT <= 1;  //206 / 122 = 1
    16'b11001110_01111011 : OUT <= 1;  //206 / 123 = 1
    16'b11001110_01111100 : OUT <= 1;  //206 / 124 = 1
    16'b11001110_01111101 : OUT <= 1;  //206 / 125 = 1
    16'b11001110_01111110 : OUT <= 1;  //206 / 126 = 1
    16'b11001110_01111111 : OUT <= 1;  //206 / 127 = 1
    16'b11001110_10000000 : OUT <= 1;  //206 / 128 = 1
    16'b11001110_10000001 : OUT <= 1;  //206 / 129 = 1
    16'b11001110_10000010 : OUT <= 1;  //206 / 130 = 1
    16'b11001110_10000011 : OUT <= 1;  //206 / 131 = 1
    16'b11001110_10000100 : OUT <= 1;  //206 / 132 = 1
    16'b11001110_10000101 : OUT <= 1;  //206 / 133 = 1
    16'b11001110_10000110 : OUT <= 1;  //206 / 134 = 1
    16'b11001110_10000111 : OUT <= 1;  //206 / 135 = 1
    16'b11001110_10001000 : OUT <= 1;  //206 / 136 = 1
    16'b11001110_10001001 : OUT <= 1;  //206 / 137 = 1
    16'b11001110_10001010 : OUT <= 1;  //206 / 138 = 1
    16'b11001110_10001011 : OUT <= 1;  //206 / 139 = 1
    16'b11001110_10001100 : OUT <= 1;  //206 / 140 = 1
    16'b11001110_10001101 : OUT <= 1;  //206 / 141 = 1
    16'b11001110_10001110 : OUT <= 1;  //206 / 142 = 1
    16'b11001110_10001111 : OUT <= 1;  //206 / 143 = 1
    16'b11001110_10010000 : OUT <= 1;  //206 / 144 = 1
    16'b11001110_10010001 : OUT <= 1;  //206 / 145 = 1
    16'b11001110_10010010 : OUT <= 1;  //206 / 146 = 1
    16'b11001110_10010011 : OUT <= 1;  //206 / 147 = 1
    16'b11001110_10010100 : OUT <= 1;  //206 / 148 = 1
    16'b11001110_10010101 : OUT <= 1;  //206 / 149 = 1
    16'b11001110_10010110 : OUT <= 1;  //206 / 150 = 1
    16'b11001110_10010111 : OUT <= 1;  //206 / 151 = 1
    16'b11001110_10011000 : OUT <= 1;  //206 / 152 = 1
    16'b11001110_10011001 : OUT <= 1;  //206 / 153 = 1
    16'b11001110_10011010 : OUT <= 1;  //206 / 154 = 1
    16'b11001110_10011011 : OUT <= 1;  //206 / 155 = 1
    16'b11001110_10011100 : OUT <= 1;  //206 / 156 = 1
    16'b11001110_10011101 : OUT <= 1;  //206 / 157 = 1
    16'b11001110_10011110 : OUT <= 1;  //206 / 158 = 1
    16'b11001110_10011111 : OUT <= 1;  //206 / 159 = 1
    16'b11001110_10100000 : OUT <= 1;  //206 / 160 = 1
    16'b11001110_10100001 : OUT <= 1;  //206 / 161 = 1
    16'b11001110_10100010 : OUT <= 1;  //206 / 162 = 1
    16'b11001110_10100011 : OUT <= 1;  //206 / 163 = 1
    16'b11001110_10100100 : OUT <= 1;  //206 / 164 = 1
    16'b11001110_10100101 : OUT <= 1;  //206 / 165 = 1
    16'b11001110_10100110 : OUT <= 1;  //206 / 166 = 1
    16'b11001110_10100111 : OUT <= 1;  //206 / 167 = 1
    16'b11001110_10101000 : OUT <= 1;  //206 / 168 = 1
    16'b11001110_10101001 : OUT <= 1;  //206 / 169 = 1
    16'b11001110_10101010 : OUT <= 1;  //206 / 170 = 1
    16'b11001110_10101011 : OUT <= 1;  //206 / 171 = 1
    16'b11001110_10101100 : OUT <= 1;  //206 / 172 = 1
    16'b11001110_10101101 : OUT <= 1;  //206 / 173 = 1
    16'b11001110_10101110 : OUT <= 1;  //206 / 174 = 1
    16'b11001110_10101111 : OUT <= 1;  //206 / 175 = 1
    16'b11001110_10110000 : OUT <= 1;  //206 / 176 = 1
    16'b11001110_10110001 : OUT <= 1;  //206 / 177 = 1
    16'b11001110_10110010 : OUT <= 1;  //206 / 178 = 1
    16'b11001110_10110011 : OUT <= 1;  //206 / 179 = 1
    16'b11001110_10110100 : OUT <= 1;  //206 / 180 = 1
    16'b11001110_10110101 : OUT <= 1;  //206 / 181 = 1
    16'b11001110_10110110 : OUT <= 1;  //206 / 182 = 1
    16'b11001110_10110111 : OUT <= 1;  //206 / 183 = 1
    16'b11001110_10111000 : OUT <= 1;  //206 / 184 = 1
    16'b11001110_10111001 : OUT <= 1;  //206 / 185 = 1
    16'b11001110_10111010 : OUT <= 1;  //206 / 186 = 1
    16'b11001110_10111011 : OUT <= 1;  //206 / 187 = 1
    16'b11001110_10111100 : OUT <= 1;  //206 / 188 = 1
    16'b11001110_10111101 : OUT <= 1;  //206 / 189 = 1
    16'b11001110_10111110 : OUT <= 1;  //206 / 190 = 1
    16'b11001110_10111111 : OUT <= 1;  //206 / 191 = 1
    16'b11001110_11000000 : OUT <= 1;  //206 / 192 = 1
    16'b11001110_11000001 : OUT <= 1;  //206 / 193 = 1
    16'b11001110_11000010 : OUT <= 1;  //206 / 194 = 1
    16'b11001110_11000011 : OUT <= 1;  //206 / 195 = 1
    16'b11001110_11000100 : OUT <= 1;  //206 / 196 = 1
    16'b11001110_11000101 : OUT <= 1;  //206 / 197 = 1
    16'b11001110_11000110 : OUT <= 1;  //206 / 198 = 1
    16'b11001110_11000111 : OUT <= 1;  //206 / 199 = 1
    16'b11001110_11001000 : OUT <= 1;  //206 / 200 = 1
    16'b11001110_11001001 : OUT <= 1;  //206 / 201 = 1
    16'b11001110_11001010 : OUT <= 1;  //206 / 202 = 1
    16'b11001110_11001011 : OUT <= 1;  //206 / 203 = 1
    16'b11001110_11001100 : OUT <= 1;  //206 / 204 = 1
    16'b11001110_11001101 : OUT <= 1;  //206 / 205 = 1
    16'b11001110_11001110 : OUT <= 1;  //206 / 206 = 1
    16'b11001110_11001111 : OUT <= 0;  //206 / 207 = 0
    16'b11001110_11010000 : OUT <= 0;  //206 / 208 = 0
    16'b11001110_11010001 : OUT <= 0;  //206 / 209 = 0
    16'b11001110_11010010 : OUT <= 0;  //206 / 210 = 0
    16'b11001110_11010011 : OUT <= 0;  //206 / 211 = 0
    16'b11001110_11010100 : OUT <= 0;  //206 / 212 = 0
    16'b11001110_11010101 : OUT <= 0;  //206 / 213 = 0
    16'b11001110_11010110 : OUT <= 0;  //206 / 214 = 0
    16'b11001110_11010111 : OUT <= 0;  //206 / 215 = 0
    16'b11001110_11011000 : OUT <= 0;  //206 / 216 = 0
    16'b11001110_11011001 : OUT <= 0;  //206 / 217 = 0
    16'b11001110_11011010 : OUT <= 0;  //206 / 218 = 0
    16'b11001110_11011011 : OUT <= 0;  //206 / 219 = 0
    16'b11001110_11011100 : OUT <= 0;  //206 / 220 = 0
    16'b11001110_11011101 : OUT <= 0;  //206 / 221 = 0
    16'b11001110_11011110 : OUT <= 0;  //206 / 222 = 0
    16'b11001110_11011111 : OUT <= 0;  //206 / 223 = 0
    16'b11001110_11100000 : OUT <= 0;  //206 / 224 = 0
    16'b11001110_11100001 : OUT <= 0;  //206 / 225 = 0
    16'b11001110_11100010 : OUT <= 0;  //206 / 226 = 0
    16'b11001110_11100011 : OUT <= 0;  //206 / 227 = 0
    16'b11001110_11100100 : OUT <= 0;  //206 / 228 = 0
    16'b11001110_11100101 : OUT <= 0;  //206 / 229 = 0
    16'b11001110_11100110 : OUT <= 0;  //206 / 230 = 0
    16'b11001110_11100111 : OUT <= 0;  //206 / 231 = 0
    16'b11001110_11101000 : OUT <= 0;  //206 / 232 = 0
    16'b11001110_11101001 : OUT <= 0;  //206 / 233 = 0
    16'b11001110_11101010 : OUT <= 0;  //206 / 234 = 0
    16'b11001110_11101011 : OUT <= 0;  //206 / 235 = 0
    16'b11001110_11101100 : OUT <= 0;  //206 / 236 = 0
    16'b11001110_11101101 : OUT <= 0;  //206 / 237 = 0
    16'b11001110_11101110 : OUT <= 0;  //206 / 238 = 0
    16'b11001110_11101111 : OUT <= 0;  //206 / 239 = 0
    16'b11001110_11110000 : OUT <= 0;  //206 / 240 = 0
    16'b11001110_11110001 : OUT <= 0;  //206 / 241 = 0
    16'b11001110_11110010 : OUT <= 0;  //206 / 242 = 0
    16'b11001110_11110011 : OUT <= 0;  //206 / 243 = 0
    16'b11001110_11110100 : OUT <= 0;  //206 / 244 = 0
    16'b11001110_11110101 : OUT <= 0;  //206 / 245 = 0
    16'b11001110_11110110 : OUT <= 0;  //206 / 246 = 0
    16'b11001110_11110111 : OUT <= 0;  //206 / 247 = 0
    16'b11001110_11111000 : OUT <= 0;  //206 / 248 = 0
    16'b11001110_11111001 : OUT <= 0;  //206 / 249 = 0
    16'b11001110_11111010 : OUT <= 0;  //206 / 250 = 0
    16'b11001110_11111011 : OUT <= 0;  //206 / 251 = 0
    16'b11001110_11111100 : OUT <= 0;  //206 / 252 = 0
    16'b11001110_11111101 : OUT <= 0;  //206 / 253 = 0
    16'b11001110_11111110 : OUT <= 0;  //206 / 254 = 0
    16'b11001110_11111111 : OUT <= 0;  //206 / 255 = 0
    16'b11001111_00000000 : OUT <= 0;  //207 / 0 = 0
    16'b11001111_00000001 : OUT <= 207;  //207 / 1 = 207
    16'b11001111_00000010 : OUT <= 103;  //207 / 2 = 103
    16'b11001111_00000011 : OUT <= 69;  //207 / 3 = 69
    16'b11001111_00000100 : OUT <= 51;  //207 / 4 = 51
    16'b11001111_00000101 : OUT <= 41;  //207 / 5 = 41
    16'b11001111_00000110 : OUT <= 34;  //207 / 6 = 34
    16'b11001111_00000111 : OUT <= 29;  //207 / 7 = 29
    16'b11001111_00001000 : OUT <= 25;  //207 / 8 = 25
    16'b11001111_00001001 : OUT <= 23;  //207 / 9 = 23
    16'b11001111_00001010 : OUT <= 20;  //207 / 10 = 20
    16'b11001111_00001011 : OUT <= 18;  //207 / 11 = 18
    16'b11001111_00001100 : OUT <= 17;  //207 / 12 = 17
    16'b11001111_00001101 : OUT <= 15;  //207 / 13 = 15
    16'b11001111_00001110 : OUT <= 14;  //207 / 14 = 14
    16'b11001111_00001111 : OUT <= 13;  //207 / 15 = 13
    16'b11001111_00010000 : OUT <= 12;  //207 / 16 = 12
    16'b11001111_00010001 : OUT <= 12;  //207 / 17 = 12
    16'b11001111_00010010 : OUT <= 11;  //207 / 18 = 11
    16'b11001111_00010011 : OUT <= 10;  //207 / 19 = 10
    16'b11001111_00010100 : OUT <= 10;  //207 / 20 = 10
    16'b11001111_00010101 : OUT <= 9;  //207 / 21 = 9
    16'b11001111_00010110 : OUT <= 9;  //207 / 22 = 9
    16'b11001111_00010111 : OUT <= 9;  //207 / 23 = 9
    16'b11001111_00011000 : OUT <= 8;  //207 / 24 = 8
    16'b11001111_00011001 : OUT <= 8;  //207 / 25 = 8
    16'b11001111_00011010 : OUT <= 7;  //207 / 26 = 7
    16'b11001111_00011011 : OUT <= 7;  //207 / 27 = 7
    16'b11001111_00011100 : OUT <= 7;  //207 / 28 = 7
    16'b11001111_00011101 : OUT <= 7;  //207 / 29 = 7
    16'b11001111_00011110 : OUT <= 6;  //207 / 30 = 6
    16'b11001111_00011111 : OUT <= 6;  //207 / 31 = 6
    16'b11001111_00100000 : OUT <= 6;  //207 / 32 = 6
    16'b11001111_00100001 : OUT <= 6;  //207 / 33 = 6
    16'b11001111_00100010 : OUT <= 6;  //207 / 34 = 6
    16'b11001111_00100011 : OUT <= 5;  //207 / 35 = 5
    16'b11001111_00100100 : OUT <= 5;  //207 / 36 = 5
    16'b11001111_00100101 : OUT <= 5;  //207 / 37 = 5
    16'b11001111_00100110 : OUT <= 5;  //207 / 38 = 5
    16'b11001111_00100111 : OUT <= 5;  //207 / 39 = 5
    16'b11001111_00101000 : OUT <= 5;  //207 / 40 = 5
    16'b11001111_00101001 : OUT <= 5;  //207 / 41 = 5
    16'b11001111_00101010 : OUT <= 4;  //207 / 42 = 4
    16'b11001111_00101011 : OUT <= 4;  //207 / 43 = 4
    16'b11001111_00101100 : OUT <= 4;  //207 / 44 = 4
    16'b11001111_00101101 : OUT <= 4;  //207 / 45 = 4
    16'b11001111_00101110 : OUT <= 4;  //207 / 46 = 4
    16'b11001111_00101111 : OUT <= 4;  //207 / 47 = 4
    16'b11001111_00110000 : OUT <= 4;  //207 / 48 = 4
    16'b11001111_00110001 : OUT <= 4;  //207 / 49 = 4
    16'b11001111_00110010 : OUT <= 4;  //207 / 50 = 4
    16'b11001111_00110011 : OUT <= 4;  //207 / 51 = 4
    16'b11001111_00110100 : OUT <= 3;  //207 / 52 = 3
    16'b11001111_00110101 : OUT <= 3;  //207 / 53 = 3
    16'b11001111_00110110 : OUT <= 3;  //207 / 54 = 3
    16'b11001111_00110111 : OUT <= 3;  //207 / 55 = 3
    16'b11001111_00111000 : OUT <= 3;  //207 / 56 = 3
    16'b11001111_00111001 : OUT <= 3;  //207 / 57 = 3
    16'b11001111_00111010 : OUT <= 3;  //207 / 58 = 3
    16'b11001111_00111011 : OUT <= 3;  //207 / 59 = 3
    16'b11001111_00111100 : OUT <= 3;  //207 / 60 = 3
    16'b11001111_00111101 : OUT <= 3;  //207 / 61 = 3
    16'b11001111_00111110 : OUT <= 3;  //207 / 62 = 3
    16'b11001111_00111111 : OUT <= 3;  //207 / 63 = 3
    16'b11001111_01000000 : OUT <= 3;  //207 / 64 = 3
    16'b11001111_01000001 : OUT <= 3;  //207 / 65 = 3
    16'b11001111_01000010 : OUT <= 3;  //207 / 66 = 3
    16'b11001111_01000011 : OUT <= 3;  //207 / 67 = 3
    16'b11001111_01000100 : OUT <= 3;  //207 / 68 = 3
    16'b11001111_01000101 : OUT <= 3;  //207 / 69 = 3
    16'b11001111_01000110 : OUT <= 2;  //207 / 70 = 2
    16'b11001111_01000111 : OUT <= 2;  //207 / 71 = 2
    16'b11001111_01001000 : OUT <= 2;  //207 / 72 = 2
    16'b11001111_01001001 : OUT <= 2;  //207 / 73 = 2
    16'b11001111_01001010 : OUT <= 2;  //207 / 74 = 2
    16'b11001111_01001011 : OUT <= 2;  //207 / 75 = 2
    16'b11001111_01001100 : OUT <= 2;  //207 / 76 = 2
    16'b11001111_01001101 : OUT <= 2;  //207 / 77 = 2
    16'b11001111_01001110 : OUT <= 2;  //207 / 78 = 2
    16'b11001111_01001111 : OUT <= 2;  //207 / 79 = 2
    16'b11001111_01010000 : OUT <= 2;  //207 / 80 = 2
    16'b11001111_01010001 : OUT <= 2;  //207 / 81 = 2
    16'b11001111_01010010 : OUT <= 2;  //207 / 82 = 2
    16'b11001111_01010011 : OUT <= 2;  //207 / 83 = 2
    16'b11001111_01010100 : OUT <= 2;  //207 / 84 = 2
    16'b11001111_01010101 : OUT <= 2;  //207 / 85 = 2
    16'b11001111_01010110 : OUT <= 2;  //207 / 86 = 2
    16'b11001111_01010111 : OUT <= 2;  //207 / 87 = 2
    16'b11001111_01011000 : OUT <= 2;  //207 / 88 = 2
    16'b11001111_01011001 : OUT <= 2;  //207 / 89 = 2
    16'b11001111_01011010 : OUT <= 2;  //207 / 90 = 2
    16'b11001111_01011011 : OUT <= 2;  //207 / 91 = 2
    16'b11001111_01011100 : OUT <= 2;  //207 / 92 = 2
    16'b11001111_01011101 : OUT <= 2;  //207 / 93 = 2
    16'b11001111_01011110 : OUT <= 2;  //207 / 94 = 2
    16'b11001111_01011111 : OUT <= 2;  //207 / 95 = 2
    16'b11001111_01100000 : OUT <= 2;  //207 / 96 = 2
    16'b11001111_01100001 : OUT <= 2;  //207 / 97 = 2
    16'b11001111_01100010 : OUT <= 2;  //207 / 98 = 2
    16'b11001111_01100011 : OUT <= 2;  //207 / 99 = 2
    16'b11001111_01100100 : OUT <= 2;  //207 / 100 = 2
    16'b11001111_01100101 : OUT <= 2;  //207 / 101 = 2
    16'b11001111_01100110 : OUT <= 2;  //207 / 102 = 2
    16'b11001111_01100111 : OUT <= 2;  //207 / 103 = 2
    16'b11001111_01101000 : OUT <= 1;  //207 / 104 = 1
    16'b11001111_01101001 : OUT <= 1;  //207 / 105 = 1
    16'b11001111_01101010 : OUT <= 1;  //207 / 106 = 1
    16'b11001111_01101011 : OUT <= 1;  //207 / 107 = 1
    16'b11001111_01101100 : OUT <= 1;  //207 / 108 = 1
    16'b11001111_01101101 : OUT <= 1;  //207 / 109 = 1
    16'b11001111_01101110 : OUT <= 1;  //207 / 110 = 1
    16'b11001111_01101111 : OUT <= 1;  //207 / 111 = 1
    16'b11001111_01110000 : OUT <= 1;  //207 / 112 = 1
    16'b11001111_01110001 : OUT <= 1;  //207 / 113 = 1
    16'b11001111_01110010 : OUT <= 1;  //207 / 114 = 1
    16'b11001111_01110011 : OUT <= 1;  //207 / 115 = 1
    16'b11001111_01110100 : OUT <= 1;  //207 / 116 = 1
    16'b11001111_01110101 : OUT <= 1;  //207 / 117 = 1
    16'b11001111_01110110 : OUT <= 1;  //207 / 118 = 1
    16'b11001111_01110111 : OUT <= 1;  //207 / 119 = 1
    16'b11001111_01111000 : OUT <= 1;  //207 / 120 = 1
    16'b11001111_01111001 : OUT <= 1;  //207 / 121 = 1
    16'b11001111_01111010 : OUT <= 1;  //207 / 122 = 1
    16'b11001111_01111011 : OUT <= 1;  //207 / 123 = 1
    16'b11001111_01111100 : OUT <= 1;  //207 / 124 = 1
    16'b11001111_01111101 : OUT <= 1;  //207 / 125 = 1
    16'b11001111_01111110 : OUT <= 1;  //207 / 126 = 1
    16'b11001111_01111111 : OUT <= 1;  //207 / 127 = 1
    16'b11001111_10000000 : OUT <= 1;  //207 / 128 = 1
    16'b11001111_10000001 : OUT <= 1;  //207 / 129 = 1
    16'b11001111_10000010 : OUT <= 1;  //207 / 130 = 1
    16'b11001111_10000011 : OUT <= 1;  //207 / 131 = 1
    16'b11001111_10000100 : OUT <= 1;  //207 / 132 = 1
    16'b11001111_10000101 : OUT <= 1;  //207 / 133 = 1
    16'b11001111_10000110 : OUT <= 1;  //207 / 134 = 1
    16'b11001111_10000111 : OUT <= 1;  //207 / 135 = 1
    16'b11001111_10001000 : OUT <= 1;  //207 / 136 = 1
    16'b11001111_10001001 : OUT <= 1;  //207 / 137 = 1
    16'b11001111_10001010 : OUT <= 1;  //207 / 138 = 1
    16'b11001111_10001011 : OUT <= 1;  //207 / 139 = 1
    16'b11001111_10001100 : OUT <= 1;  //207 / 140 = 1
    16'b11001111_10001101 : OUT <= 1;  //207 / 141 = 1
    16'b11001111_10001110 : OUT <= 1;  //207 / 142 = 1
    16'b11001111_10001111 : OUT <= 1;  //207 / 143 = 1
    16'b11001111_10010000 : OUT <= 1;  //207 / 144 = 1
    16'b11001111_10010001 : OUT <= 1;  //207 / 145 = 1
    16'b11001111_10010010 : OUT <= 1;  //207 / 146 = 1
    16'b11001111_10010011 : OUT <= 1;  //207 / 147 = 1
    16'b11001111_10010100 : OUT <= 1;  //207 / 148 = 1
    16'b11001111_10010101 : OUT <= 1;  //207 / 149 = 1
    16'b11001111_10010110 : OUT <= 1;  //207 / 150 = 1
    16'b11001111_10010111 : OUT <= 1;  //207 / 151 = 1
    16'b11001111_10011000 : OUT <= 1;  //207 / 152 = 1
    16'b11001111_10011001 : OUT <= 1;  //207 / 153 = 1
    16'b11001111_10011010 : OUT <= 1;  //207 / 154 = 1
    16'b11001111_10011011 : OUT <= 1;  //207 / 155 = 1
    16'b11001111_10011100 : OUT <= 1;  //207 / 156 = 1
    16'b11001111_10011101 : OUT <= 1;  //207 / 157 = 1
    16'b11001111_10011110 : OUT <= 1;  //207 / 158 = 1
    16'b11001111_10011111 : OUT <= 1;  //207 / 159 = 1
    16'b11001111_10100000 : OUT <= 1;  //207 / 160 = 1
    16'b11001111_10100001 : OUT <= 1;  //207 / 161 = 1
    16'b11001111_10100010 : OUT <= 1;  //207 / 162 = 1
    16'b11001111_10100011 : OUT <= 1;  //207 / 163 = 1
    16'b11001111_10100100 : OUT <= 1;  //207 / 164 = 1
    16'b11001111_10100101 : OUT <= 1;  //207 / 165 = 1
    16'b11001111_10100110 : OUT <= 1;  //207 / 166 = 1
    16'b11001111_10100111 : OUT <= 1;  //207 / 167 = 1
    16'b11001111_10101000 : OUT <= 1;  //207 / 168 = 1
    16'b11001111_10101001 : OUT <= 1;  //207 / 169 = 1
    16'b11001111_10101010 : OUT <= 1;  //207 / 170 = 1
    16'b11001111_10101011 : OUT <= 1;  //207 / 171 = 1
    16'b11001111_10101100 : OUT <= 1;  //207 / 172 = 1
    16'b11001111_10101101 : OUT <= 1;  //207 / 173 = 1
    16'b11001111_10101110 : OUT <= 1;  //207 / 174 = 1
    16'b11001111_10101111 : OUT <= 1;  //207 / 175 = 1
    16'b11001111_10110000 : OUT <= 1;  //207 / 176 = 1
    16'b11001111_10110001 : OUT <= 1;  //207 / 177 = 1
    16'b11001111_10110010 : OUT <= 1;  //207 / 178 = 1
    16'b11001111_10110011 : OUT <= 1;  //207 / 179 = 1
    16'b11001111_10110100 : OUT <= 1;  //207 / 180 = 1
    16'b11001111_10110101 : OUT <= 1;  //207 / 181 = 1
    16'b11001111_10110110 : OUT <= 1;  //207 / 182 = 1
    16'b11001111_10110111 : OUT <= 1;  //207 / 183 = 1
    16'b11001111_10111000 : OUT <= 1;  //207 / 184 = 1
    16'b11001111_10111001 : OUT <= 1;  //207 / 185 = 1
    16'b11001111_10111010 : OUT <= 1;  //207 / 186 = 1
    16'b11001111_10111011 : OUT <= 1;  //207 / 187 = 1
    16'b11001111_10111100 : OUT <= 1;  //207 / 188 = 1
    16'b11001111_10111101 : OUT <= 1;  //207 / 189 = 1
    16'b11001111_10111110 : OUT <= 1;  //207 / 190 = 1
    16'b11001111_10111111 : OUT <= 1;  //207 / 191 = 1
    16'b11001111_11000000 : OUT <= 1;  //207 / 192 = 1
    16'b11001111_11000001 : OUT <= 1;  //207 / 193 = 1
    16'b11001111_11000010 : OUT <= 1;  //207 / 194 = 1
    16'b11001111_11000011 : OUT <= 1;  //207 / 195 = 1
    16'b11001111_11000100 : OUT <= 1;  //207 / 196 = 1
    16'b11001111_11000101 : OUT <= 1;  //207 / 197 = 1
    16'b11001111_11000110 : OUT <= 1;  //207 / 198 = 1
    16'b11001111_11000111 : OUT <= 1;  //207 / 199 = 1
    16'b11001111_11001000 : OUT <= 1;  //207 / 200 = 1
    16'b11001111_11001001 : OUT <= 1;  //207 / 201 = 1
    16'b11001111_11001010 : OUT <= 1;  //207 / 202 = 1
    16'b11001111_11001011 : OUT <= 1;  //207 / 203 = 1
    16'b11001111_11001100 : OUT <= 1;  //207 / 204 = 1
    16'b11001111_11001101 : OUT <= 1;  //207 / 205 = 1
    16'b11001111_11001110 : OUT <= 1;  //207 / 206 = 1
    16'b11001111_11001111 : OUT <= 1;  //207 / 207 = 1
    16'b11001111_11010000 : OUT <= 0;  //207 / 208 = 0
    16'b11001111_11010001 : OUT <= 0;  //207 / 209 = 0
    16'b11001111_11010010 : OUT <= 0;  //207 / 210 = 0
    16'b11001111_11010011 : OUT <= 0;  //207 / 211 = 0
    16'b11001111_11010100 : OUT <= 0;  //207 / 212 = 0
    16'b11001111_11010101 : OUT <= 0;  //207 / 213 = 0
    16'b11001111_11010110 : OUT <= 0;  //207 / 214 = 0
    16'b11001111_11010111 : OUT <= 0;  //207 / 215 = 0
    16'b11001111_11011000 : OUT <= 0;  //207 / 216 = 0
    16'b11001111_11011001 : OUT <= 0;  //207 / 217 = 0
    16'b11001111_11011010 : OUT <= 0;  //207 / 218 = 0
    16'b11001111_11011011 : OUT <= 0;  //207 / 219 = 0
    16'b11001111_11011100 : OUT <= 0;  //207 / 220 = 0
    16'b11001111_11011101 : OUT <= 0;  //207 / 221 = 0
    16'b11001111_11011110 : OUT <= 0;  //207 / 222 = 0
    16'b11001111_11011111 : OUT <= 0;  //207 / 223 = 0
    16'b11001111_11100000 : OUT <= 0;  //207 / 224 = 0
    16'b11001111_11100001 : OUT <= 0;  //207 / 225 = 0
    16'b11001111_11100010 : OUT <= 0;  //207 / 226 = 0
    16'b11001111_11100011 : OUT <= 0;  //207 / 227 = 0
    16'b11001111_11100100 : OUT <= 0;  //207 / 228 = 0
    16'b11001111_11100101 : OUT <= 0;  //207 / 229 = 0
    16'b11001111_11100110 : OUT <= 0;  //207 / 230 = 0
    16'b11001111_11100111 : OUT <= 0;  //207 / 231 = 0
    16'b11001111_11101000 : OUT <= 0;  //207 / 232 = 0
    16'b11001111_11101001 : OUT <= 0;  //207 / 233 = 0
    16'b11001111_11101010 : OUT <= 0;  //207 / 234 = 0
    16'b11001111_11101011 : OUT <= 0;  //207 / 235 = 0
    16'b11001111_11101100 : OUT <= 0;  //207 / 236 = 0
    16'b11001111_11101101 : OUT <= 0;  //207 / 237 = 0
    16'b11001111_11101110 : OUT <= 0;  //207 / 238 = 0
    16'b11001111_11101111 : OUT <= 0;  //207 / 239 = 0
    16'b11001111_11110000 : OUT <= 0;  //207 / 240 = 0
    16'b11001111_11110001 : OUT <= 0;  //207 / 241 = 0
    16'b11001111_11110010 : OUT <= 0;  //207 / 242 = 0
    16'b11001111_11110011 : OUT <= 0;  //207 / 243 = 0
    16'b11001111_11110100 : OUT <= 0;  //207 / 244 = 0
    16'b11001111_11110101 : OUT <= 0;  //207 / 245 = 0
    16'b11001111_11110110 : OUT <= 0;  //207 / 246 = 0
    16'b11001111_11110111 : OUT <= 0;  //207 / 247 = 0
    16'b11001111_11111000 : OUT <= 0;  //207 / 248 = 0
    16'b11001111_11111001 : OUT <= 0;  //207 / 249 = 0
    16'b11001111_11111010 : OUT <= 0;  //207 / 250 = 0
    16'b11001111_11111011 : OUT <= 0;  //207 / 251 = 0
    16'b11001111_11111100 : OUT <= 0;  //207 / 252 = 0
    16'b11001111_11111101 : OUT <= 0;  //207 / 253 = 0
    16'b11001111_11111110 : OUT <= 0;  //207 / 254 = 0
    16'b11001111_11111111 : OUT <= 0;  //207 / 255 = 0
    16'b11010000_00000000 : OUT <= 0;  //208 / 0 = 0
    16'b11010000_00000001 : OUT <= 208;  //208 / 1 = 208
    16'b11010000_00000010 : OUT <= 104;  //208 / 2 = 104
    16'b11010000_00000011 : OUT <= 69;  //208 / 3 = 69
    16'b11010000_00000100 : OUT <= 52;  //208 / 4 = 52
    16'b11010000_00000101 : OUT <= 41;  //208 / 5 = 41
    16'b11010000_00000110 : OUT <= 34;  //208 / 6 = 34
    16'b11010000_00000111 : OUT <= 29;  //208 / 7 = 29
    16'b11010000_00001000 : OUT <= 26;  //208 / 8 = 26
    16'b11010000_00001001 : OUT <= 23;  //208 / 9 = 23
    16'b11010000_00001010 : OUT <= 20;  //208 / 10 = 20
    16'b11010000_00001011 : OUT <= 18;  //208 / 11 = 18
    16'b11010000_00001100 : OUT <= 17;  //208 / 12 = 17
    16'b11010000_00001101 : OUT <= 16;  //208 / 13 = 16
    16'b11010000_00001110 : OUT <= 14;  //208 / 14 = 14
    16'b11010000_00001111 : OUT <= 13;  //208 / 15 = 13
    16'b11010000_00010000 : OUT <= 13;  //208 / 16 = 13
    16'b11010000_00010001 : OUT <= 12;  //208 / 17 = 12
    16'b11010000_00010010 : OUT <= 11;  //208 / 18 = 11
    16'b11010000_00010011 : OUT <= 10;  //208 / 19 = 10
    16'b11010000_00010100 : OUT <= 10;  //208 / 20 = 10
    16'b11010000_00010101 : OUT <= 9;  //208 / 21 = 9
    16'b11010000_00010110 : OUT <= 9;  //208 / 22 = 9
    16'b11010000_00010111 : OUT <= 9;  //208 / 23 = 9
    16'b11010000_00011000 : OUT <= 8;  //208 / 24 = 8
    16'b11010000_00011001 : OUT <= 8;  //208 / 25 = 8
    16'b11010000_00011010 : OUT <= 8;  //208 / 26 = 8
    16'b11010000_00011011 : OUT <= 7;  //208 / 27 = 7
    16'b11010000_00011100 : OUT <= 7;  //208 / 28 = 7
    16'b11010000_00011101 : OUT <= 7;  //208 / 29 = 7
    16'b11010000_00011110 : OUT <= 6;  //208 / 30 = 6
    16'b11010000_00011111 : OUT <= 6;  //208 / 31 = 6
    16'b11010000_00100000 : OUT <= 6;  //208 / 32 = 6
    16'b11010000_00100001 : OUT <= 6;  //208 / 33 = 6
    16'b11010000_00100010 : OUT <= 6;  //208 / 34 = 6
    16'b11010000_00100011 : OUT <= 5;  //208 / 35 = 5
    16'b11010000_00100100 : OUT <= 5;  //208 / 36 = 5
    16'b11010000_00100101 : OUT <= 5;  //208 / 37 = 5
    16'b11010000_00100110 : OUT <= 5;  //208 / 38 = 5
    16'b11010000_00100111 : OUT <= 5;  //208 / 39 = 5
    16'b11010000_00101000 : OUT <= 5;  //208 / 40 = 5
    16'b11010000_00101001 : OUT <= 5;  //208 / 41 = 5
    16'b11010000_00101010 : OUT <= 4;  //208 / 42 = 4
    16'b11010000_00101011 : OUT <= 4;  //208 / 43 = 4
    16'b11010000_00101100 : OUT <= 4;  //208 / 44 = 4
    16'b11010000_00101101 : OUT <= 4;  //208 / 45 = 4
    16'b11010000_00101110 : OUT <= 4;  //208 / 46 = 4
    16'b11010000_00101111 : OUT <= 4;  //208 / 47 = 4
    16'b11010000_00110000 : OUT <= 4;  //208 / 48 = 4
    16'b11010000_00110001 : OUT <= 4;  //208 / 49 = 4
    16'b11010000_00110010 : OUT <= 4;  //208 / 50 = 4
    16'b11010000_00110011 : OUT <= 4;  //208 / 51 = 4
    16'b11010000_00110100 : OUT <= 4;  //208 / 52 = 4
    16'b11010000_00110101 : OUT <= 3;  //208 / 53 = 3
    16'b11010000_00110110 : OUT <= 3;  //208 / 54 = 3
    16'b11010000_00110111 : OUT <= 3;  //208 / 55 = 3
    16'b11010000_00111000 : OUT <= 3;  //208 / 56 = 3
    16'b11010000_00111001 : OUT <= 3;  //208 / 57 = 3
    16'b11010000_00111010 : OUT <= 3;  //208 / 58 = 3
    16'b11010000_00111011 : OUT <= 3;  //208 / 59 = 3
    16'b11010000_00111100 : OUT <= 3;  //208 / 60 = 3
    16'b11010000_00111101 : OUT <= 3;  //208 / 61 = 3
    16'b11010000_00111110 : OUT <= 3;  //208 / 62 = 3
    16'b11010000_00111111 : OUT <= 3;  //208 / 63 = 3
    16'b11010000_01000000 : OUT <= 3;  //208 / 64 = 3
    16'b11010000_01000001 : OUT <= 3;  //208 / 65 = 3
    16'b11010000_01000010 : OUT <= 3;  //208 / 66 = 3
    16'b11010000_01000011 : OUT <= 3;  //208 / 67 = 3
    16'b11010000_01000100 : OUT <= 3;  //208 / 68 = 3
    16'b11010000_01000101 : OUT <= 3;  //208 / 69 = 3
    16'b11010000_01000110 : OUT <= 2;  //208 / 70 = 2
    16'b11010000_01000111 : OUT <= 2;  //208 / 71 = 2
    16'b11010000_01001000 : OUT <= 2;  //208 / 72 = 2
    16'b11010000_01001001 : OUT <= 2;  //208 / 73 = 2
    16'b11010000_01001010 : OUT <= 2;  //208 / 74 = 2
    16'b11010000_01001011 : OUT <= 2;  //208 / 75 = 2
    16'b11010000_01001100 : OUT <= 2;  //208 / 76 = 2
    16'b11010000_01001101 : OUT <= 2;  //208 / 77 = 2
    16'b11010000_01001110 : OUT <= 2;  //208 / 78 = 2
    16'b11010000_01001111 : OUT <= 2;  //208 / 79 = 2
    16'b11010000_01010000 : OUT <= 2;  //208 / 80 = 2
    16'b11010000_01010001 : OUT <= 2;  //208 / 81 = 2
    16'b11010000_01010010 : OUT <= 2;  //208 / 82 = 2
    16'b11010000_01010011 : OUT <= 2;  //208 / 83 = 2
    16'b11010000_01010100 : OUT <= 2;  //208 / 84 = 2
    16'b11010000_01010101 : OUT <= 2;  //208 / 85 = 2
    16'b11010000_01010110 : OUT <= 2;  //208 / 86 = 2
    16'b11010000_01010111 : OUT <= 2;  //208 / 87 = 2
    16'b11010000_01011000 : OUT <= 2;  //208 / 88 = 2
    16'b11010000_01011001 : OUT <= 2;  //208 / 89 = 2
    16'b11010000_01011010 : OUT <= 2;  //208 / 90 = 2
    16'b11010000_01011011 : OUT <= 2;  //208 / 91 = 2
    16'b11010000_01011100 : OUT <= 2;  //208 / 92 = 2
    16'b11010000_01011101 : OUT <= 2;  //208 / 93 = 2
    16'b11010000_01011110 : OUT <= 2;  //208 / 94 = 2
    16'b11010000_01011111 : OUT <= 2;  //208 / 95 = 2
    16'b11010000_01100000 : OUT <= 2;  //208 / 96 = 2
    16'b11010000_01100001 : OUT <= 2;  //208 / 97 = 2
    16'b11010000_01100010 : OUT <= 2;  //208 / 98 = 2
    16'b11010000_01100011 : OUT <= 2;  //208 / 99 = 2
    16'b11010000_01100100 : OUT <= 2;  //208 / 100 = 2
    16'b11010000_01100101 : OUT <= 2;  //208 / 101 = 2
    16'b11010000_01100110 : OUT <= 2;  //208 / 102 = 2
    16'b11010000_01100111 : OUT <= 2;  //208 / 103 = 2
    16'b11010000_01101000 : OUT <= 2;  //208 / 104 = 2
    16'b11010000_01101001 : OUT <= 1;  //208 / 105 = 1
    16'b11010000_01101010 : OUT <= 1;  //208 / 106 = 1
    16'b11010000_01101011 : OUT <= 1;  //208 / 107 = 1
    16'b11010000_01101100 : OUT <= 1;  //208 / 108 = 1
    16'b11010000_01101101 : OUT <= 1;  //208 / 109 = 1
    16'b11010000_01101110 : OUT <= 1;  //208 / 110 = 1
    16'b11010000_01101111 : OUT <= 1;  //208 / 111 = 1
    16'b11010000_01110000 : OUT <= 1;  //208 / 112 = 1
    16'b11010000_01110001 : OUT <= 1;  //208 / 113 = 1
    16'b11010000_01110010 : OUT <= 1;  //208 / 114 = 1
    16'b11010000_01110011 : OUT <= 1;  //208 / 115 = 1
    16'b11010000_01110100 : OUT <= 1;  //208 / 116 = 1
    16'b11010000_01110101 : OUT <= 1;  //208 / 117 = 1
    16'b11010000_01110110 : OUT <= 1;  //208 / 118 = 1
    16'b11010000_01110111 : OUT <= 1;  //208 / 119 = 1
    16'b11010000_01111000 : OUT <= 1;  //208 / 120 = 1
    16'b11010000_01111001 : OUT <= 1;  //208 / 121 = 1
    16'b11010000_01111010 : OUT <= 1;  //208 / 122 = 1
    16'b11010000_01111011 : OUT <= 1;  //208 / 123 = 1
    16'b11010000_01111100 : OUT <= 1;  //208 / 124 = 1
    16'b11010000_01111101 : OUT <= 1;  //208 / 125 = 1
    16'b11010000_01111110 : OUT <= 1;  //208 / 126 = 1
    16'b11010000_01111111 : OUT <= 1;  //208 / 127 = 1
    16'b11010000_10000000 : OUT <= 1;  //208 / 128 = 1
    16'b11010000_10000001 : OUT <= 1;  //208 / 129 = 1
    16'b11010000_10000010 : OUT <= 1;  //208 / 130 = 1
    16'b11010000_10000011 : OUT <= 1;  //208 / 131 = 1
    16'b11010000_10000100 : OUT <= 1;  //208 / 132 = 1
    16'b11010000_10000101 : OUT <= 1;  //208 / 133 = 1
    16'b11010000_10000110 : OUT <= 1;  //208 / 134 = 1
    16'b11010000_10000111 : OUT <= 1;  //208 / 135 = 1
    16'b11010000_10001000 : OUT <= 1;  //208 / 136 = 1
    16'b11010000_10001001 : OUT <= 1;  //208 / 137 = 1
    16'b11010000_10001010 : OUT <= 1;  //208 / 138 = 1
    16'b11010000_10001011 : OUT <= 1;  //208 / 139 = 1
    16'b11010000_10001100 : OUT <= 1;  //208 / 140 = 1
    16'b11010000_10001101 : OUT <= 1;  //208 / 141 = 1
    16'b11010000_10001110 : OUT <= 1;  //208 / 142 = 1
    16'b11010000_10001111 : OUT <= 1;  //208 / 143 = 1
    16'b11010000_10010000 : OUT <= 1;  //208 / 144 = 1
    16'b11010000_10010001 : OUT <= 1;  //208 / 145 = 1
    16'b11010000_10010010 : OUT <= 1;  //208 / 146 = 1
    16'b11010000_10010011 : OUT <= 1;  //208 / 147 = 1
    16'b11010000_10010100 : OUT <= 1;  //208 / 148 = 1
    16'b11010000_10010101 : OUT <= 1;  //208 / 149 = 1
    16'b11010000_10010110 : OUT <= 1;  //208 / 150 = 1
    16'b11010000_10010111 : OUT <= 1;  //208 / 151 = 1
    16'b11010000_10011000 : OUT <= 1;  //208 / 152 = 1
    16'b11010000_10011001 : OUT <= 1;  //208 / 153 = 1
    16'b11010000_10011010 : OUT <= 1;  //208 / 154 = 1
    16'b11010000_10011011 : OUT <= 1;  //208 / 155 = 1
    16'b11010000_10011100 : OUT <= 1;  //208 / 156 = 1
    16'b11010000_10011101 : OUT <= 1;  //208 / 157 = 1
    16'b11010000_10011110 : OUT <= 1;  //208 / 158 = 1
    16'b11010000_10011111 : OUT <= 1;  //208 / 159 = 1
    16'b11010000_10100000 : OUT <= 1;  //208 / 160 = 1
    16'b11010000_10100001 : OUT <= 1;  //208 / 161 = 1
    16'b11010000_10100010 : OUT <= 1;  //208 / 162 = 1
    16'b11010000_10100011 : OUT <= 1;  //208 / 163 = 1
    16'b11010000_10100100 : OUT <= 1;  //208 / 164 = 1
    16'b11010000_10100101 : OUT <= 1;  //208 / 165 = 1
    16'b11010000_10100110 : OUT <= 1;  //208 / 166 = 1
    16'b11010000_10100111 : OUT <= 1;  //208 / 167 = 1
    16'b11010000_10101000 : OUT <= 1;  //208 / 168 = 1
    16'b11010000_10101001 : OUT <= 1;  //208 / 169 = 1
    16'b11010000_10101010 : OUT <= 1;  //208 / 170 = 1
    16'b11010000_10101011 : OUT <= 1;  //208 / 171 = 1
    16'b11010000_10101100 : OUT <= 1;  //208 / 172 = 1
    16'b11010000_10101101 : OUT <= 1;  //208 / 173 = 1
    16'b11010000_10101110 : OUT <= 1;  //208 / 174 = 1
    16'b11010000_10101111 : OUT <= 1;  //208 / 175 = 1
    16'b11010000_10110000 : OUT <= 1;  //208 / 176 = 1
    16'b11010000_10110001 : OUT <= 1;  //208 / 177 = 1
    16'b11010000_10110010 : OUT <= 1;  //208 / 178 = 1
    16'b11010000_10110011 : OUT <= 1;  //208 / 179 = 1
    16'b11010000_10110100 : OUT <= 1;  //208 / 180 = 1
    16'b11010000_10110101 : OUT <= 1;  //208 / 181 = 1
    16'b11010000_10110110 : OUT <= 1;  //208 / 182 = 1
    16'b11010000_10110111 : OUT <= 1;  //208 / 183 = 1
    16'b11010000_10111000 : OUT <= 1;  //208 / 184 = 1
    16'b11010000_10111001 : OUT <= 1;  //208 / 185 = 1
    16'b11010000_10111010 : OUT <= 1;  //208 / 186 = 1
    16'b11010000_10111011 : OUT <= 1;  //208 / 187 = 1
    16'b11010000_10111100 : OUT <= 1;  //208 / 188 = 1
    16'b11010000_10111101 : OUT <= 1;  //208 / 189 = 1
    16'b11010000_10111110 : OUT <= 1;  //208 / 190 = 1
    16'b11010000_10111111 : OUT <= 1;  //208 / 191 = 1
    16'b11010000_11000000 : OUT <= 1;  //208 / 192 = 1
    16'b11010000_11000001 : OUT <= 1;  //208 / 193 = 1
    16'b11010000_11000010 : OUT <= 1;  //208 / 194 = 1
    16'b11010000_11000011 : OUT <= 1;  //208 / 195 = 1
    16'b11010000_11000100 : OUT <= 1;  //208 / 196 = 1
    16'b11010000_11000101 : OUT <= 1;  //208 / 197 = 1
    16'b11010000_11000110 : OUT <= 1;  //208 / 198 = 1
    16'b11010000_11000111 : OUT <= 1;  //208 / 199 = 1
    16'b11010000_11001000 : OUT <= 1;  //208 / 200 = 1
    16'b11010000_11001001 : OUT <= 1;  //208 / 201 = 1
    16'b11010000_11001010 : OUT <= 1;  //208 / 202 = 1
    16'b11010000_11001011 : OUT <= 1;  //208 / 203 = 1
    16'b11010000_11001100 : OUT <= 1;  //208 / 204 = 1
    16'b11010000_11001101 : OUT <= 1;  //208 / 205 = 1
    16'b11010000_11001110 : OUT <= 1;  //208 / 206 = 1
    16'b11010000_11001111 : OUT <= 1;  //208 / 207 = 1
    16'b11010000_11010000 : OUT <= 1;  //208 / 208 = 1
    16'b11010000_11010001 : OUT <= 0;  //208 / 209 = 0
    16'b11010000_11010010 : OUT <= 0;  //208 / 210 = 0
    16'b11010000_11010011 : OUT <= 0;  //208 / 211 = 0
    16'b11010000_11010100 : OUT <= 0;  //208 / 212 = 0
    16'b11010000_11010101 : OUT <= 0;  //208 / 213 = 0
    16'b11010000_11010110 : OUT <= 0;  //208 / 214 = 0
    16'b11010000_11010111 : OUT <= 0;  //208 / 215 = 0
    16'b11010000_11011000 : OUT <= 0;  //208 / 216 = 0
    16'b11010000_11011001 : OUT <= 0;  //208 / 217 = 0
    16'b11010000_11011010 : OUT <= 0;  //208 / 218 = 0
    16'b11010000_11011011 : OUT <= 0;  //208 / 219 = 0
    16'b11010000_11011100 : OUT <= 0;  //208 / 220 = 0
    16'b11010000_11011101 : OUT <= 0;  //208 / 221 = 0
    16'b11010000_11011110 : OUT <= 0;  //208 / 222 = 0
    16'b11010000_11011111 : OUT <= 0;  //208 / 223 = 0
    16'b11010000_11100000 : OUT <= 0;  //208 / 224 = 0
    16'b11010000_11100001 : OUT <= 0;  //208 / 225 = 0
    16'b11010000_11100010 : OUT <= 0;  //208 / 226 = 0
    16'b11010000_11100011 : OUT <= 0;  //208 / 227 = 0
    16'b11010000_11100100 : OUT <= 0;  //208 / 228 = 0
    16'b11010000_11100101 : OUT <= 0;  //208 / 229 = 0
    16'b11010000_11100110 : OUT <= 0;  //208 / 230 = 0
    16'b11010000_11100111 : OUT <= 0;  //208 / 231 = 0
    16'b11010000_11101000 : OUT <= 0;  //208 / 232 = 0
    16'b11010000_11101001 : OUT <= 0;  //208 / 233 = 0
    16'b11010000_11101010 : OUT <= 0;  //208 / 234 = 0
    16'b11010000_11101011 : OUT <= 0;  //208 / 235 = 0
    16'b11010000_11101100 : OUT <= 0;  //208 / 236 = 0
    16'b11010000_11101101 : OUT <= 0;  //208 / 237 = 0
    16'b11010000_11101110 : OUT <= 0;  //208 / 238 = 0
    16'b11010000_11101111 : OUT <= 0;  //208 / 239 = 0
    16'b11010000_11110000 : OUT <= 0;  //208 / 240 = 0
    16'b11010000_11110001 : OUT <= 0;  //208 / 241 = 0
    16'b11010000_11110010 : OUT <= 0;  //208 / 242 = 0
    16'b11010000_11110011 : OUT <= 0;  //208 / 243 = 0
    16'b11010000_11110100 : OUT <= 0;  //208 / 244 = 0
    16'b11010000_11110101 : OUT <= 0;  //208 / 245 = 0
    16'b11010000_11110110 : OUT <= 0;  //208 / 246 = 0
    16'b11010000_11110111 : OUT <= 0;  //208 / 247 = 0
    16'b11010000_11111000 : OUT <= 0;  //208 / 248 = 0
    16'b11010000_11111001 : OUT <= 0;  //208 / 249 = 0
    16'b11010000_11111010 : OUT <= 0;  //208 / 250 = 0
    16'b11010000_11111011 : OUT <= 0;  //208 / 251 = 0
    16'b11010000_11111100 : OUT <= 0;  //208 / 252 = 0
    16'b11010000_11111101 : OUT <= 0;  //208 / 253 = 0
    16'b11010000_11111110 : OUT <= 0;  //208 / 254 = 0
    16'b11010000_11111111 : OUT <= 0;  //208 / 255 = 0
    16'b11010001_00000000 : OUT <= 0;  //209 / 0 = 0
    16'b11010001_00000001 : OUT <= 209;  //209 / 1 = 209
    16'b11010001_00000010 : OUT <= 104;  //209 / 2 = 104
    16'b11010001_00000011 : OUT <= 69;  //209 / 3 = 69
    16'b11010001_00000100 : OUT <= 52;  //209 / 4 = 52
    16'b11010001_00000101 : OUT <= 41;  //209 / 5 = 41
    16'b11010001_00000110 : OUT <= 34;  //209 / 6 = 34
    16'b11010001_00000111 : OUT <= 29;  //209 / 7 = 29
    16'b11010001_00001000 : OUT <= 26;  //209 / 8 = 26
    16'b11010001_00001001 : OUT <= 23;  //209 / 9 = 23
    16'b11010001_00001010 : OUT <= 20;  //209 / 10 = 20
    16'b11010001_00001011 : OUT <= 19;  //209 / 11 = 19
    16'b11010001_00001100 : OUT <= 17;  //209 / 12 = 17
    16'b11010001_00001101 : OUT <= 16;  //209 / 13 = 16
    16'b11010001_00001110 : OUT <= 14;  //209 / 14 = 14
    16'b11010001_00001111 : OUT <= 13;  //209 / 15 = 13
    16'b11010001_00010000 : OUT <= 13;  //209 / 16 = 13
    16'b11010001_00010001 : OUT <= 12;  //209 / 17 = 12
    16'b11010001_00010010 : OUT <= 11;  //209 / 18 = 11
    16'b11010001_00010011 : OUT <= 11;  //209 / 19 = 11
    16'b11010001_00010100 : OUT <= 10;  //209 / 20 = 10
    16'b11010001_00010101 : OUT <= 9;  //209 / 21 = 9
    16'b11010001_00010110 : OUT <= 9;  //209 / 22 = 9
    16'b11010001_00010111 : OUT <= 9;  //209 / 23 = 9
    16'b11010001_00011000 : OUT <= 8;  //209 / 24 = 8
    16'b11010001_00011001 : OUT <= 8;  //209 / 25 = 8
    16'b11010001_00011010 : OUT <= 8;  //209 / 26 = 8
    16'b11010001_00011011 : OUT <= 7;  //209 / 27 = 7
    16'b11010001_00011100 : OUT <= 7;  //209 / 28 = 7
    16'b11010001_00011101 : OUT <= 7;  //209 / 29 = 7
    16'b11010001_00011110 : OUT <= 6;  //209 / 30 = 6
    16'b11010001_00011111 : OUT <= 6;  //209 / 31 = 6
    16'b11010001_00100000 : OUT <= 6;  //209 / 32 = 6
    16'b11010001_00100001 : OUT <= 6;  //209 / 33 = 6
    16'b11010001_00100010 : OUT <= 6;  //209 / 34 = 6
    16'b11010001_00100011 : OUT <= 5;  //209 / 35 = 5
    16'b11010001_00100100 : OUT <= 5;  //209 / 36 = 5
    16'b11010001_00100101 : OUT <= 5;  //209 / 37 = 5
    16'b11010001_00100110 : OUT <= 5;  //209 / 38 = 5
    16'b11010001_00100111 : OUT <= 5;  //209 / 39 = 5
    16'b11010001_00101000 : OUT <= 5;  //209 / 40 = 5
    16'b11010001_00101001 : OUT <= 5;  //209 / 41 = 5
    16'b11010001_00101010 : OUT <= 4;  //209 / 42 = 4
    16'b11010001_00101011 : OUT <= 4;  //209 / 43 = 4
    16'b11010001_00101100 : OUT <= 4;  //209 / 44 = 4
    16'b11010001_00101101 : OUT <= 4;  //209 / 45 = 4
    16'b11010001_00101110 : OUT <= 4;  //209 / 46 = 4
    16'b11010001_00101111 : OUT <= 4;  //209 / 47 = 4
    16'b11010001_00110000 : OUT <= 4;  //209 / 48 = 4
    16'b11010001_00110001 : OUT <= 4;  //209 / 49 = 4
    16'b11010001_00110010 : OUT <= 4;  //209 / 50 = 4
    16'b11010001_00110011 : OUT <= 4;  //209 / 51 = 4
    16'b11010001_00110100 : OUT <= 4;  //209 / 52 = 4
    16'b11010001_00110101 : OUT <= 3;  //209 / 53 = 3
    16'b11010001_00110110 : OUT <= 3;  //209 / 54 = 3
    16'b11010001_00110111 : OUT <= 3;  //209 / 55 = 3
    16'b11010001_00111000 : OUT <= 3;  //209 / 56 = 3
    16'b11010001_00111001 : OUT <= 3;  //209 / 57 = 3
    16'b11010001_00111010 : OUT <= 3;  //209 / 58 = 3
    16'b11010001_00111011 : OUT <= 3;  //209 / 59 = 3
    16'b11010001_00111100 : OUT <= 3;  //209 / 60 = 3
    16'b11010001_00111101 : OUT <= 3;  //209 / 61 = 3
    16'b11010001_00111110 : OUT <= 3;  //209 / 62 = 3
    16'b11010001_00111111 : OUT <= 3;  //209 / 63 = 3
    16'b11010001_01000000 : OUT <= 3;  //209 / 64 = 3
    16'b11010001_01000001 : OUT <= 3;  //209 / 65 = 3
    16'b11010001_01000010 : OUT <= 3;  //209 / 66 = 3
    16'b11010001_01000011 : OUT <= 3;  //209 / 67 = 3
    16'b11010001_01000100 : OUT <= 3;  //209 / 68 = 3
    16'b11010001_01000101 : OUT <= 3;  //209 / 69 = 3
    16'b11010001_01000110 : OUT <= 2;  //209 / 70 = 2
    16'b11010001_01000111 : OUT <= 2;  //209 / 71 = 2
    16'b11010001_01001000 : OUT <= 2;  //209 / 72 = 2
    16'b11010001_01001001 : OUT <= 2;  //209 / 73 = 2
    16'b11010001_01001010 : OUT <= 2;  //209 / 74 = 2
    16'b11010001_01001011 : OUT <= 2;  //209 / 75 = 2
    16'b11010001_01001100 : OUT <= 2;  //209 / 76 = 2
    16'b11010001_01001101 : OUT <= 2;  //209 / 77 = 2
    16'b11010001_01001110 : OUT <= 2;  //209 / 78 = 2
    16'b11010001_01001111 : OUT <= 2;  //209 / 79 = 2
    16'b11010001_01010000 : OUT <= 2;  //209 / 80 = 2
    16'b11010001_01010001 : OUT <= 2;  //209 / 81 = 2
    16'b11010001_01010010 : OUT <= 2;  //209 / 82 = 2
    16'b11010001_01010011 : OUT <= 2;  //209 / 83 = 2
    16'b11010001_01010100 : OUT <= 2;  //209 / 84 = 2
    16'b11010001_01010101 : OUT <= 2;  //209 / 85 = 2
    16'b11010001_01010110 : OUT <= 2;  //209 / 86 = 2
    16'b11010001_01010111 : OUT <= 2;  //209 / 87 = 2
    16'b11010001_01011000 : OUT <= 2;  //209 / 88 = 2
    16'b11010001_01011001 : OUT <= 2;  //209 / 89 = 2
    16'b11010001_01011010 : OUT <= 2;  //209 / 90 = 2
    16'b11010001_01011011 : OUT <= 2;  //209 / 91 = 2
    16'b11010001_01011100 : OUT <= 2;  //209 / 92 = 2
    16'b11010001_01011101 : OUT <= 2;  //209 / 93 = 2
    16'b11010001_01011110 : OUT <= 2;  //209 / 94 = 2
    16'b11010001_01011111 : OUT <= 2;  //209 / 95 = 2
    16'b11010001_01100000 : OUT <= 2;  //209 / 96 = 2
    16'b11010001_01100001 : OUT <= 2;  //209 / 97 = 2
    16'b11010001_01100010 : OUT <= 2;  //209 / 98 = 2
    16'b11010001_01100011 : OUT <= 2;  //209 / 99 = 2
    16'b11010001_01100100 : OUT <= 2;  //209 / 100 = 2
    16'b11010001_01100101 : OUT <= 2;  //209 / 101 = 2
    16'b11010001_01100110 : OUT <= 2;  //209 / 102 = 2
    16'b11010001_01100111 : OUT <= 2;  //209 / 103 = 2
    16'b11010001_01101000 : OUT <= 2;  //209 / 104 = 2
    16'b11010001_01101001 : OUT <= 1;  //209 / 105 = 1
    16'b11010001_01101010 : OUT <= 1;  //209 / 106 = 1
    16'b11010001_01101011 : OUT <= 1;  //209 / 107 = 1
    16'b11010001_01101100 : OUT <= 1;  //209 / 108 = 1
    16'b11010001_01101101 : OUT <= 1;  //209 / 109 = 1
    16'b11010001_01101110 : OUT <= 1;  //209 / 110 = 1
    16'b11010001_01101111 : OUT <= 1;  //209 / 111 = 1
    16'b11010001_01110000 : OUT <= 1;  //209 / 112 = 1
    16'b11010001_01110001 : OUT <= 1;  //209 / 113 = 1
    16'b11010001_01110010 : OUT <= 1;  //209 / 114 = 1
    16'b11010001_01110011 : OUT <= 1;  //209 / 115 = 1
    16'b11010001_01110100 : OUT <= 1;  //209 / 116 = 1
    16'b11010001_01110101 : OUT <= 1;  //209 / 117 = 1
    16'b11010001_01110110 : OUT <= 1;  //209 / 118 = 1
    16'b11010001_01110111 : OUT <= 1;  //209 / 119 = 1
    16'b11010001_01111000 : OUT <= 1;  //209 / 120 = 1
    16'b11010001_01111001 : OUT <= 1;  //209 / 121 = 1
    16'b11010001_01111010 : OUT <= 1;  //209 / 122 = 1
    16'b11010001_01111011 : OUT <= 1;  //209 / 123 = 1
    16'b11010001_01111100 : OUT <= 1;  //209 / 124 = 1
    16'b11010001_01111101 : OUT <= 1;  //209 / 125 = 1
    16'b11010001_01111110 : OUT <= 1;  //209 / 126 = 1
    16'b11010001_01111111 : OUT <= 1;  //209 / 127 = 1
    16'b11010001_10000000 : OUT <= 1;  //209 / 128 = 1
    16'b11010001_10000001 : OUT <= 1;  //209 / 129 = 1
    16'b11010001_10000010 : OUT <= 1;  //209 / 130 = 1
    16'b11010001_10000011 : OUT <= 1;  //209 / 131 = 1
    16'b11010001_10000100 : OUT <= 1;  //209 / 132 = 1
    16'b11010001_10000101 : OUT <= 1;  //209 / 133 = 1
    16'b11010001_10000110 : OUT <= 1;  //209 / 134 = 1
    16'b11010001_10000111 : OUT <= 1;  //209 / 135 = 1
    16'b11010001_10001000 : OUT <= 1;  //209 / 136 = 1
    16'b11010001_10001001 : OUT <= 1;  //209 / 137 = 1
    16'b11010001_10001010 : OUT <= 1;  //209 / 138 = 1
    16'b11010001_10001011 : OUT <= 1;  //209 / 139 = 1
    16'b11010001_10001100 : OUT <= 1;  //209 / 140 = 1
    16'b11010001_10001101 : OUT <= 1;  //209 / 141 = 1
    16'b11010001_10001110 : OUT <= 1;  //209 / 142 = 1
    16'b11010001_10001111 : OUT <= 1;  //209 / 143 = 1
    16'b11010001_10010000 : OUT <= 1;  //209 / 144 = 1
    16'b11010001_10010001 : OUT <= 1;  //209 / 145 = 1
    16'b11010001_10010010 : OUT <= 1;  //209 / 146 = 1
    16'b11010001_10010011 : OUT <= 1;  //209 / 147 = 1
    16'b11010001_10010100 : OUT <= 1;  //209 / 148 = 1
    16'b11010001_10010101 : OUT <= 1;  //209 / 149 = 1
    16'b11010001_10010110 : OUT <= 1;  //209 / 150 = 1
    16'b11010001_10010111 : OUT <= 1;  //209 / 151 = 1
    16'b11010001_10011000 : OUT <= 1;  //209 / 152 = 1
    16'b11010001_10011001 : OUT <= 1;  //209 / 153 = 1
    16'b11010001_10011010 : OUT <= 1;  //209 / 154 = 1
    16'b11010001_10011011 : OUT <= 1;  //209 / 155 = 1
    16'b11010001_10011100 : OUT <= 1;  //209 / 156 = 1
    16'b11010001_10011101 : OUT <= 1;  //209 / 157 = 1
    16'b11010001_10011110 : OUT <= 1;  //209 / 158 = 1
    16'b11010001_10011111 : OUT <= 1;  //209 / 159 = 1
    16'b11010001_10100000 : OUT <= 1;  //209 / 160 = 1
    16'b11010001_10100001 : OUT <= 1;  //209 / 161 = 1
    16'b11010001_10100010 : OUT <= 1;  //209 / 162 = 1
    16'b11010001_10100011 : OUT <= 1;  //209 / 163 = 1
    16'b11010001_10100100 : OUT <= 1;  //209 / 164 = 1
    16'b11010001_10100101 : OUT <= 1;  //209 / 165 = 1
    16'b11010001_10100110 : OUT <= 1;  //209 / 166 = 1
    16'b11010001_10100111 : OUT <= 1;  //209 / 167 = 1
    16'b11010001_10101000 : OUT <= 1;  //209 / 168 = 1
    16'b11010001_10101001 : OUT <= 1;  //209 / 169 = 1
    16'b11010001_10101010 : OUT <= 1;  //209 / 170 = 1
    16'b11010001_10101011 : OUT <= 1;  //209 / 171 = 1
    16'b11010001_10101100 : OUT <= 1;  //209 / 172 = 1
    16'b11010001_10101101 : OUT <= 1;  //209 / 173 = 1
    16'b11010001_10101110 : OUT <= 1;  //209 / 174 = 1
    16'b11010001_10101111 : OUT <= 1;  //209 / 175 = 1
    16'b11010001_10110000 : OUT <= 1;  //209 / 176 = 1
    16'b11010001_10110001 : OUT <= 1;  //209 / 177 = 1
    16'b11010001_10110010 : OUT <= 1;  //209 / 178 = 1
    16'b11010001_10110011 : OUT <= 1;  //209 / 179 = 1
    16'b11010001_10110100 : OUT <= 1;  //209 / 180 = 1
    16'b11010001_10110101 : OUT <= 1;  //209 / 181 = 1
    16'b11010001_10110110 : OUT <= 1;  //209 / 182 = 1
    16'b11010001_10110111 : OUT <= 1;  //209 / 183 = 1
    16'b11010001_10111000 : OUT <= 1;  //209 / 184 = 1
    16'b11010001_10111001 : OUT <= 1;  //209 / 185 = 1
    16'b11010001_10111010 : OUT <= 1;  //209 / 186 = 1
    16'b11010001_10111011 : OUT <= 1;  //209 / 187 = 1
    16'b11010001_10111100 : OUT <= 1;  //209 / 188 = 1
    16'b11010001_10111101 : OUT <= 1;  //209 / 189 = 1
    16'b11010001_10111110 : OUT <= 1;  //209 / 190 = 1
    16'b11010001_10111111 : OUT <= 1;  //209 / 191 = 1
    16'b11010001_11000000 : OUT <= 1;  //209 / 192 = 1
    16'b11010001_11000001 : OUT <= 1;  //209 / 193 = 1
    16'b11010001_11000010 : OUT <= 1;  //209 / 194 = 1
    16'b11010001_11000011 : OUT <= 1;  //209 / 195 = 1
    16'b11010001_11000100 : OUT <= 1;  //209 / 196 = 1
    16'b11010001_11000101 : OUT <= 1;  //209 / 197 = 1
    16'b11010001_11000110 : OUT <= 1;  //209 / 198 = 1
    16'b11010001_11000111 : OUT <= 1;  //209 / 199 = 1
    16'b11010001_11001000 : OUT <= 1;  //209 / 200 = 1
    16'b11010001_11001001 : OUT <= 1;  //209 / 201 = 1
    16'b11010001_11001010 : OUT <= 1;  //209 / 202 = 1
    16'b11010001_11001011 : OUT <= 1;  //209 / 203 = 1
    16'b11010001_11001100 : OUT <= 1;  //209 / 204 = 1
    16'b11010001_11001101 : OUT <= 1;  //209 / 205 = 1
    16'b11010001_11001110 : OUT <= 1;  //209 / 206 = 1
    16'b11010001_11001111 : OUT <= 1;  //209 / 207 = 1
    16'b11010001_11010000 : OUT <= 1;  //209 / 208 = 1
    16'b11010001_11010001 : OUT <= 1;  //209 / 209 = 1
    16'b11010001_11010010 : OUT <= 0;  //209 / 210 = 0
    16'b11010001_11010011 : OUT <= 0;  //209 / 211 = 0
    16'b11010001_11010100 : OUT <= 0;  //209 / 212 = 0
    16'b11010001_11010101 : OUT <= 0;  //209 / 213 = 0
    16'b11010001_11010110 : OUT <= 0;  //209 / 214 = 0
    16'b11010001_11010111 : OUT <= 0;  //209 / 215 = 0
    16'b11010001_11011000 : OUT <= 0;  //209 / 216 = 0
    16'b11010001_11011001 : OUT <= 0;  //209 / 217 = 0
    16'b11010001_11011010 : OUT <= 0;  //209 / 218 = 0
    16'b11010001_11011011 : OUT <= 0;  //209 / 219 = 0
    16'b11010001_11011100 : OUT <= 0;  //209 / 220 = 0
    16'b11010001_11011101 : OUT <= 0;  //209 / 221 = 0
    16'b11010001_11011110 : OUT <= 0;  //209 / 222 = 0
    16'b11010001_11011111 : OUT <= 0;  //209 / 223 = 0
    16'b11010001_11100000 : OUT <= 0;  //209 / 224 = 0
    16'b11010001_11100001 : OUT <= 0;  //209 / 225 = 0
    16'b11010001_11100010 : OUT <= 0;  //209 / 226 = 0
    16'b11010001_11100011 : OUT <= 0;  //209 / 227 = 0
    16'b11010001_11100100 : OUT <= 0;  //209 / 228 = 0
    16'b11010001_11100101 : OUT <= 0;  //209 / 229 = 0
    16'b11010001_11100110 : OUT <= 0;  //209 / 230 = 0
    16'b11010001_11100111 : OUT <= 0;  //209 / 231 = 0
    16'b11010001_11101000 : OUT <= 0;  //209 / 232 = 0
    16'b11010001_11101001 : OUT <= 0;  //209 / 233 = 0
    16'b11010001_11101010 : OUT <= 0;  //209 / 234 = 0
    16'b11010001_11101011 : OUT <= 0;  //209 / 235 = 0
    16'b11010001_11101100 : OUT <= 0;  //209 / 236 = 0
    16'b11010001_11101101 : OUT <= 0;  //209 / 237 = 0
    16'b11010001_11101110 : OUT <= 0;  //209 / 238 = 0
    16'b11010001_11101111 : OUT <= 0;  //209 / 239 = 0
    16'b11010001_11110000 : OUT <= 0;  //209 / 240 = 0
    16'b11010001_11110001 : OUT <= 0;  //209 / 241 = 0
    16'b11010001_11110010 : OUT <= 0;  //209 / 242 = 0
    16'b11010001_11110011 : OUT <= 0;  //209 / 243 = 0
    16'b11010001_11110100 : OUT <= 0;  //209 / 244 = 0
    16'b11010001_11110101 : OUT <= 0;  //209 / 245 = 0
    16'b11010001_11110110 : OUT <= 0;  //209 / 246 = 0
    16'b11010001_11110111 : OUT <= 0;  //209 / 247 = 0
    16'b11010001_11111000 : OUT <= 0;  //209 / 248 = 0
    16'b11010001_11111001 : OUT <= 0;  //209 / 249 = 0
    16'b11010001_11111010 : OUT <= 0;  //209 / 250 = 0
    16'b11010001_11111011 : OUT <= 0;  //209 / 251 = 0
    16'b11010001_11111100 : OUT <= 0;  //209 / 252 = 0
    16'b11010001_11111101 : OUT <= 0;  //209 / 253 = 0
    16'b11010001_11111110 : OUT <= 0;  //209 / 254 = 0
    16'b11010001_11111111 : OUT <= 0;  //209 / 255 = 0
    16'b11010010_00000000 : OUT <= 0;  //210 / 0 = 0
    16'b11010010_00000001 : OUT <= 210;  //210 / 1 = 210
    16'b11010010_00000010 : OUT <= 105;  //210 / 2 = 105
    16'b11010010_00000011 : OUT <= 70;  //210 / 3 = 70
    16'b11010010_00000100 : OUT <= 52;  //210 / 4 = 52
    16'b11010010_00000101 : OUT <= 42;  //210 / 5 = 42
    16'b11010010_00000110 : OUT <= 35;  //210 / 6 = 35
    16'b11010010_00000111 : OUT <= 30;  //210 / 7 = 30
    16'b11010010_00001000 : OUT <= 26;  //210 / 8 = 26
    16'b11010010_00001001 : OUT <= 23;  //210 / 9 = 23
    16'b11010010_00001010 : OUT <= 21;  //210 / 10 = 21
    16'b11010010_00001011 : OUT <= 19;  //210 / 11 = 19
    16'b11010010_00001100 : OUT <= 17;  //210 / 12 = 17
    16'b11010010_00001101 : OUT <= 16;  //210 / 13 = 16
    16'b11010010_00001110 : OUT <= 15;  //210 / 14 = 15
    16'b11010010_00001111 : OUT <= 14;  //210 / 15 = 14
    16'b11010010_00010000 : OUT <= 13;  //210 / 16 = 13
    16'b11010010_00010001 : OUT <= 12;  //210 / 17 = 12
    16'b11010010_00010010 : OUT <= 11;  //210 / 18 = 11
    16'b11010010_00010011 : OUT <= 11;  //210 / 19 = 11
    16'b11010010_00010100 : OUT <= 10;  //210 / 20 = 10
    16'b11010010_00010101 : OUT <= 10;  //210 / 21 = 10
    16'b11010010_00010110 : OUT <= 9;  //210 / 22 = 9
    16'b11010010_00010111 : OUT <= 9;  //210 / 23 = 9
    16'b11010010_00011000 : OUT <= 8;  //210 / 24 = 8
    16'b11010010_00011001 : OUT <= 8;  //210 / 25 = 8
    16'b11010010_00011010 : OUT <= 8;  //210 / 26 = 8
    16'b11010010_00011011 : OUT <= 7;  //210 / 27 = 7
    16'b11010010_00011100 : OUT <= 7;  //210 / 28 = 7
    16'b11010010_00011101 : OUT <= 7;  //210 / 29 = 7
    16'b11010010_00011110 : OUT <= 7;  //210 / 30 = 7
    16'b11010010_00011111 : OUT <= 6;  //210 / 31 = 6
    16'b11010010_00100000 : OUT <= 6;  //210 / 32 = 6
    16'b11010010_00100001 : OUT <= 6;  //210 / 33 = 6
    16'b11010010_00100010 : OUT <= 6;  //210 / 34 = 6
    16'b11010010_00100011 : OUT <= 6;  //210 / 35 = 6
    16'b11010010_00100100 : OUT <= 5;  //210 / 36 = 5
    16'b11010010_00100101 : OUT <= 5;  //210 / 37 = 5
    16'b11010010_00100110 : OUT <= 5;  //210 / 38 = 5
    16'b11010010_00100111 : OUT <= 5;  //210 / 39 = 5
    16'b11010010_00101000 : OUT <= 5;  //210 / 40 = 5
    16'b11010010_00101001 : OUT <= 5;  //210 / 41 = 5
    16'b11010010_00101010 : OUT <= 5;  //210 / 42 = 5
    16'b11010010_00101011 : OUT <= 4;  //210 / 43 = 4
    16'b11010010_00101100 : OUT <= 4;  //210 / 44 = 4
    16'b11010010_00101101 : OUT <= 4;  //210 / 45 = 4
    16'b11010010_00101110 : OUT <= 4;  //210 / 46 = 4
    16'b11010010_00101111 : OUT <= 4;  //210 / 47 = 4
    16'b11010010_00110000 : OUT <= 4;  //210 / 48 = 4
    16'b11010010_00110001 : OUT <= 4;  //210 / 49 = 4
    16'b11010010_00110010 : OUT <= 4;  //210 / 50 = 4
    16'b11010010_00110011 : OUT <= 4;  //210 / 51 = 4
    16'b11010010_00110100 : OUT <= 4;  //210 / 52 = 4
    16'b11010010_00110101 : OUT <= 3;  //210 / 53 = 3
    16'b11010010_00110110 : OUT <= 3;  //210 / 54 = 3
    16'b11010010_00110111 : OUT <= 3;  //210 / 55 = 3
    16'b11010010_00111000 : OUT <= 3;  //210 / 56 = 3
    16'b11010010_00111001 : OUT <= 3;  //210 / 57 = 3
    16'b11010010_00111010 : OUT <= 3;  //210 / 58 = 3
    16'b11010010_00111011 : OUT <= 3;  //210 / 59 = 3
    16'b11010010_00111100 : OUT <= 3;  //210 / 60 = 3
    16'b11010010_00111101 : OUT <= 3;  //210 / 61 = 3
    16'b11010010_00111110 : OUT <= 3;  //210 / 62 = 3
    16'b11010010_00111111 : OUT <= 3;  //210 / 63 = 3
    16'b11010010_01000000 : OUT <= 3;  //210 / 64 = 3
    16'b11010010_01000001 : OUT <= 3;  //210 / 65 = 3
    16'b11010010_01000010 : OUT <= 3;  //210 / 66 = 3
    16'b11010010_01000011 : OUT <= 3;  //210 / 67 = 3
    16'b11010010_01000100 : OUT <= 3;  //210 / 68 = 3
    16'b11010010_01000101 : OUT <= 3;  //210 / 69 = 3
    16'b11010010_01000110 : OUT <= 3;  //210 / 70 = 3
    16'b11010010_01000111 : OUT <= 2;  //210 / 71 = 2
    16'b11010010_01001000 : OUT <= 2;  //210 / 72 = 2
    16'b11010010_01001001 : OUT <= 2;  //210 / 73 = 2
    16'b11010010_01001010 : OUT <= 2;  //210 / 74 = 2
    16'b11010010_01001011 : OUT <= 2;  //210 / 75 = 2
    16'b11010010_01001100 : OUT <= 2;  //210 / 76 = 2
    16'b11010010_01001101 : OUT <= 2;  //210 / 77 = 2
    16'b11010010_01001110 : OUT <= 2;  //210 / 78 = 2
    16'b11010010_01001111 : OUT <= 2;  //210 / 79 = 2
    16'b11010010_01010000 : OUT <= 2;  //210 / 80 = 2
    16'b11010010_01010001 : OUT <= 2;  //210 / 81 = 2
    16'b11010010_01010010 : OUT <= 2;  //210 / 82 = 2
    16'b11010010_01010011 : OUT <= 2;  //210 / 83 = 2
    16'b11010010_01010100 : OUT <= 2;  //210 / 84 = 2
    16'b11010010_01010101 : OUT <= 2;  //210 / 85 = 2
    16'b11010010_01010110 : OUT <= 2;  //210 / 86 = 2
    16'b11010010_01010111 : OUT <= 2;  //210 / 87 = 2
    16'b11010010_01011000 : OUT <= 2;  //210 / 88 = 2
    16'b11010010_01011001 : OUT <= 2;  //210 / 89 = 2
    16'b11010010_01011010 : OUT <= 2;  //210 / 90 = 2
    16'b11010010_01011011 : OUT <= 2;  //210 / 91 = 2
    16'b11010010_01011100 : OUT <= 2;  //210 / 92 = 2
    16'b11010010_01011101 : OUT <= 2;  //210 / 93 = 2
    16'b11010010_01011110 : OUT <= 2;  //210 / 94 = 2
    16'b11010010_01011111 : OUT <= 2;  //210 / 95 = 2
    16'b11010010_01100000 : OUT <= 2;  //210 / 96 = 2
    16'b11010010_01100001 : OUT <= 2;  //210 / 97 = 2
    16'b11010010_01100010 : OUT <= 2;  //210 / 98 = 2
    16'b11010010_01100011 : OUT <= 2;  //210 / 99 = 2
    16'b11010010_01100100 : OUT <= 2;  //210 / 100 = 2
    16'b11010010_01100101 : OUT <= 2;  //210 / 101 = 2
    16'b11010010_01100110 : OUT <= 2;  //210 / 102 = 2
    16'b11010010_01100111 : OUT <= 2;  //210 / 103 = 2
    16'b11010010_01101000 : OUT <= 2;  //210 / 104 = 2
    16'b11010010_01101001 : OUT <= 2;  //210 / 105 = 2
    16'b11010010_01101010 : OUT <= 1;  //210 / 106 = 1
    16'b11010010_01101011 : OUT <= 1;  //210 / 107 = 1
    16'b11010010_01101100 : OUT <= 1;  //210 / 108 = 1
    16'b11010010_01101101 : OUT <= 1;  //210 / 109 = 1
    16'b11010010_01101110 : OUT <= 1;  //210 / 110 = 1
    16'b11010010_01101111 : OUT <= 1;  //210 / 111 = 1
    16'b11010010_01110000 : OUT <= 1;  //210 / 112 = 1
    16'b11010010_01110001 : OUT <= 1;  //210 / 113 = 1
    16'b11010010_01110010 : OUT <= 1;  //210 / 114 = 1
    16'b11010010_01110011 : OUT <= 1;  //210 / 115 = 1
    16'b11010010_01110100 : OUT <= 1;  //210 / 116 = 1
    16'b11010010_01110101 : OUT <= 1;  //210 / 117 = 1
    16'b11010010_01110110 : OUT <= 1;  //210 / 118 = 1
    16'b11010010_01110111 : OUT <= 1;  //210 / 119 = 1
    16'b11010010_01111000 : OUT <= 1;  //210 / 120 = 1
    16'b11010010_01111001 : OUT <= 1;  //210 / 121 = 1
    16'b11010010_01111010 : OUT <= 1;  //210 / 122 = 1
    16'b11010010_01111011 : OUT <= 1;  //210 / 123 = 1
    16'b11010010_01111100 : OUT <= 1;  //210 / 124 = 1
    16'b11010010_01111101 : OUT <= 1;  //210 / 125 = 1
    16'b11010010_01111110 : OUT <= 1;  //210 / 126 = 1
    16'b11010010_01111111 : OUT <= 1;  //210 / 127 = 1
    16'b11010010_10000000 : OUT <= 1;  //210 / 128 = 1
    16'b11010010_10000001 : OUT <= 1;  //210 / 129 = 1
    16'b11010010_10000010 : OUT <= 1;  //210 / 130 = 1
    16'b11010010_10000011 : OUT <= 1;  //210 / 131 = 1
    16'b11010010_10000100 : OUT <= 1;  //210 / 132 = 1
    16'b11010010_10000101 : OUT <= 1;  //210 / 133 = 1
    16'b11010010_10000110 : OUT <= 1;  //210 / 134 = 1
    16'b11010010_10000111 : OUT <= 1;  //210 / 135 = 1
    16'b11010010_10001000 : OUT <= 1;  //210 / 136 = 1
    16'b11010010_10001001 : OUT <= 1;  //210 / 137 = 1
    16'b11010010_10001010 : OUT <= 1;  //210 / 138 = 1
    16'b11010010_10001011 : OUT <= 1;  //210 / 139 = 1
    16'b11010010_10001100 : OUT <= 1;  //210 / 140 = 1
    16'b11010010_10001101 : OUT <= 1;  //210 / 141 = 1
    16'b11010010_10001110 : OUT <= 1;  //210 / 142 = 1
    16'b11010010_10001111 : OUT <= 1;  //210 / 143 = 1
    16'b11010010_10010000 : OUT <= 1;  //210 / 144 = 1
    16'b11010010_10010001 : OUT <= 1;  //210 / 145 = 1
    16'b11010010_10010010 : OUT <= 1;  //210 / 146 = 1
    16'b11010010_10010011 : OUT <= 1;  //210 / 147 = 1
    16'b11010010_10010100 : OUT <= 1;  //210 / 148 = 1
    16'b11010010_10010101 : OUT <= 1;  //210 / 149 = 1
    16'b11010010_10010110 : OUT <= 1;  //210 / 150 = 1
    16'b11010010_10010111 : OUT <= 1;  //210 / 151 = 1
    16'b11010010_10011000 : OUT <= 1;  //210 / 152 = 1
    16'b11010010_10011001 : OUT <= 1;  //210 / 153 = 1
    16'b11010010_10011010 : OUT <= 1;  //210 / 154 = 1
    16'b11010010_10011011 : OUT <= 1;  //210 / 155 = 1
    16'b11010010_10011100 : OUT <= 1;  //210 / 156 = 1
    16'b11010010_10011101 : OUT <= 1;  //210 / 157 = 1
    16'b11010010_10011110 : OUT <= 1;  //210 / 158 = 1
    16'b11010010_10011111 : OUT <= 1;  //210 / 159 = 1
    16'b11010010_10100000 : OUT <= 1;  //210 / 160 = 1
    16'b11010010_10100001 : OUT <= 1;  //210 / 161 = 1
    16'b11010010_10100010 : OUT <= 1;  //210 / 162 = 1
    16'b11010010_10100011 : OUT <= 1;  //210 / 163 = 1
    16'b11010010_10100100 : OUT <= 1;  //210 / 164 = 1
    16'b11010010_10100101 : OUT <= 1;  //210 / 165 = 1
    16'b11010010_10100110 : OUT <= 1;  //210 / 166 = 1
    16'b11010010_10100111 : OUT <= 1;  //210 / 167 = 1
    16'b11010010_10101000 : OUT <= 1;  //210 / 168 = 1
    16'b11010010_10101001 : OUT <= 1;  //210 / 169 = 1
    16'b11010010_10101010 : OUT <= 1;  //210 / 170 = 1
    16'b11010010_10101011 : OUT <= 1;  //210 / 171 = 1
    16'b11010010_10101100 : OUT <= 1;  //210 / 172 = 1
    16'b11010010_10101101 : OUT <= 1;  //210 / 173 = 1
    16'b11010010_10101110 : OUT <= 1;  //210 / 174 = 1
    16'b11010010_10101111 : OUT <= 1;  //210 / 175 = 1
    16'b11010010_10110000 : OUT <= 1;  //210 / 176 = 1
    16'b11010010_10110001 : OUT <= 1;  //210 / 177 = 1
    16'b11010010_10110010 : OUT <= 1;  //210 / 178 = 1
    16'b11010010_10110011 : OUT <= 1;  //210 / 179 = 1
    16'b11010010_10110100 : OUT <= 1;  //210 / 180 = 1
    16'b11010010_10110101 : OUT <= 1;  //210 / 181 = 1
    16'b11010010_10110110 : OUT <= 1;  //210 / 182 = 1
    16'b11010010_10110111 : OUT <= 1;  //210 / 183 = 1
    16'b11010010_10111000 : OUT <= 1;  //210 / 184 = 1
    16'b11010010_10111001 : OUT <= 1;  //210 / 185 = 1
    16'b11010010_10111010 : OUT <= 1;  //210 / 186 = 1
    16'b11010010_10111011 : OUT <= 1;  //210 / 187 = 1
    16'b11010010_10111100 : OUT <= 1;  //210 / 188 = 1
    16'b11010010_10111101 : OUT <= 1;  //210 / 189 = 1
    16'b11010010_10111110 : OUT <= 1;  //210 / 190 = 1
    16'b11010010_10111111 : OUT <= 1;  //210 / 191 = 1
    16'b11010010_11000000 : OUT <= 1;  //210 / 192 = 1
    16'b11010010_11000001 : OUT <= 1;  //210 / 193 = 1
    16'b11010010_11000010 : OUT <= 1;  //210 / 194 = 1
    16'b11010010_11000011 : OUT <= 1;  //210 / 195 = 1
    16'b11010010_11000100 : OUT <= 1;  //210 / 196 = 1
    16'b11010010_11000101 : OUT <= 1;  //210 / 197 = 1
    16'b11010010_11000110 : OUT <= 1;  //210 / 198 = 1
    16'b11010010_11000111 : OUT <= 1;  //210 / 199 = 1
    16'b11010010_11001000 : OUT <= 1;  //210 / 200 = 1
    16'b11010010_11001001 : OUT <= 1;  //210 / 201 = 1
    16'b11010010_11001010 : OUT <= 1;  //210 / 202 = 1
    16'b11010010_11001011 : OUT <= 1;  //210 / 203 = 1
    16'b11010010_11001100 : OUT <= 1;  //210 / 204 = 1
    16'b11010010_11001101 : OUT <= 1;  //210 / 205 = 1
    16'b11010010_11001110 : OUT <= 1;  //210 / 206 = 1
    16'b11010010_11001111 : OUT <= 1;  //210 / 207 = 1
    16'b11010010_11010000 : OUT <= 1;  //210 / 208 = 1
    16'b11010010_11010001 : OUT <= 1;  //210 / 209 = 1
    16'b11010010_11010010 : OUT <= 1;  //210 / 210 = 1
    16'b11010010_11010011 : OUT <= 0;  //210 / 211 = 0
    16'b11010010_11010100 : OUT <= 0;  //210 / 212 = 0
    16'b11010010_11010101 : OUT <= 0;  //210 / 213 = 0
    16'b11010010_11010110 : OUT <= 0;  //210 / 214 = 0
    16'b11010010_11010111 : OUT <= 0;  //210 / 215 = 0
    16'b11010010_11011000 : OUT <= 0;  //210 / 216 = 0
    16'b11010010_11011001 : OUT <= 0;  //210 / 217 = 0
    16'b11010010_11011010 : OUT <= 0;  //210 / 218 = 0
    16'b11010010_11011011 : OUT <= 0;  //210 / 219 = 0
    16'b11010010_11011100 : OUT <= 0;  //210 / 220 = 0
    16'b11010010_11011101 : OUT <= 0;  //210 / 221 = 0
    16'b11010010_11011110 : OUT <= 0;  //210 / 222 = 0
    16'b11010010_11011111 : OUT <= 0;  //210 / 223 = 0
    16'b11010010_11100000 : OUT <= 0;  //210 / 224 = 0
    16'b11010010_11100001 : OUT <= 0;  //210 / 225 = 0
    16'b11010010_11100010 : OUT <= 0;  //210 / 226 = 0
    16'b11010010_11100011 : OUT <= 0;  //210 / 227 = 0
    16'b11010010_11100100 : OUT <= 0;  //210 / 228 = 0
    16'b11010010_11100101 : OUT <= 0;  //210 / 229 = 0
    16'b11010010_11100110 : OUT <= 0;  //210 / 230 = 0
    16'b11010010_11100111 : OUT <= 0;  //210 / 231 = 0
    16'b11010010_11101000 : OUT <= 0;  //210 / 232 = 0
    16'b11010010_11101001 : OUT <= 0;  //210 / 233 = 0
    16'b11010010_11101010 : OUT <= 0;  //210 / 234 = 0
    16'b11010010_11101011 : OUT <= 0;  //210 / 235 = 0
    16'b11010010_11101100 : OUT <= 0;  //210 / 236 = 0
    16'b11010010_11101101 : OUT <= 0;  //210 / 237 = 0
    16'b11010010_11101110 : OUT <= 0;  //210 / 238 = 0
    16'b11010010_11101111 : OUT <= 0;  //210 / 239 = 0
    16'b11010010_11110000 : OUT <= 0;  //210 / 240 = 0
    16'b11010010_11110001 : OUT <= 0;  //210 / 241 = 0
    16'b11010010_11110010 : OUT <= 0;  //210 / 242 = 0
    16'b11010010_11110011 : OUT <= 0;  //210 / 243 = 0
    16'b11010010_11110100 : OUT <= 0;  //210 / 244 = 0
    16'b11010010_11110101 : OUT <= 0;  //210 / 245 = 0
    16'b11010010_11110110 : OUT <= 0;  //210 / 246 = 0
    16'b11010010_11110111 : OUT <= 0;  //210 / 247 = 0
    16'b11010010_11111000 : OUT <= 0;  //210 / 248 = 0
    16'b11010010_11111001 : OUT <= 0;  //210 / 249 = 0
    16'b11010010_11111010 : OUT <= 0;  //210 / 250 = 0
    16'b11010010_11111011 : OUT <= 0;  //210 / 251 = 0
    16'b11010010_11111100 : OUT <= 0;  //210 / 252 = 0
    16'b11010010_11111101 : OUT <= 0;  //210 / 253 = 0
    16'b11010010_11111110 : OUT <= 0;  //210 / 254 = 0
    16'b11010010_11111111 : OUT <= 0;  //210 / 255 = 0
    16'b11010011_00000000 : OUT <= 0;  //211 / 0 = 0
    16'b11010011_00000001 : OUT <= 211;  //211 / 1 = 211
    16'b11010011_00000010 : OUT <= 105;  //211 / 2 = 105
    16'b11010011_00000011 : OUT <= 70;  //211 / 3 = 70
    16'b11010011_00000100 : OUT <= 52;  //211 / 4 = 52
    16'b11010011_00000101 : OUT <= 42;  //211 / 5 = 42
    16'b11010011_00000110 : OUT <= 35;  //211 / 6 = 35
    16'b11010011_00000111 : OUT <= 30;  //211 / 7 = 30
    16'b11010011_00001000 : OUT <= 26;  //211 / 8 = 26
    16'b11010011_00001001 : OUT <= 23;  //211 / 9 = 23
    16'b11010011_00001010 : OUT <= 21;  //211 / 10 = 21
    16'b11010011_00001011 : OUT <= 19;  //211 / 11 = 19
    16'b11010011_00001100 : OUT <= 17;  //211 / 12 = 17
    16'b11010011_00001101 : OUT <= 16;  //211 / 13 = 16
    16'b11010011_00001110 : OUT <= 15;  //211 / 14 = 15
    16'b11010011_00001111 : OUT <= 14;  //211 / 15 = 14
    16'b11010011_00010000 : OUT <= 13;  //211 / 16 = 13
    16'b11010011_00010001 : OUT <= 12;  //211 / 17 = 12
    16'b11010011_00010010 : OUT <= 11;  //211 / 18 = 11
    16'b11010011_00010011 : OUT <= 11;  //211 / 19 = 11
    16'b11010011_00010100 : OUT <= 10;  //211 / 20 = 10
    16'b11010011_00010101 : OUT <= 10;  //211 / 21 = 10
    16'b11010011_00010110 : OUT <= 9;  //211 / 22 = 9
    16'b11010011_00010111 : OUT <= 9;  //211 / 23 = 9
    16'b11010011_00011000 : OUT <= 8;  //211 / 24 = 8
    16'b11010011_00011001 : OUT <= 8;  //211 / 25 = 8
    16'b11010011_00011010 : OUT <= 8;  //211 / 26 = 8
    16'b11010011_00011011 : OUT <= 7;  //211 / 27 = 7
    16'b11010011_00011100 : OUT <= 7;  //211 / 28 = 7
    16'b11010011_00011101 : OUT <= 7;  //211 / 29 = 7
    16'b11010011_00011110 : OUT <= 7;  //211 / 30 = 7
    16'b11010011_00011111 : OUT <= 6;  //211 / 31 = 6
    16'b11010011_00100000 : OUT <= 6;  //211 / 32 = 6
    16'b11010011_00100001 : OUT <= 6;  //211 / 33 = 6
    16'b11010011_00100010 : OUT <= 6;  //211 / 34 = 6
    16'b11010011_00100011 : OUT <= 6;  //211 / 35 = 6
    16'b11010011_00100100 : OUT <= 5;  //211 / 36 = 5
    16'b11010011_00100101 : OUT <= 5;  //211 / 37 = 5
    16'b11010011_00100110 : OUT <= 5;  //211 / 38 = 5
    16'b11010011_00100111 : OUT <= 5;  //211 / 39 = 5
    16'b11010011_00101000 : OUT <= 5;  //211 / 40 = 5
    16'b11010011_00101001 : OUT <= 5;  //211 / 41 = 5
    16'b11010011_00101010 : OUT <= 5;  //211 / 42 = 5
    16'b11010011_00101011 : OUT <= 4;  //211 / 43 = 4
    16'b11010011_00101100 : OUT <= 4;  //211 / 44 = 4
    16'b11010011_00101101 : OUT <= 4;  //211 / 45 = 4
    16'b11010011_00101110 : OUT <= 4;  //211 / 46 = 4
    16'b11010011_00101111 : OUT <= 4;  //211 / 47 = 4
    16'b11010011_00110000 : OUT <= 4;  //211 / 48 = 4
    16'b11010011_00110001 : OUT <= 4;  //211 / 49 = 4
    16'b11010011_00110010 : OUT <= 4;  //211 / 50 = 4
    16'b11010011_00110011 : OUT <= 4;  //211 / 51 = 4
    16'b11010011_00110100 : OUT <= 4;  //211 / 52 = 4
    16'b11010011_00110101 : OUT <= 3;  //211 / 53 = 3
    16'b11010011_00110110 : OUT <= 3;  //211 / 54 = 3
    16'b11010011_00110111 : OUT <= 3;  //211 / 55 = 3
    16'b11010011_00111000 : OUT <= 3;  //211 / 56 = 3
    16'b11010011_00111001 : OUT <= 3;  //211 / 57 = 3
    16'b11010011_00111010 : OUT <= 3;  //211 / 58 = 3
    16'b11010011_00111011 : OUT <= 3;  //211 / 59 = 3
    16'b11010011_00111100 : OUT <= 3;  //211 / 60 = 3
    16'b11010011_00111101 : OUT <= 3;  //211 / 61 = 3
    16'b11010011_00111110 : OUT <= 3;  //211 / 62 = 3
    16'b11010011_00111111 : OUT <= 3;  //211 / 63 = 3
    16'b11010011_01000000 : OUT <= 3;  //211 / 64 = 3
    16'b11010011_01000001 : OUT <= 3;  //211 / 65 = 3
    16'b11010011_01000010 : OUT <= 3;  //211 / 66 = 3
    16'b11010011_01000011 : OUT <= 3;  //211 / 67 = 3
    16'b11010011_01000100 : OUT <= 3;  //211 / 68 = 3
    16'b11010011_01000101 : OUT <= 3;  //211 / 69 = 3
    16'b11010011_01000110 : OUT <= 3;  //211 / 70 = 3
    16'b11010011_01000111 : OUT <= 2;  //211 / 71 = 2
    16'b11010011_01001000 : OUT <= 2;  //211 / 72 = 2
    16'b11010011_01001001 : OUT <= 2;  //211 / 73 = 2
    16'b11010011_01001010 : OUT <= 2;  //211 / 74 = 2
    16'b11010011_01001011 : OUT <= 2;  //211 / 75 = 2
    16'b11010011_01001100 : OUT <= 2;  //211 / 76 = 2
    16'b11010011_01001101 : OUT <= 2;  //211 / 77 = 2
    16'b11010011_01001110 : OUT <= 2;  //211 / 78 = 2
    16'b11010011_01001111 : OUT <= 2;  //211 / 79 = 2
    16'b11010011_01010000 : OUT <= 2;  //211 / 80 = 2
    16'b11010011_01010001 : OUT <= 2;  //211 / 81 = 2
    16'b11010011_01010010 : OUT <= 2;  //211 / 82 = 2
    16'b11010011_01010011 : OUT <= 2;  //211 / 83 = 2
    16'b11010011_01010100 : OUT <= 2;  //211 / 84 = 2
    16'b11010011_01010101 : OUT <= 2;  //211 / 85 = 2
    16'b11010011_01010110 : OUT <= 2;  //211 / 86 = 2
    16'b11010011_01010111 : OUT <= 2;  //211 / 87 = 2
    16'b11010011_01011000 : OUT <= 2;  //211 / 88 = 2
    16'b11010011_01011001 : OUT <= 2;  //211 / 89 = 2
    16'b11010011_01011010 : OUT <= 2;  //211 / 90 = 2
    16'b11010011_01011011 : OUT <= 2;  //211 / 91 = 2
    16'b11010011_01011100 : OUT <= 2;  //211 / 92 = 2
    16'b11010011_01011101 : OUT <= 2;  //211 / 93 = 2
    16'b11010011_01011110 : OUT <= 2;  //211 / 94 = 2
    16'b11010011_01011111 : OUT <= 2;  //211 / 95 = 2
    16'b11010011_01100000 : OUT <= 2;  //211 / 96 = 2
    16'b11010011_01100001 : OUT <= 2;  //211 / 97 = 2
    16'b11010011_01100010 : OUT <= 2;  //211 / 98 = 2
    16'b11010011_01100011 : OUT <= 2;  //211 / 99 = 2
    16'b11010011_01100100 : OUT <= 2;  //211 / 100 = 2
    16'b11010011_01100101 : OUT <= 2;  //211 / 101 = 2
    16'b11010011_01100110 : OUT <= 2;  //211 / 102 = 2
    16'b11010011_01100111 : OUT <= 2;  //211 / 103 = 2
    16'b11010011_01101000 : OUT <= 2;  //211 / 104 = 2
    16'b11010011_01101001 : OUT <= 2;  //211 / 105 = 2
    16'b11010011_01101010 : OUT <= 1;  //211 / 106 = 1
    16'b11010011_01101011 : OUT <= 1;  //211 / 107 = 1
    16'b11010011_01101100 : OUT <= 1;  //211 / 108 = 1
    16'b11010011_01101101 : OUT <= 1;  //211 / 109 = 1
    16'b11010011_01101110 : OUT <= 1;  //211 / 110 = 1
    16'b11010011_01101111 : OUT <= 1;  //211 / 111 = 1
    16'b11010011_01110000 : OUT <= 1;  //211 / 112 = 1
    16'b11010011_01110001 : OUT <= 1;  //211 / 113 = 1
    16'b11010011_01110010 : OUT <= 1;  //211 / 114 = 1
    16'b11010011_01110011 : OUT <= 1;  //211 / 115 = 1
    16'b11010011_01110100 : OUT <= 1;  //211 / 116 = 1
    16'b11010011_01110101 : OUT <= 1;  //211 / 117 = 1
    16'b11010011_01110110 : OUT <= 1;  //211 / 118 = 1
    16'b11010011_01110111 : OUT <= 1;  //211 / 119 = 1
    16'b11010011_01111000 : OUT <= 1;  //211 / 120 = 1
    16'b11010011_01111001 : OUT <= 1;  //211 / 121 = 1
    16'b11010011_01111010 : OUT <= 1;  //211 / 122 = 1
    16'b11010011_01111011 : OUT <= 1;  //211 / 123 = 1
    16'b11010011_01111100 : OUT <= 1;  //211 / 124 = 1
    16'b11010011_01111101 : OUT <= 1;  //211 / 125 = 1
    16'b11010011_01111110 : OUT <= 1;  //211 / 126 = 1
    16'b11010011_01111111 : OUT <= 1;  //211 / 127 = 1
    16'b11010011_10000000 : OUT <= 1;  //211 / 128 = 1
    16'b11010011_10000001 : OUT <= 1;  //211 / 129 = 1
    16'b11010011_10000010 : OUT <= 1;  //211 / 130 = 1
    16'b11010011_10000011 : OUT <= 1;  //211 / 131 = 1
    16'b11010011_10000100 : OUT <= 1;  //211 / 132 = 1
    16'b11010011_10000101 : OUT <= 1;  //211 / 133 = 1
    16'b11010011_10000110 : OUT <= 1;  //211 / 134 = 1
    16'b11010011_10000111 : OUT <= 1;  //211 / 135 = 1
    16'b11010011_10001000 : OUT <= 1;  //211 / 136 = 1
    16'b11010011_10001001 : OUT <= 1;  //211 / 137 = 1
    16'b11010011_10001010 : OUT <= 1;  //211 / 138 = 1
    16'b11010011_10001011 : OUT <= 1;  //211 / 139 = 1
    16'b11010011_10001100 : OUT <= 1;  //211 / 140 = 1
    16'b11010011_10001101 : OUT <= 1;  //211 / 141 = 1
    16'b11010011_10001110 : OUT <= 1;  //211 / 142 = 1
    16'b11010011_10001111 : OUT <= 1;  //211 / 143 = 1
    16'b11010011_10010000 : OUT <= 1;  //211 / 144 = 1
    16'b11010011_10010001 : OUT <= 1;  //211 / 145 = 1
    16'b11010011_10010010 : OUT <= 1;  //211 / 146 = 1
    16'b11010011_10010011 : OUT <= 1;  //211 / 147 = 1
    16'b11010011_10010100 : OUT <= 1;  //211 / 148 = 1
    16'b11010011_10010101 : OUT <= 1;  //211 / 149 = 1
    16'b11010011_10010110 : OUT <= 1;  //211 / 150 = 1
    16'b11010011_10010111 : OUT <= 1;  //211 / 151 = 1
    16'b11010011_10011000 : OUT <= 1;  //211 / 152 = 1
    16'b11010011_10011001 : OUT <= 1;  //211 / 153 = 1
    16'b11010011_10011010 : OUT <= 1;  //211 / 154 = 1
    16'b11010011_10011011 : OUT <= 1;  //211 / 155 = 1
    16'b11010011_10011100 : OUT <= 1;  //211 / 156 = 1
    16'b11010011_10011101 : OUT <= 1;  //211 / 157 = 1
    16'b11010011_10011110 : OUT <= 1;  //211 / 158 = 1
    16'b11010011_10011111 : OUT <= 1;  //211 / 159 = 1
    16'b11010011_10100000 : OUT <= 1;  //211 / 160 = 1
    16'b11010011_10100001 : OUT <= 1;  //211 / 161 = 1
    16'b11010011_10100010 : OUT <= 1;  //211 / 162 = 1
    16'b11010011_10100011 : OUT <= 1;  //211 / 163 = 1
    16'b11010011_10100100 : OUT <= 1;  //211 / 164 = 1
    16'b11010011_10100101 : OUT <= 1;  //211 / 165 = 1
    16'b11010011_10100110 : OUT <= 1;  //211 / 166 = 1
    16'b11010011_10100111 : OUT <= 1;  //211 / 167 = 1
    16'b11010011_10101000 : OUT <= 1;  //211 / 168 = 1
    16'b11010011_10101001 : OUT <= 1;  //211 / 169 = 1
    16'b11010011_10101010 : OUT <= 1;  //211 / 170 = 1
    16'b11010011_10101011 : OUT <= 1;  //211 / 171 = 1
    16'b11010011_10101100 : OUT <= 1;  //211 / 172 = 1
    16'b11010011_10101101 : OUT <= 1;  //211 / 173 = 1
    16'b11010011_10101110 : OUT <= 1;  //211 / 174 = 1
    16'b11010011_10101111 : OUT <= 1;  //211 / 175 = 1
    16'b11010011_10110000 : OUT <= 1;  //211 / 176 = 1
    16'b11010011_10110001 : OUT <= 1;  //211 / 177 = 1
    16'b11010011_10110010 : OUT <= 1;  //211 / 178 = 1
    16'b11010011_10110011 : OUT <= 1;  //211 / 179 = 1
    16'b11010011_10110100 : OUT <= 1;  //211 / 180 = 1
    16'b11010011_10110101 : OUT <= 1;  //211 / 181 = 1
    16'b11010011_10110110 : OUT <= 1;  //211 / 182 = 1
    16'b11010011_10110111 : OUT <= 1;  //211 / 183 = 1
    16'b11010011_10111000 : OUT <= 1;  //211 / 184 = 1
    16'b11010011_10111001 : OUT <= 1;  //211 / 185 = 1
    16'b11010011_10111010 : OUT <= 1;  //211 / 186 = 1
    16'b11010011_10111011 : OUT <= 1;  //211 / 187 = 1
    16'b11010011_10111100 : OUT <= 1;  //211 / 188 = 1
    16'b11010011_10111101 : OUT <= 1;  //211 / 189 = 1
    16'b11010011_10111110 : OUT <= 1;  //211 / 190 = 1
    16'b11010011_10111111 : OUT <= 1;  //211 / 191 = 1
    16'b11010011_11000000 : OUT <= 1;  //211 / 192 = 1
    16'b11010011_11000001 : OUT <= 1;  //211 / 193 = 1
    16'b11010011_11000010 : OUT <= 1;  //211 / 194 = 1
    16'b11010011_11000011 : OUT <= 1;  //211 / 195 = 1
    16'b11010011_11000100 : OUT <= 1;  //211 / 196 = 1
    16'b11010011_11000101 : OUT <= 1;  //211 / 197 = 1
    16'b11010011_11000110 : OUT <= 1;  //211 / 198 = 1
    16'b11010011_11000111 : OUT <= 1;  //211 / 199 = 1
    16'b11010011_11001000 : OUT <= 1;  //211 / 200 = 1
    16'b11010011_11001001 : OUT <= 1;  //211 / 201 = 1
    16'b11010011_11001010 : OUT <= 1;  //211 / 202 = 1
    16'b11010011_11001011 : OUT <= 1;  //211 / 203 = 1
    16'b11010011_11001100 : OUT <= 1;  //211 / 204 = 1
    16'b11010011_11001101 : OUT <= 1;  //211 / 205 = 1
    16'b11010011_11001110 : OUT <= 1;  //211 / 206 = 1
    16'b11010011_11001111 : OUT <= 1;  //211 / 207 = 1
    16'b11010011_11010000 : OUT <= 1;  //211 / 208 = 1
    16'b11010011_11010001 : OUT <= 1;  //211 / 209 = 1
    16'b11010011_11010010 : OUT <= 1;  //211 / 210 = 1
    16'b11010011_11010011 : OUT <= 1;  //211 / 211 = 1
    16'b11010011_11010100 : OUT <= 0;  //211 / 212 = 0
    16'b11010011_11010101 : OUT <= 0;  //211 / 213 = 0
    16'b11010011_11010110 : OUT <= 0;  //211 / 214 = 0
    16'b11010011_11010111 : OUT <= 0;  //211 / 215 = 0
    16'b11010011_11011000 : OUT <= 0;  //211 / 216 = 0
    16'b11010011_11011001 : OUT <= 0;  //211 / 217 = 0
    16'b11010011_11011010 : OUT <= 0;  //211 / 218 = 0
    16'b11010011_11011011 : OUT <= 0;  //211 / 219 = 0
    16'b11010011_11011100 : OUT <= 0;  //211 / 220 = 0
    16'b11010011_11011101 : OUT <= 0;  //211 / 221 = 0
    16'b11010011_11011110 : OUT <= 0;  //211 / 222 = 0
    16'b11010011_11011111 : OUT <= 0;  //211 / 223 = 0
    16'b11010011_11100000 : OUT <= 0;  //211 / 224 = 0
    16'b11010011_11100001 : OUT <= 0;  //211 / 225 = 0
    16'b11010011_11100010 : OUT <= 0;  //211 / 226 = 0
    16'b11010011_11100011 : OUT <= 0;  //211 / 227 = 0
    16'b11010011_11100100 : OUT <= 0;  //211 / 228 = 0
    16'b11010011_11100101 : OUT <= 0;  //211 / 229 = 0
    16'b11010011_11100110 : OUT <= 0;  //211 / 230 = 0
    16'b11010011_11100111 : OUT <= 0;  //211 / 231 = 0
    16'b11010011_11101000 : OUT <= 0;  //211 / 232 = 0
    16'b11010011_11101001 : OUT <= 0;  //211 / 233 = 0
    16'b11010011_11101010 : OUT <= 0;  //211 / 234 = 0
    16'b11010011_11101011 : OUT <= 0;  //211 / 235 = 0
    16'b11010011_11101100 : OUT <= 0;  //211 / 236 = 0
    16'b11010011_11101101 : OUT <= 0;  //211 / 237 = 0
    16'b11010011_11101110 : OUT <= 0;  //211 / 238 = 0
    16'b11010011_11101111 : OUT <= 0;  //211 / 239 = 0
    16'b11010011_11110000 : OUT <= 0;  //211 / 240 = 0
    16'b11010011_11110001 : OUT <= 0;  //211 / 241 = 0
    16'b11010011_11110010 : OUT <= 0;  //211 / 242 = 0
    16'b11010011_11110011 : OUT <= 0;  //211 / 243 = 0
    16'b11010011_11110100 : OUT <= 0;  //211 / 244 = 0
    16'b11010011_11110101 : OUT <= 0;  //211 / 245 = 0
    16'b11010011_11110110 : OUT <= 0;  //211 / 246 = 0
    16'b11010011_11110111 : OUT <= 0;  //211 / 247 = 0
    16'b11010011_11111000 : OUT <= 0;  //211 / 248 = 0
    16'b11010011_11111001 : OUT <= 0;  //211 / 249 = 0
    16'b11010011_11111010 : OUT <= 0;  //211 / 250 = 0
    16'b11010011_11111011 : OUT <= 0;  //211 / 251 = 0
    16'b11010011_11111100 : OUT <= 0;  //211 / 252 = 0
    16'b11010011_11111101 : OUT <= 0;  //211 / 253 = 0
    16'b11010011_11111110 : OUT <= 0;  //211 / 254 = 0
    16'b11010011_11111111 : OUT <= 0;  //211 / 255 = 0
    16'b11010100_00000000 : OUT <= 0;  //212 / 0 = 0
    16'b11010100_00000001 : OUT <= 212;  //212 / 1 = 212
    16'b11010100_00000010 : OUT <= 106;  //212 / 2 = 106
    16'b11010100_00000011 : OUT <= 70;  //212 / 3 = 70
    16'b11010100_00000100 : OUT <= 53;  //212 / 4 = 53
    16'b11010100_00000101 : OUT <= 42;  //212 / 5 = 42
    16'b11010100_00000110 : OUT <= 35;  //212 / 6 = 35
    16'b11010100_00000111 : OUT <= 30;  //212 / 7 = 30
    16'b11010100_00001000 : OUT <= 26;  //212 / 8 = 26
    16'b11010100_00001001 : OUT <= 23;  //212 / 9 = 23
    16'b11010100_00001010 : OUT <= 21;  //212 / 10 = 21
    16'b11010100_00001011 : OUT <= 19;  //212 / 11 = 19
    16'b11010100_00001100 : OUT <= 17;  //212 / 12 = 17
    16'b11010100_00001101 : OUT <= 16;  //212 / 13 = 16
    16'b11010100_00001110 : OUT <= 15;  //212 / 14 = 15
    16'b11010100_00001111 : OUT <= 14;  //212 / 15 = 14
    16'b11010100_00010000 : OUT <= 13;  //212 / 16 = 13
    16'b11010100_00010001 : OUT <= 12;  //212 / 17 = 12
    16'b11010100_00010010 : OUT <= 11;  //212 / 18 = 11
    16'b11010100_00010011 : OUT <= 11;  //212 / 19 = 11
    16'b11010100_00010100 : OUT <= 10;  //212 / 20 = 10
    16'b11010100_00010101 : OUT <= 10;  //212 / 21 = 10
    16'b11010100_00010110 : OUT <= 9;  //212 / 22 = 9
    16'b11010100_00010111 : OUT <= 9;  //212 / 23 = 9
    16'b11010100_00011000 : OUT <= 8;  //212 / 24 = 8
    16'b11010100_00011001 : OUT <= 8;  //212 / 25 = 8
    16'b11010100_00011010 : OUT <= 8;  //212 / 26 = 8
    16'b11010100_00011011 : OUT <= 7;  //212 / 27 = 7
    16'b11010100_00011100 : OUT <= 7;  //212 / 28 = 7
    16'b11010100_00011101 : OUT <= 7;  //212 / 29 = 7
    16'b11010100_00011110 : OUT <= 7;  //212 / 30 = 7
    16'b11010100_00011111 : OUT <= 6;  //212 / 31 = 6
    16'b11010100_00100000 : OUT <= 6;  //212 / 32 = 6
    16'b11010100_00100001 : OUT <= 6;  //212 / 33 = 6
    16'b11010100_00100010 : OUT <= 6;  //212 / 34 = 6
    16'b11010100_00100011 : OUT <= 6;  //212 / 35 = 6
    16'b11010100_00100100 : OUT <= 5;  //212 / 36 = 5
    16'b11010100_00100101 : OUT <= 5;  //212 / 37 = 5
    16'b11010100_00100110 : OUT <= 5;  //212 / 38 = 5
    16'b11010100_00100111 : OUT <= 5;  //212 / 39 = 5
    16'b11010100_00101000 : OUT <= 5;  //212 / 40 = 5
    16'b11010100_00101001 : OUT <= 5;  //212 / 41 = 5
    16'b11010100_00101010 : OUT <= 5;  //212 / 42 = 5
    16'b11010100_00101011 : OUT <= 4;  //212 / 43 = 4
    16'b11010100_00101100 : OUT <= 4;  //212 / 44 = 4
    16'b11010100_00101101 : OUT <= 4;  //212 / 45 = 4
    16'b11010100_00101110 : OUT <= 4;  //212 / 46 = 4
    16'b11010100_00101111 : OUT <= 4;  //212 / 47 = 4
    16'b11010100_00110000 : OUT <= 4;  //212 / 48 = 4
    16'b11010100_00110001 : OUT <= 4;  //212 / 49 = 4
    16'b11010100_00110010 : OUT <= 4;  //212 / 50 = 4
    16'b11010100_00110011 : OUT <= 4;  //212 / 51 = 4
    16'b11010100_00110100 : OUT <= 4;  //212 / 52 = 4
    16'b11010100_00110101 : OUT <= 4;  //212 / 53 = 4
    16'b11010100_00110110 : OUT <= 3;  //212 / 54 = 3
    16'b11010100_00110111 : OUT <= 3;  //212 / 55 = 3
    16'b11010100_00111000 : OUT <= 3;  //212 / 56 = 3
    16'b11010100_00111001 : OUT <= 3;  //212 / 57 = 3
    16'b11010100_00111010 : OUT <= 3;  //212 / 58 = 3
    16'b11010100_00111011 : OUT <= 3;  //212 / 59 = 3
    16'b11010100_00111100 : OUT <= 3;  //212 / 60 = 3
    16'b11010100_00111101 : OUT <= 3;  //212 / 61 = 3
    16'b11010100_00111110 : OUT <= 3;  //212 / 62 = 3
    16'b11010100_00111111 : OUT <= 3;  //212 / 63 = 3
    16'b11010100_01000000 : OUT <= 3;  //212 / 64 = 3
    16'b11010100_01000001 : OUT <= 3;  //212 / 65 = 3
    16'b11010100_01000010 : OUT <= 3;  //212 / 66 = 3
    16'b11010100_01000011 : OUT <= 3;  //212 / 67 = 3
    16'b11010100_01000100 : OUT <= 3;  //212 / 68 = 3
    16'b11010100_01000101 : OUT <= 3;  //212 / 69 = 3
    16'b11010100_01000110 : OUT <= 3;  //212 / 70 = 3
    16'b11010100_01000111 : OUT <= 2;  //212 / 71 = 2
    16'b11010100_01001000 : OUT <= 2;  //212 / 72 = 2
    16'b11010100_01001001 : OUT <= 2;  //212 / 73 = 2
    16'b11010100_01001010 : OUT <= 2;  //212 / 74 = 2
    16'b11010100_01001011 : OUT <= 2;  //212 / 75 = 2
    16'b11010100_01001100 : OUT <= 2;  //212 / 76 = 2
    16'b11010100_01001101 : OUT <= 2;  //212 / 77 = 2
    16'b11010100_01001110 : OUT <= 2;  //212 / 78 = 2
    16'b11010100_01001111 : OUT <= 2;  //212 / 79 = 2
    16'b11010100_01010000 : OUT <= 2;  //212 / 80 = 2
    16'b11010100_01010001 : OUT <= 2;  //212 / 81 = 2
    16'b11010100_01010010 : OUT <= 2;  //212 / 82 = 2
    16'b11010100_01010011 : OUT <= 2;  //212 / 83 = 2
    16'b11010100_01010100 : OUT <= 2;  //212 / 84 = 2
    16'b11010100_01010101 : OUT <= 2;  //212 / 85 = 2
    16'b11010100_01010110 : OUT <= 2;  //212 / 86 = 2
    16'b11010100_01010111 : OUT <= 2;  //212 / 87 = 2
    16'b11010100_01011000 : OUT <= 2;  //212 / 88 = 2
    16'b11010100_01011001 : OUT <= 2;  //212 / 89 = 2
    16'b11010100_01011010 : OUT <= 2;  //212 / 90 = 2
    16'b11010100_01011011 : OUT <= 2;  //212 / 91 = 2
    16'b11010100_01011100 : OUT <= 2;  //212 / 92 = 2
    16'b11010100_01011101 : OUT <= 2;  //212 / 93 = 2
    16'b11010100_01011110 : OUT <= 2;  //212 / 94 = 2
    16'b11010100_01011111 : OUT <= 2;  //212 / 95 = 2
    16'b11010100_01100000 : OUT <= 2;  //212 / 96 = 2
    16'b11010100_01100001 : OUT <= 2;  //212 / 97 = 2
    16'b11010100_01100010 : OUT <= 2;  //212 / 98 = 2
    16'b11010100_01100011 : OUT <= 2;  //212 / 99 = 2
    16'b11010100_01100100 : OUT <= 2;  //212 / 100 = 2
    16'b11010100_01100101 : OUT <= 2;  //212 / 101 = 2
    16'b11010100_01100110 : OUT <= 2;  //212 / 102 = 2
    16'b11010100_01100111 : OUT <= 2;  //212 / 103 = 2
    16'b11010100_01101000 : OUT <= 2;  //212 / 104 = 2
    16'b11010100_01101001 : OUT <= 2;  //212 / 105 = 2
    16'b11010100_01101010 : OUT <= 2;  //212 / 106 = 2
    16'b11010100_01101011 : OUT <= 1;  //212 / 107 = 1
    16'b11010100_01101100 : OUT <= 1;  //212 / 108 = 1
    16'b11010100_01101101 : OUT <= 1;  //212 / 109 = 1
    16'b11010100_01101110 : OUT <= 1;  //212 / 110 = 1
    16'b11010100_01101111 : OUT <= 1;  //212 / 111 = 1
    16'b11010100_01110000 : OUT <= 1;  //212 / 112 = 1
    16'b11010100_01110001 : OUT <= 1;  //212 / 113 = 1
    16'b11010100_01110010 : OUT <= 1;  //212 / 114 = 1
    16'b11010100_01110011 : OUT <= 1;  //212 / 115 = 1
    16'b11010100_01110100 : OUT <= 1;  //212 / 116 = 1
    16'b11010100_01110101 : OUT <= 1;  //212 / 117 = 1
    16'b11010100_01110110 : OUT <= 1;  //212 / 118 = 1
    16'b11010100_01110111 : OUT <= 1;  //212 / 119 = 1
    16'b11010100_01111000 : OUT <= 1;  //212 / 120 = 1
    16'b11010100_01111001 : OUT <= 1;  //212 / 121 = 1
    16'b11010100_01111010 : OUT <= 1;  //212 / 122 = 1
    16'b11010100_01111011 : OUT <= 1;  //212 / 123 = 1
    16'b11010100_01111100 : OUT <= 1;  //212 / 124 = 1
    16'b11010100_01111101 : OUT <= 1;  //212 / 125 = 1
    16'b11010100_01111110 : OUT <= 1;  //212 / 126 = 1
    16'b11010100_01111111 : OUT <= 1;  //212 / 127 = 1
    16'b11010100_10000000 : OUT <= 1;  //212 / 128 = 1
    16'b11010100_10000001 : OUT <= 1;  //212 / 129 = 1
    16'b11010100_10000010 : OUT <= 1;  //212 / 130 = 1
    16'b11010100_10000011 : OUT <= 1;  //212 / 131 = 1
    16'b11010100_10000100 : OUT <= 1;  //212 / 132 = 1
    16'b11010100_10000101 : OUT <= 1;  //212 / 133 = 1
    16'b11010100_10000110 : OUT <= 1;  //212 / 134 = 1
    16'b11010100_10000111 : OUT <= 1;  //212 / 135 = 1
    16'b11010100_10001000 : OUT <= 1;  //212 / 136 = 1
    16'b11010100_10001001 : OUT <= 1;  //212 / 137 = 1
    16'b11010100_10001010 : OUT <= 1;  //212 / 138 = 1
    16'b11010100_10001011 : OUT <= 1;  //212 / 139 = 1
    16'b11010100_10001100 : OUT <= 1;  //212 / 140 = 1
    16'b11010100_10001101 : OUT <= 1;  //212 / 141 = 1
    16'b11010100_10001110 : OUT <= 1;  //212 / 142 = 1
    16'b11010100_10001111 : OUT <= 1;  //212 / 143 = 1
    16'b11010100_10010000 : OUT <= 1;  //212 / 144 = 1
    16'b11010100_10010001 : OUT <= 1;  //212 / 145 = 1
    16'b11010100_10010010 : OUT <= 1;  //212 / 146 = 1
    16'b11010100_10010011 : OUT <= 1;  //212 / 147 = 1
    16'b11010100_10010100 : OUT <= 1;  //212 / 148 = 1
    16'b11010100_10010101 : OUT <= 1;  //212 / 149 = 1
    16'b11010100_10010110 : OUT <= 1;  //212 / 150 = 1
    16'b11010100_10010111 : OUT <= 1;  //212 / 151 = 1
    16'b11010100_10011000 : OUT <= 1;  //212 / 152 = 1
    16'b11010100_10011001 : OUT <= 1;  //212 / 153 = 1
    16'b11010100_10011010 : OUT <= 1;  //212 / 154 = 1
    16'b11010100_10011011 : OUT <= 1;  //212 / 155 = 1
    16'b11010100_10011100 : OUT <= 1;  //212 / 156 = 1
    16'b11010100_10011101 : OUT <= 1;  //212 / 157 = 1
    16'b11010100_10011110 : OUT <= 1;  //212 / 158 = 1
    16'b11010100_10011111 : OUT <= 1;  //212 / 159 = 1
    16'b11010100_10100000 : OUT <= 1;  //212 / 160 = 1
    16'b11010100_10100001 : OUT <= 1;  //212 / 161 = 1
    16'b11010100_10100010 : OUT <= 1;  //212 / 162 = 1
    16'b11010100_10100011 : OUT <= 1;  //212 / 163 = 1
    16'b11010100_10100100 : OUT <= 1;  //212 / 164 = 1
    16'b11010100_10100101 : OUT <= 1;  //212 / 165 = 1
    16'b11010100_10100110 : OUT <= 1;  //212 / 166 = 1
    16'b11010100_10100111 : OUT <= 1;  //212 / 167 = 1
    16'b11010100_10101000 : OUT <= 1;  //212 / 168 = 1
    16'b11010100_10101001 : OUT <= 1;  //212 / 169 = 1
    16'b11010100_10101010 : OUT <= 1;  //212 / 170 = 1
    16'b11010100_10101011 : OUT <= 1;  //212 / 171 = 1
    16'b11010100_10101100 : OUT <= 1;  //212 / 172 = 1
    16'b11010100_10101101 : OUT <= 1;  //212 / 173 = 1
    16'b11010100_10101110 : OUT <= 1;  //212 / 174 = 1
    16'b11010100_10101111 : OUT <= 1;  //212 / 175 = 1
    16'b11010100_10110000 : OUT <= 1;  //212 / 176 = 1
    16'b11010100_10110001 : OUT <= 1;  //212 / 177 = 1
    16'b11010100_10110010 : OUT <= 1;  //212 / 178 = 1
    16'b11010100_10110011 : OUT <= 1;  //212 / 179 = 1
    16'b11010100_10110100 : OUT <= 1;  //212 / 180 = 1
    16'b11010100_10110101 : OUT <= 1;  //212 / 181 = 1
    16'b11010100_10110110 : OUT <= 1;  //212 / 182 = 1
    16'b11010100_10110111 : OUT <= 1;  //212 / 183 = 1
    16'b11010100_10111000 : OUT <= 1;  //212 / 184 = 1
    16'b11010100_10111001 : OUT <= 1;  //212 / 185 = 1
    16'b11010100_10111010 : OUT <= 1;  //212 / 186 = 1
    16'b11010100_10111011 : OUT <= 1;  //212 / 187 = 1
    16'b11010100_10111100 : OUT <= 1;  //212 / 188 = 1
    16'b11010100_10111101 : OUT <= 1;  //212 / 189 = 1
    16'b11010100_10111110 : OUT <= 1;  //212 / 190 = 1
    16'b11010100_10111111 : OUT <= 1;  //212 / 191 = 1
    16'b11010100_11000000 : OUT <= 1;  //212 / 192 = 1
    16'b11010100_11000001 : OUT <= 1;  //212 / 193 = 1
    16'b11010100_11000010 : OUT <= 1;  //212 / 194 = 1
    16'b11010100_11000011 : OUT <= 1;  //212 / 195 = 1
    16'b11010100_11000100 : OUT <= 1;  //212 / 196 = 1
    16'b11010100_11000101 : OUT <= 1;  //212 / 197 = 1
    16'b11010100_11000110 : OUT <= 1;  //212 / 198 = 1
    16'b11010100_11000111 : OUT <= 1;  //212 / 199 = 1
    16'b11010100_11001000 : OUT <= 1;  //212 / 200 = 1
    16'b11010100_11001001 : OUT <= 1;  //212 / 201 = 1
    16'b11010100_11001010 : OUT <= 1;  //212 / 202 = 1
    16'b11010100_11001011 : OUT <= 1;  //212 / 203 = 1
    16'b11010100_11001100 : OUT <= 1;  //212 / 204 = 1
    16'b11010100_11001101 : OUT <= 1;  //212 / 205 = 1
    16'b11010100_11001110 : OUT <= 1;  //212 / 206 = 1
    16'b11010100_11001111 : OUT <= 1;  //212 / 207 = 1
    16'b11010100_11010000 : OUT <= 1;  //212 / 208 = 1
    16'b11010100_11010001 : OUT <= 1;  //212 / 209 = 1
    16'b11010100_11010010 : OUT <= 1;  //212 / 210 = 1
    16'b11010100_11010011 : OUT <= 1;  //212 / 211 = 1
    16'b11010100_11010100 : OUT <= 1;  //212 / 212 = 1
    16'b11010100_11010101 : OUT <= 0;  //212 / 213 = 0
    16'b11010100_11010110 : OUT <= 0;  //212 / 214 = 0
    16'b11010100_11010111 : OUT <= 0;  //212 / 215 = 0
    16'b11010100_11011000 : OUT <= 0;  //212 / 216 = 0
    16'b11010100_11011001 : OUT <= 0;  //212 / 217 = 0
    16'b11010100_11011010 : OUT <= 0;  //212 / 218 = 0
    16'b11010100_11011011 : OUT <= 0;  //212 / 219 = 0
    16'b11010100_11011100 : OUT <= 0;  //212 / 220 = 0
    16'b11010100_11011101 : OUT <= 0;  //212 / 221 = 0
    16'b11010100_11011110 : OUT <= 0;  //212 / 222 = 0
    16'b11010100_11011111 : OUT <= 0;  //212 / 223 = 0
    16'b11010100_11100000 : OUT <= 0;  //212 / 224 = 0
    16'b11010100_11100001 : OUT <= 0;  //212 / 225 = 0
    16'b11010100_11100010 : OUT <= 0;  //212 / 226 = 0
    16'b11010100_11100011 : OUT <= 0;  //212 / 227 = 0
    16'b11010100_11100100 : OUT <= 0;  //212 / 228 = 0
    16'b11010100_11100101 : OUT <= 0;  //212 / 229 = 0
    16'b11010100_11100110 : OUT <= 0;  //212 / 230 = 0
    16'b11010100_11100111 : OUT <= 0;  //212 / 231 = 0
    16'b11010100_11101000 : OUT <= 0;  //212 / 232 = 0
    16'b11010100_11101001 : OUT <= 0;  //212 / 233 = 0
    16'b11010100_11101010 : OUT <= 0;  //212 / 234 = 0
    16'b11010100_11101011 : OUT <= 0;  //212 / 235 = 0
    16'b11010100_11101100 : OUT <= 0;  //212 / 236 = 0
    16'b11010100_11101101 : OUT <= 0;  //212 / 237 = 0
    16'b11010100_11101110 : OUT <= 0;  //212 / 238 = 0
    16'b11010100_11101111 : OUT <= 0;  //212 / 239 = 0
    16'b11010100_11110000 : OUT <= 0;  //212 / 240 = 0
    16'b11010100_11110001 : OUT <= 0;  //212 / 241 = 0
    16'b11010100_11110010 : OUT <= 0;  //212 / 242 = 0
    16'b11010100_11110011 : OUT <= 0;  //212 / 243 = 0
    16'b11010100_11110100 : OUT <= 0;  //212 / 244 = 0
    16'b11010100_11110101 : OUT <= 0;  //212 / 245 = 0
    16'b11010100_11110110 : OUT <= 0;  //212 / 246 = 0
    16'b11010100_11110111 : OUT <= 0;  //212 / 247 = 0
    16'b11010100_11111000 : OUT <= 0;  //212 / 248 = 0
    16'b11010100_11111001 : OUT <= 0;  //212 / 249 = 0
    16'b11010100_11111010 : OUT <= 0;  //212 / 250 = 0
    16'b11010100_11111011 : OUT <= 0;  //212 / 251 = 0
    16'b11010100_11111100 : OUT <= 0;  //212 / 252 = 0
    16'b11010100_11111101 : OUT <= 0;  //212 / 253 = 0
    16'b11010100_11111110 : OUT <= 0;  //212 / 254 = 0
    16'b11010100_11111111 : OUT <= 0;  //212 / 255 = 0
    16'b11010101_00000000 : OUT <= 0;  //213 / 0 = 0
    16'b11010101_00000001 : OUT <= 213;  //213 / 1 = 213
    16'b11010101_00000010 : OUT <= 106;  //213 / 2 = 106
    16'b11010101_00000011 : OUT <= 71;  //213 / 3 = 71
    16'b11010101_00000100 : OUT <= 53;  //213 / 4 = 53
    16'b11010101_00000101 : OUT <= 42;  //213 / 5 = 42
    16'b11010101_00000110 : OUT <= 35;  //213 / 6 = 35
    16'b11010101_00000111 : OUT <= 30;  //213 / 7 = 30
    16'b11010101_00001000 : OUT <= 26;  //213 / 8 = 26
    16'b11010101_00001001 : OUT <= 23;  //213 / 9 = 23
    16'b11010101_00001010 : OUT <= 21;  //213 / 10 = 21
    16'b11010101_00001011 : OUT <= 19;  //213 / 11 = 19
    16'b11010101_00001100 : OUT <= 17;  //213 / 12 = 17
    16'b11010101_00001101 : OUT <= 16;  //213 / 13 = 16
    16'b11010101_00001110 : OUT <= 15;  //213 / 14 = 15
    16'b11010101_00001111 : OUT <= 14;  //213 / 15 = 14
    16'b11010101_00010000 : OUT <= 13;  //213 / 16 = 13
    16'b11010101_00010001 : OUT <= 12;  //213 / 17 = 12
    16'b11010101_00010010 : OUT <= 11;  //213 / 18 = 11
    16'b11010101_00010011 : OUT <= 11;  //213 / 19 = 11
    16'b11010101_00010100 : OUT <= 10;  //213 / 20 = 10
    16'b11010101_00010101 : OUT <= 10;  //213 / 21 = 10
    16'b11010101_00010110 : OUT <= 9;  //213 / 22 = 9
    16'b11010101_00010111 : OUT <= 9;  //213 / 23 = 9
    16'b11010101_00011000 : OUT <= 8;  //213 / 24 = 8
    16'b11010101_00011001 : OUT <= 8;  //213 / 25 = 8
    16'b11010101_00011010 : OUT <= 8;  //213 / 26 = 8
    16'b11010101_00011011 : OUT <= 7;  //213 / 27 = 7
    16'b11010101_00011100 : OUT <= 7;  //213 / 28 = 7
    16'b11010101_00011101 : OUT <= 7;  //213 / 29 = 7
    16'b11010101_00011110 : OUT <= 7;  //213 / 30 = 7
    16'b11010101_00011111 : OUT <= 6;  //213 / 31 = 6
    16'b11010101_00100000 : OUT <= 6;  //213 / 32 = 6
    16'b11010101_00100001 : OUT <= 6;  //213 / 33 = 6
    16'b11010101_00100010 : OUT <= 6;  //213 / 34 = 6
    16'b11010101_00100011 : OUT <= 6;  //213 / 35 = 6
    16'b11010101_00100100 : OUT <= 5;  //213 / 36 = 5
    16'b11010101_00100101 : OUT <= 5;  //213 / 37 = 5
    16'b11010101_00100110 : OUT <= 5;  //213 / 38 = 5
    16'b11010101_00100111 : OUT <= 5;  //213 / 39 = 5
    16'b11010101_00101000 : OUT <= 5;  //213 / 40 = 5
    16'b11010101_00101001 : OUT <= 5;  //213 / 41 = 5
    16'b11010101_00101010 : OUT <= 5;  //213 / 42 = 5
    16'b11010101_00101011 : OUT <= 4;  //213 / 43 = 4
    16'b11010101_00101100 : OUT <= 4;  //213 / 44 = 4
    16'b11010101_00101101 : OUT <= 4;  //213 / 45 = 4
    16'b11010101_00101110 : OUT <= 4;  //213 / 46 = 4
    16'b11010101_00101111 : OUT <= 4;  //213 / 47 = 4
    16'b11010101_00110000 : OUT <= 4;  //213 / 48 = 4
    16'b11010101_00110001 : OUT <= 4;  //213 / 49 = 4
    16'b11010101_00110010 : OUT <= 4;  //213 / 50 = 4
    16'b11010101_00110011 : OUT <= 4;  //213 / 51 = 4
    16'b11010101_00110100 : OUT <= 4;  //213 / 52 = 4
    16'b11010101_00110101 : OUT <= 4;  //213 / 53 = 4
    16'b11010101_00110110 : OUT <= 3;  //213 / 54 = 3
    16'b11010101_00110111 : OUT <= 3;  //213 / 55 = 3
    16'b11010101_00111000 : OUT <= 3;  //213 / 56 = 3
    16'b11010101_00111001 : OUT <= 3;  //213 / 57 = 3
    16'b11010101_00111010 : OUT <= 3;  //213 / 58 = 3
    16'b11010101_00111011 : OUT <= 3;  //213 / 59 = 3
    16'b11010101_00111100 : OUT <= 3;  //213 / 60 = 3
    16'b11010101_00111101 : OUT <= 3;  //213 / 61 = 3
    16'b11010101_00111110 : OUT <= 3;  //213 / 62 = 3
    16'b11010101_00111111 : OUT <= 3;  //213 / 63 = 3
    16'b11010101_01000000 : OUT <= 3;  //213 / 64 = 3
    16'b11010101_01000001 : OUT <= 3;  //213 / 65 = 3
    16'b11010101_01000010 : OUT <= 3;  //213 / 66 = 3
    16'b11010101_01000011 : OUT <= 3;  //213 / 67 = 3
    16'b11010101_01000100 : OUT <= 3;  //213 / 68 = 3
    16'b11010101_01000101 : OUT <= 3;  //213 / 69 = 3
    16'b11010101_01000110 : OUT <= 3;  //213 / 70 = 3
    16'b11010101_01000111 : OUT <= 3;  //213 / 71 = 3
    16'b11010101_01001000 : OUT <= 2;  //213 / 72 = 2
    16'b11010101_01001001 : OUT <= 2;  //213 / 73 = 2
    16'b11010101_01001010 : OUT <= 2;  //213 / 74 = 2
    16'b11010101_01001011 : OUT <= 2;  //213 / 75 = 2
    16'b11010101_01001100 : OUT <= 2;  //213 / 76 = 2
    16'b11010101_01001101 : OUT <= 2;  //213 / 77 = 2
    16'b11010101_01001110 : OUT <= 2;  //213 / 78 = 2
    16'b11010101_01001111 : OUT <= 2;  //213 / 79 = 2
    16'b11010101_01010000 : OUT <= 2;  //213 / 80 = 2
    16'b11010101_01010001 : OUT <= 2;  //213 / 81 = 2
    16'b11010101_01010010 : OUT <= 2;  //213 / 82 = 2
    16'b11010101_01010011 : OUT <= 2;  //213 / 83 = 2
    16'b11010101_01010100 : OUT <= 2;  //213 / 84 = 2
    16'b11010101_01010101 : OUT <= 2;  //213 / 85 = 2
    16'b11010101_01010110 : OUT <= 2;  //213 / 86 = 2
    16'b11010101_01010111 : OUT <= 2;  //213 / 87 = 2
    16'b11010101_01011000 : OUT <= 2;  //213 / 88 = 2
    16'b11010101_01011001 : OUT <= 2;  //213 / 89 = 2
    16'b11010101_01011010 : OUT <= 2;  //213 / 90 = 2
    16'b11010101_01011011 : OUT <= 2;  //213 / 91 = 2
    16'b11010101_01011100 : OUT <= 2;  //213 / 92 = 2
    16'b11010101_01011101 : OUT <= 2;  //213 / 93 = 2
    16'b11010101_01011110 : OUT <= 2;  //213 / 94 = 2
    16'b11010101_01011111 : OUT <= 2;  //213 / 95 = 2
    16'b11010101_01100000 : OUT <= 2;  //213 / 96 = 2
    16'b11010101_01100001 : OUT <= 2;  //213 / 97 = 2
    16'b11010101_01100010 : OUT <= 2;  //213 / 98 = 2
    16'b11010101_01100011 : OUT <= 2;  //213 / 99 = 2
    16'b11010101_01100100 : OUT <= 2;  //213 / 100 = 2
    16'b11010101_01100101 : OUT <= 2;  //213 / 101 = 2
    16'b11010101_01100110 : OUT <= 2;  //213 / 102 = 2
    16'b11010101_01100111 : OUT <= 2;  //213 / 103 = 2
    16'b11010101_01101000 : OUT <= 2;  //213 / 104 = 2
    16'b11010101_01101001 : OUT <= 2;  //213 / 105 = 2
    16'b11010101_01101010 : OUT <= 2;  //213 / 106 = 2
    16'b11010101_01101011 : OUT <= 1;  //213 / 107 = 1
    16'b11010101_01101100 : OUT <= 1;  //213 / 108 = 1
    16'b11010101_01101101 : OUT <= 1;  //213 / 109 = 1
    16'b11010101_01101110 : OUT <= 1;  //213 / 110 = 1
    16'b11010101_01101111 : OUT <= 1;  //213 / 111 = 1
    16'b11010101_01110000 : OUT <= 1;  //213 / 112 = 1
    16'b11010101_01110001 : OUT <= 1;  //213 / 113 = 1
    16'b11010101_01110010 : OUT <= 1;  //213 / 114 = 1
    16'b11010101_01110011 : OUT <= 1;  //213 / 115 = 1
    16'b11010101_01110100 : OUT <= 1;  //213 / 116 = 1
    16'b11010101_01110101 : OUT <= 1;  //213 / 117 = 1
    16'b11010101_01110110 : OUT <= 1;  //213 / 118 = 1
    16'b11010101_01110111 : OUT <= 1;  //213 / 119 = 1
    16'b11010101_01111000 : OUT <= 1;  //213 / 120 = 1
    16'b11010101_01111001 : OUT <= 1;  //213 / 121 = 1
    16'b11010101_01111010 : OUT <= 1;  //213 / 122 = 1
    16'b11010101_01111011 : OUT <= 1;  //213 / 123 = 1
    16'b11010101_01111100 : OUT <= 1;  //213 / 124 = 1
    16'b11010101_01111101 : OUT <= 1;  //213 / 125 = 1
    16'b11010101_01111110 : OUT <= 1;  //213 / 126 = 1
    16'b11010101_01111111 : OUT <= 1;  //213 / 127 = 1
    16'b11010101_10000000 : OUT <= 1;  //213 / 128 = 1
    16'b11010101_10000001 : OUT <= 1;  //213 / 129 = 1
    16'b11010101_10000010 : OUT <= 1;  //213 / 130 = 1
    16'b11010101_10000011 : OUT <= 1;  //213 / 131 = 1
    16'b11010101_10000100 : OUT <= 1;  //213 / 132 = 1
    16'b11010101_10000101 : OUT <= 1;  //213 / 133 = 1
    16'b11010101_10000110 : OUT <= 1;  //213 / 134 = 1
    16'b11010101_10000111 : OUT <= 1;  //213 / 135 = 1
    16'b11010101_10001000 : OUT <= 1;  //213 / 136 = 1
    16'b11010101_10001001 : OUT <= 1;  //213 / 137 = 1
    16'b11010101_10001010 : OUT <= 1;  //213 / 138 = 1
    16'b11010101_10001011 : OUT <= 1;  //213 / 139 = 1
    16'b11010101_10001100 : OUT <= 1;  //213 / 140 = 1
    16'b11010101_10001101 : OUT <= 1;  //213 / 141 = 1
    16'b11010101_10001110 : OUT <= 1;  //213 / 142 = 1
    16'b11010101_10001111 : OUT <= 1;  //213 / 143 = 1
    16'b11010101_10010000 : OUT <= 1;  //213 / 144 = 1
    16'b11010101_10010001 : OUT <= 1;  //213 / 145 = 1
    16'b11010101_10010010 : OUT <= 1;  //213 / 146 = 1
    16'b11010101_10010011 : OUT <= 1;  //213 / 147 = 1
    16'b11010101_10010100 : OUT <= 1;  //213 / 148 = 1
    16'b11010101_10010101 : OUT <= 1;  //213 / 149 = 1
    16'b11010101_10010110 : OUT <= 1;  //213 / 150 = 1
    16'b11010101_10010111 : OUT <= 1;  //213 / 151 = 1
    16'b11010101_10011000 : OUT <= 1;  //213 / 152 = 1
    16'b11010101_10011001 : OUT <= 1;  //213 / 153 = 1
    16'b11010101_10011010 : OUT <= 1;  //213 / 154 = 1
    16'b11010101_10011011 : OUT <= 1;  //213 / 155 = 1
    16'b11010101_10011100 : OUT <= 1;  //213 / 156 = 1
    16'b11010101_10011101 : OUT <= 1;  //213 / 157 = 1
    16'b11010101_10011110 : OUT <= 1;  //213 / 158 = 1
    16'b11010101_10011111 : OUT <= 1;  //213 / 159 = 1
    16'b11010101_10100000 : OUT <= 1;  //213 / 160 = 1
    16'b11010101_10100001 : OUT <= 1;  //213 / 161 = 1
    16'b11010101_10100010 : OUT <= 1;  //213 / 162 = 1
    16'b11010101_10100011 : OUT <= 1;  //213 / 163 = 1
    16'b11010101_10100100 : OUT <= 1;  //213 / 164 = 1
    16'b11010101_10100101 : OUT <= 1;  //213 / 165 = 1
    16'b11010101_10100110 : OUT <= 1;  //213 / 166 = 1
    16'b11010101_10100111 : OUT <= 1;  //213 / 167 = 1
    16'b11010101_10101000 : OUT <= 1;  //213 / 168 = 1
    16'b11010101_10101001 : OUT <= 1;  //213 / 169 = 1
    16'b11010101_10101010 : OUT <= 1;  //213 / 170 = 1
    16'b11010101_10101011 : OUT <= 1;  //213 / 171 = 1
    16'b11010101_10101100 : OUT <= 1;  //213 / 172 = 1
    16'b11010101_10101101 : OUT <= 1;  //213 / 173 = 1
    16'b11010101_10101110 : OUT <= 1;  //213 / 174 = 1
    16'b11010101_10101111 : OUT <= 1;  //213 / 175 = 1
    16'b11010101_10110000 : OUT <= 1;  //213 / 176 = 1
    16'b11010101_10110001 : OUT <= 1;  //213 / 177 = 1
    16'b11010101_10110010 : OUT <= 1;  //213 / 178 = 1
    16'b11010101_10110011 : OUT <= 1;  //213 / 179 = 1
    16'b11010101_10110100 : OUT <= 1;  //213 / 180 = 1
    16'b11010101_10110101 : OUT <= 1;  //213 / 181 = 1
    16'b11010101_10110110 : OUT <= 1;  //213 / 182 = 1
    16'b11010101_10110111 : OUT <= 1;  //213 / 183 = 1
    16'b11010101_10111000 : OUT <= 1;  //213 / 184 = 1
    16'b11010101_10111001 : OUT <= 1;  //213 / 185 = 1
    16'b11010101_10111010 : OUT <= 1;  //213 / 186 = 1
    16'b11010101_10111011 : OUT <= 1;  //213 / 187 = 1
    16'b11010101_10111100 : OUT <= 1;  //213 / 188 = 1
    16'b11010101_10111101 : OUT <= 1;  //213 / 189 = 1
    16'b11010101_10111110 : OUT <= 1;  //213 / 190 = 1
    16'b11010101_10111111 : OUT <= 1;  //213 / 191 = 1
    16'b11010101_11000000 : OUT <= 1;  //213 / 192 = 1
    16'b11010101_11000001 : OUT <= 1;  //213 / 193 = 1
    16'b11010101_11000010 : OUT <= 1;  //213 / 194 = 1
    16'b11010101_11000011 : OUT <= 1;  //213 / 195 = 1
    16'b11010101_11000100 : OUT <= 1;  //213 / 196 = 1
    16'b11010101_11000101 : OUT <= 1;  //213 / 197 = 1
    16'b11010101_11000110 : OUT <= 1;  //213 / 198 = 1
    16'b11010101_11000111 : OUT <= 1;  //213 / 199 = 1
    16'b11010101_11001000 : OUT <= 1;  //213 / 200 = 1
    16'b11010101_11001001 : OUT <= 1;  //213 / 201 = 1
    16'b11010101_11001010 : OUT <= 1;  //213 / 202 = 1
    16'b11010101_11001011 : OUT <= 1;  //213 / 203 = 1
    16'b11010101_11001100 : OUT <= 1;  //213 / 204 = 1
    16'b11010101_11001101 : OUT <= 1;  //213 / 205 = 1
    16'b11010101_11001110 : OUT <= 1;  //213 / 206 = 1
    16'b11010101_11001111 : OUT <= 1;  //213 / 207 = 1
    16'b11010101_11010000 : OUT <= 1;  //213 / 208 = 1
    16'b11010101_11010001 : OUT <= 1;  //213 / 209 = 1
    16'b11010101_11010010 : OUT <= 1;  //213 / 210 = 1
    16'b11010101_11010011 : OUT <= 1;  //213 / 211 = 1
    16'b11010101_11010100 : OUT <= 1;  //213 / 212 = 1
    16'b11010101_11010101 : OUT <= 1;  //213 / 213 = 1
    16'b11010101_11010110 : OUT <= 0;  //213 / 214 = 0
    16'b11010101_11010111 : OUT <= 0;  //213 / 215 = 0
    16'b11010101_11011000 : OUT <= 0;  //213 / 216 = 0
    16'b11010101_11011001 : OUT <= 0;  //213 / 217 = 0
    16'b11010101_11011010 : OUT <= 0;  //213 / 218 = 0
    16'b11010101_11011011 : OUT <= 0;  //213 / 219 = 0
    16'b11010101_11011100 : OUT <= 0;  //213 / 220 = 0
    16'b11010101_11011101 : OUT <= 0;  //213 / 221 = 0
    16'b11010101_11011110 : OUT <= 0;  //213 / 222 = 0
    16'b11010101_11011111 : OUT <= 0;  //213 / 223 = 0
    16'b11010101_11100000 : OUT <= 0;  //213 / 224 = 0
    16'b11010101_11100001 : OUT <= 0;  //213 / 225 = 0
    16'b11010101_11100010 : OUT <= 0;  //213 / 226 = 0
    16'b11010101_11100011 : OUT <= 0;  //213 / 227 = 0
    16'b11010101_11100100 : OUT <= 0;  //213 / 228 = 0
    16'b11010101_11100101 : OUT <= 0;  //213 / 229 = 0
    16'b11010101_11100110 : OUT <= 0;  //213 / 230 = 0
    16'b11010101_11100111 : OUT <= 0;  //213 / 231 = 0
    16'b11010101_11101000 : OUT <= 0;  //213 / 232 = 0
    16'b11010101_11101001 : OUT <= 0;  //213 / 233 = 0
    16'b11010101_11101010 : OUT <= 0;  //213 / 234 = 0
    16'b11010101_11101011 : OUT <= 0;  //213 / 235 = 0
    16'b11010101_11101100 : OUT <= 0;  //213 / 236 = 0
    16'b11010101_11101101 : OUT <= 0;  //213 / 237 = 0
    16'b11010101_11101110 : OUT <= 0;  //213 / 238 = 0
    16'b11010101_11101111 : OUT <= 0;  //213 / 239 = 0
    16'b11010101_11110000 : OUT <= 0;  //213 / 240 = 0
    16'b11010101_11110001 : OUT <= 0;  //213 / 241 = 0
    16'b11010101_11110010 : OUT <= 0;  //213 / 242 = 0
    16'b11010101_11110011 : OUT <= 0;  //213 / 243 = 0
    16'b11010101_11110100 : OUT <= 0;  //213 / 244 = 0
    16'b11010101_11110101 : OUT <= 0;  //213 / 245 = 0
    16'b11010101_11110110 : OUT <= 0;  //213 / 246 = 0
    16'b11010101_11110111 : OUT <= 0;  //213 / 247 = 0
    16'b11010101_11111000 : OUT <= 0;  //213 / 248 = 0
    16'b11010101_11111001 : OUT <= 0;  //213 / 249 = 0
    16'b11010101_11111010 : OUT <= 0;  //213 / 250 = 0
    16'b11010101_11111011 : OUT <= 0;  //213 / 251 = 0
    16'b11010101_11111100 : OUT <= 0;  //213 / 252 = 0
    16'b11010101_11111101 : OUT <= 0;  //213 / 253 = 0
    16'b11010101_11111110 : OUT <= 0;  //213 / 254 = 0
    16'b11010101_11111111 : OUT <= 0;  //213 / 255 = 0
    16'b11010110_00000000 : OUT <= 0;  //214 / 0 = 0
    16'b11010110_00000001 : OUT <= 214;  //214 / 1 = 214
    16'b11010110_00000010 : OUT <= 107;  //214 / 2 = 107
    16'b11010110_00000011 : OUT <= 71;  //214 / 3 = 71
    16'b11010110_00000100 : OUT <= 53;  //214 / 4 = 53
    16'b11010110_00000101 : OUT <= 42;  //214 / 5 = 42
    16'b11010110_00000110 : OUT <= 35;  //214 / 6 = 35
    16'b11010110_00000111 : OUT <= 30;  //214 / 7 = 30
    16'b11010110_00001000 : OUT <= 26;  //214 / 8 = 26
    16'b11010110_00001001 : OUT <= 23;  //214 / 9 = 23
    16'b11010110_00001010 : OUT <= 21;  //214 / 10 = 21
    16'b11010110_00001011 : OUT <= 19;  //214 / 11 = 19
    16'b11010110_00001100 : OUT <= 17;  //214 / 12 = 17
    16'b11010110_00001101 : OUT <= 16;  //214 / 13 = 16
    16'b11010110_00001110 : OUT <= 15;  //214 / 14 = 15
    16'b11010110_00001111 : OUT <= 14;  //214 / 15 = 14
    16'b11010110_00010000 : OUT <= 13;  //214 / 16 = 13
    16'b11010110_00010001 : OUT <= 12;  //214 / 17 = 12
    16'b11010110_00010010 : OUT <= 11;  //214 / 18 = 11
    16'b11010110_00010011 : OUT <= 11;  //214 / 19 = 11
    16'b11010110_00010100 : OUT <= 10;  //214 / 20 = 10
    16'b11010110_00010101 : OUT <= 10;  //214 / 21 = 10
    16'b11010110_00010110 : OUT <= 9;  //214 / 22 = 9
    16'b11010110_00010111 : OUT <= 9;  //214 / 23 = 9
    16'b11010110_00011000 : OUT <= 8;  //214 / 24 = 8
    16'b11010110_00011001 : OUT <= 8;  //214 / 25 = 8
    16'b11010110_00011010 : OUT <= 8;  //214 / 26 = 8
    16'b11010110_00011011 : OUT <= 7;  //214 / 27 = 7
    16'b11010110_00011100 : OUT <= 7;  //214 / 28 = 7
    16'b11010110_00011101 : OUT <= 7;  //214 / 29 = 7
    16'b11010110_00011110 : OUT <= 7;  //214 / 30 = 7
    16'b11010110_00011111 : OUT <= 6;  //214 / 31 = 6
    16'b11010110_00100000 : OUT <= 6;  //214 / 32 = 6
    16'b11010110_00100001 : OUT <= 6;  //214 / 33 = 6
    16'b11010110_00100010 : OUT <= 6;  //214 / 34 = 6
    16'b11010110_00100011 : OUT <= 6;  //214 / 35 = 6
    16'b11010110_00100100 : OUT <= 5;  //214 / 36 = 5
    16'b11010110_00100101 : OUT <= 5;  //214 / 37 = 5
    16'b11010110_00100110 : OUT <= 5;  //214 / 38 = 5
    16'b11010110_00100111 : OUT <= 5;  //214 / 39 = 5
    16'b11010110_00101000 : OUT <= 5;  //214 / 40 = 5
    16'b11010110_00101001 : OUT <= 5;  //214 / 41 = 5
    16'b11010110_00101010 : OUT <= 5;  //214 / 42 = 5
    16'b11010110_00101011 : OUT <= 4;  //214 / 43 = 4
    16'b11010110_00101100 : OUT <= 4;  //214 / 44 = 4
    16'b11010110_00101101 : OUT <= 4;  //214 / 45 = 4
    16'b11010110_00101110 : OUT <= 4;  //214 / 46 = 4
    16'b11010110_00101111 : OUT <= 4;  //214 / 47 = 4
    16'b11010110_00110000 : OUT <= 4;  //214 / 48 = 4
    16'b11010110_00110001 : OUT <= 4;  //214 / 49 = 4
    16'b11010110_00110010 : OUT <= 4;  //214 / 50 = 4
    16'b11010110_00110011 : OUT <= 4;  //214 / 51 = 4
    16'b11010110_00110100 : OUT <= 4;  //214 / 52 = 4
    16'b11010110_00110101 : OUT <= 4;  //214 / 53 = 4
    16'b11010110_00110110 : OUT <= 3;  //214 / 54 = 3
    16'b11010110_00110111 : OUT <= 3;  //214 / 55 = 3
    16'b11010110_00111000 : OUT <= 3;  //214 / 56 = 3
    16'b11010110_00111001 : OUT <= 3;  //214 / 57 = 3
    16'b11010110_00111010 : OUT <= 3;  //214 / 58 = 3
    16'b11010110_00111011 : OUT <= 3;  //214 / 59 = 3
    16'b11010110_00111100 : OUT <= 3;  //214 / 60 = 3
    16'b11010110_00111101 : OUT <= 3;  //214 / 61 = 3
    16'b11010110_00111110 : OUT <= 3;  //214 / 62 = 3
    16'b11010110_00111111 : OUT <= 3;  //214 / 63 = 3
    16'b11010110_01000000 : OUT <= 3;  //214 / 64 = 3
    16'b11010110_01000001 : OUT <= 3;  //214 / 65 = 3
    16'b11010110_01000010 : OUT <= 3;  //214 / 66 = 3
    16'b11010110_01000011 : OUT <= 3;  //214 / 67 = 3
    16'b11010110_01000100 : OUT <= 3;  //214 / 68 = 3
    16'b11010110_01000101 : OUT <= 3;  //214 / 69 = 3
    16'b11010110_01000110 : OUT <= 3;  //214 / 70 = 3
    16'b11010110_01000111 : OUT <= 3;  //214 / 71 = 3
    16'b11010110_01001000 : OUT <= 2;  //214 / 72 = 2
    16'b11010110_01001001 : OUT <= 2;  //214 / 73 = 2
    16'b11010110_01001010 : OUT <= 2;  //214 / 74 = 2
    16'b11010110_01001011 : OUT <= 2;  //214 / 75 = 2
    16'b11010110_01001100 : OUT <= 2;  //214 / 76 = 2
    16'b11010110_01001101 : OUT <= 2;  //214 / 77 = 2
    16'b11010110_01001110 : OUT <= 2;  //214 / 78 = 2
    16'b11010110_01001111 : OUT <= 2;  //214 / 79 = 2
    16'b11010110_01010000 : OUT <= 2;  //214 / 80 = 2
    16'b11010110_01010001 : OUT <= 2;  //214 / 81 = 2
    16'b11010110_01010010 : OUT <= 2;  //214 / 82 = 2
    16'b11010110_01010011 : OUT <= 2;  //214 / 83 = 2
    16'b11010110_01010100 : OUT <= 2;  //214 / 84 = 2
    16'b11010110_01010101 : OUT <= 2;  //214 / 85 = 2
    16'b11010110_01010110 : OUT <= 2;  //214 / 86 = 2
    16'b11010110_01010111 : OUT <= 2;  //214 / 87 = 2
    16'b11010110_01011000 : OUT <= 2;  //214 / 88 = 2
    16'b11010110_01011001 : OUT <= 2;  //214 / 89 = 2
    16'b11010110_01011010 : OUT <= 2;  //214 / 90 = 2
    16'b11010110_01011011 : OUT <= 2;  //214 / 91 = 2
    16'b11010110_01011100 : OUT <= 2;  //214 / 92 = 2
    16'b11010110_01011101 : OUT <= 2;  //214 / 93 = 2
    16'b11010110_01011110 : OUT <= 2;  //214 / 94 = 2
    16'b11010110_01011111 : OUT <= 2;  //214 / 95 = 2
    16'b11010110_01100000 : OUT <= 2;  //214 / 96 = 2
    16'b11010110_01100001 : OUT <= 2;  //214 / 97 = 2
    16'b11010110_01100010 : OUT <= 2;  //214 / 98 = 2
    16'b11010110_01100011 : OUT <= 2;  //214 / 99 = 2
    16'b11010110_01100100 : OUT <= 2;  //214 / 100 = 2
    16'b11010110_01100101 : OUT <= 2;  //214 / 101 = 2
    16'b11010110_01100110 : OUT <= 2;  //214 / 102 = 2
    16'b11010110_01100111 : OUT <= 2;  //214 / 103 = 2
    16'b11010110_01101000 : OUT <= 2;  //214 / 104 = 2
    16'b11010110_01101001 : OUT <= 2;  //214 / 105 = 2
    16'b11010110_01101010 : OUT <= 2;  //214 / 106 = 2
    16'b11010110_01101011 : OUT <= 2;  //214 / 107 = 2
    16'b11010110_01101100 : OUT <= 1;  //214 / 108 = 1
    16'b11010110_01101101 : OUT <= 1;  //214 / 109 = 1
    16'b11010110_01101110 : OUT <= 1;  //214 / 110 = 1
    16'b11010110_01101111 : OUT <= 1;  //214 / 111 = 1
    16'b11010110_01110000 : OUT <= 1;  //214 / 112 = 1
    16'b11010110_01110001 : OUT <= 1;  //214 / 113 = 1
    16'b11010110_01110010 : OUT <= 1;  //214 / 114 = 1
    16'b11010110_01110011 : OUT <= 1;  //214 / 115 = 1
    16'b11010110_01110100 : OUT <= 1;  //214 / 116 = 1
    16'b11010110_01110101 : OUT <= 1;  //214 / 117 = 1
    16'b11010110_01110110 : OUT <= 1;  //214 / 118 = 1
    16'b11010110_01110111 : OUT <= 1;  //214 / 119 = 1
    16'b11010110_01111000 : OUT <= 1;  //214 / 120 = 1
    16'b11010110_01111001 : OUT <= 1;  //214 / 121 = 1
    16'b11010110_01111010 : OUT <= 1;  //214 / 122 = 1
    16'b11010110_01111011 : OUT <= 1;  //214 / 123 = 1
    16'b11010110_01111100 : OUT <= 1;  //214 / 124 = 1
    16'b11010110_01111101 : OUT <= 1;  //214 / 125 = 1
    16'b11010110_01111110 : OUT <= 1;  //214 / 126 = 1
    16'b11010110_01111111 : OUT <= 1;  //214 / 127 = 1
    16'b11010110_10000000 : OUT <= 1;  //214 / 128 = 1
    16'b11010110_10000001 : OUT <= 1;  //214 / 129 = 1
    16'b11010110_10000010 : OUT <= 1;  //214 / 130 = 1
    16'b11010110_10000011 : OUT <= 1;  //214 / 131 = 1
    16'b11010110_10000100 : OUT <= 1;  //214 / 132 = 1
    16'b11010110_10000101 : OUT <= 1;  //214 / 133 = 1
    16'b11010110_10000110 : OUT <= 1;  //214 / 134 = 1
    16'b11010110_10000111 : OUT <= 1;  //214 / 135 = 1
    16'b11010110_10001000 : OUT <= 1;  //214 / 136 = 1
    16'b11010110_10001001 : OUT <= 1;  //214 / 137 = 1
    16'b11010110_10001010 : OUT <= 1;  //214 / 138 = 1
    16'b11010110_10001011 : OUT <= 1;  //214 / 139 = 1
    16'b11010110_10001100 : OUT <= 1;  //214 / 140 = 1
    16'b11010110_10001101 : OUT <= 1;  //214 / 141 = 1
    16'b11010110_10001110 : OUT <= 1;  //214 / 142 = 1
    16'b11010110_10001111 : OUT <= 1;  //214 / 143 = 1
    16'b11010110_10010000 : OUT <= 1;  //214 / 144 = 1
    16'b11010110_10010001 : OUT <= 1;  //214 / 145 = 1
    16'b11010110_10010010 : OUT <= 1;  //214 / 146 = 1
    16'b11010110_10010011 : OUT <= 1;  //214 / 147 = 1
    16'b11010110_10010100 : OUT <= 1;  //214 / 148 = 1
    16'b11010110_10010101 : OUT <= 1;  //214 / 149 = 1
    16'b11010110_10010110 : OUT <= 1;  //214 / 150 = 1
    16'b11010110_10010111 : OUT <= 1;  //214 / 151 = 1
    16'b11010110_10011000 : OUT <= 1;  //214 / 152 = 1
    16'b11010110_10011001 : OUT <= 1;  //214 / 153 = 1
    16'b11010110_10011010 : OUT <= 1;  //214 / 154 = 1
    16'b11010110_10011011 : OUT <= 1;  //214 / 155 = 1
    16'b11010110_10011100 : OUT <= 1;  //214 / 156 = 1
    16'b11010110_10011101 : OUT <= 1;  //214 / 157 = 1
    16'b11010110_10011110 : OUT <= 1;  //214 / 158 = 1
    16'b11010110_10011111 : OUT <= 1;  //214 / 159 = 1
    16'b11010110_10100000 : OUT <= 1;  //214 / 160 = 1
    16'b11010110_10100001 : OUT <= 1;  //214 / 161 = 1
    16'b11010110_10100010 : OUT <= 1;  //214 / 162 = 1
    16'b11010110_10100011 : OUT <= 1;  //214 / 163 = 1
    16'b11010110_10100100 : OUT <= 1;  //214 / 164 = 1
    16'b11010110_10100101 : OUT <= 1;  //214 / 165 = 1
    16'b11010110_10100110 : OUT <= 1;  //214 / 166 = 1
    16'b11010110_10100111 : OUT <= 1;  //214 / 167 = 1
    16'b11010110_10101000 : OUT <= 1;  //214 / 168 = 1
    16'b11010110_10101001 : OUT <= 1;  //214 / 169 = 1
    16'b11010110_10101010 : OUT <= 1;  //214 / 170 = 1
    16'b11010110_10101011 : OUT <= 1;  //214 / 171 = 1
    16'b11010110_10101100 : OUT <= 1;  //214 / 172 = 1
    16'b11010110_10101101 : OUT <= 1;  //214 / 173 = 1
    16'b11010110_10101110 : OUT <= 1;  //214 / 174 = 1
    16'b11010110_10101111 : OUT <= 1;  //214 / 175 = 1
    16'b11010110_10110000 : OUT <= 1;  //214 / 176 = 1
    16'b11010110_10110001 : OUT <= 1;  //214 / 177 = 1
    16'b11010110_10110010 : OUT <= 1;  //214 / 178 = 1
    16'b11010110_10110011 : OUT <= 1;  //214 / 179 = 1
    16'b11010110_10110100 : OUT <= 1;  //214 / 180 = 1
    16'b11010110_10110101 : OUT <= 1;  //214 / 181 = 1
    16'b11010110_10110110 : OUT <= 1;  //214 / 182 = 1
    16'b11010110_10110111 : OUT <= 1;  //214 / 183 = 1
    16'b11010110_10111000 : OUT <= 1;  //214 / 184 = 1
    16'b11010110_10111001 : OUT <= 1;  //214 / 185 = 1
    16'b11010110_10111010 : OUT <= 1;  //214 / 186 = 1
    16'b11010110_10111011 : OUT <= 1;  //214 / 187 = 1
    16'b11010110_10111100 : OUT <= 1;  //214 / 188 = 1
    16'b11010110_10111101 : OUT <= 1;  //214 / 189 = 1
    16'b11010110_10111110 : OUT <= 1;  //214 / 190 = 1
    16'b11010110_10111111 : OUT <= 1;  //214 / 191 = 1
    16'b11010110_11000000 : OUT <= 1;  //214 / 192 = 1
    16'b11010110_11000001 : OUT <= 1;  //214 / 193 = 1
    16'b11010110_11000010 : OUT <= 1;  //214 / 194 = 1
    16'b11010110_11000011 : OUT <= 1;  //214 / 195 = 1
    16'b11010110_11000100 : OUT <= 1;  //214 / 196 = 1
    16'b11010110_11000101 : OUT <= 1;  //214 / 197 = 1
    16'b11010110_11000110 : OUT <= 1;  //214 / 198 = 1
    16'b11010110_11000111 : OUT <= 1;  //214 / 199 = 1
    16'b11010110_11001000 : OUT <= 1;  //214 / 200 = 1
    16'b11010110_11001001 : OUT <= 1;  //214 / 201 = 1
    16'b11010110_11001010 : OUT <= 1;  //214 / 202 = 1
    16'b11010110_11001011 : OUT <= 1;  //214 / 203 = 1
    16'b11010110_11001100 : OUT <= 1;  //214 / 204 = 1
    16'b11010110_11001101 : OUT <= 1;  //214 / 205 = 1
    16'b11010110_11001110 : OUT <= 1;  //214 / 206 = 1
    16'b11010110_11001111 : OUT <= 1;  //214 / 207 = 1
    16'b11010110_11010000 : OUT <= 1;  //214 / 208 = 1
    16'b11010110_11010001 : OUT <= 1;  //214 / 209 = 1
    16'b11010110_11010010 : OUT <= 1;  //214 / 210 = 1
    16'b11010110_11010011 : OUT <= 1;  //214 / 211 = 1
    16'b11010110_11010100 : OUT <= 1;  //214 / 212 = 1
    16'b11010110_11010101 : OUT <= 1;  //214 / 213 = 1
    16'b11010110_11010110 : OUT <= 1;  //214 / 214 = 1
    16'b11010110_11010111 : OUT <= 0;  //214 / 215 = 0
    16'b11010110_11011000 : OUT <= 0;  //214 / 216 = 0
    16'b11010110_11011001 : OUT <= 0;  //214 / 217 = 0
    16'b11010110_11011010 : OUT <= 0;  //214 / 218 = 0
    16'b11010110_11011011 : OUT <= 0;  //214 / 219 = 0
    16'b11010110_11011100 : OUT <= 0;  //214 / 220 = 0
    16'b11010110_11011101 : OUT <= 0;  //214 / 221 = 0
    16'b11010110_11011110 : OUT <= 0;  //214 / 222 = 0
    16'b11010110_11011111 : OUT <= 0;  //214 / 223 = 0
    16'b11010110_11100000 : OUT <= 0;  //214 / 224 = 0
    16'b11010110_11100001 : OUT <= 0;  //214 / 225 = 0
    16'b11010110_11100010 : OUT <= 0;  //214 / 226 = 0
    16'b11010110_11100011 : OUT <= 0;  //214 / 227 = 0
    16'b11010110_11100100 : OUT <= 0;  //214 / 228 = 0
    16'b11010110_11100101 : OUT <= 0;  //214 / 229 = 0
    16'b11010110_11100110 : OUT <= 0;  //214 / 230 = 0
    16'b11010110_11100111 : OUT <= 0;  //214 / 231 = 0
    16'b11010110_11101000 : OUT <= 0;  //214 / 232 = 0
    16'b11010110_11101001 : OUT <= 0;  //214 / 233 = 0
    16'b11010110_11101010 : OUT <= 0;  //214 / 234 = 0
    16'b11010110_11101011 : OUT <= 0;  //214 / 235 = 0
    16'b11010110_11101100 : OUT <= 0;  //214 / 236 = 0
    16'b11010110_11101101 : OUT <= 0;  //214 / 237 = 0
    16'b11010110_11101110 : OUT <= 0;  //214 / 238 = 0
    16'b11010110_11101111 : OUT <= 0;  //214 / 239 = 0
    16'b11010110_11110000 : OUT <= 0;  //214 / 240 = 0
    16'b11010110_11110001 : OUT <= 0;  //214 / 241 = 0
    16'b11010110_11110010 : OUT <= 0;  //214 / 242 = 0
    16'b11010110_11110011 : OUT <= 0;  //214 / 243 = 0
    16'b11010110_11110100 : OUT <= 0;  //214 / 244 = 0
    16'b11010110_11110101 : OUT <= 0;  //214 / 245 = 0
    16'b11010110_11110110 : OUT <= 0;  //214 / 246 = 0
    16'b11010110_11110111 : OUT <= 0;  //214 / 247 = 0
    16'b11010110_11111000 : OUT <= 0;  //214 / 248 = 0
    16'b11010110_11111001 : OUT <= 0;  //214 / 249 = 0
    16'b11010110_11111010 : OUT <= 0;  //214 / 250 = 0
    16'b11010110_11111011 : OUT <= 0;  //214 / 251 = 0
    16'b11010110_11111100 : OUT <= 0;  //214 / 252 = 0
    16'b11010110_11111101 : OUT <= 0;  //214 / 253 = 0
    16'b11010110_11111110 : OUT <= 0;  //214 / 254 = 0
    16'b11010110_11111111 : OUT <= 0;  //214 / 255 = 0
    16'b11010111_00000000 : OUT <= 0;  //215 / 0 = 0
    16'b11010111_00000001 : OUT <= 215;  //215 / 1 = 215
    16'b11010111_00000010 : OUT <= 107;  //215 / 2 = 107
    16'b11010111_00000011 : OUT <= 71;  //215 / 3 = 71
    16'b11010111_00000100 : OUT <= 53;  //215 / 4 = 53
    16'b11010111_00000101 : OUT <= 43;  //215 / 5 = 43
    16'b11010111_00000110 : OUT <= 35;  //215 / 6 = 35
    16'b11010111_00000111 : OUT <= 30;  //215 / 7 = 30
    16'b11010111_00001000 : OUT <= 26;  //215 / 8 = 26
    16'b11010111_00001001 : OUT <= 23;  //215 / 9 = 23
    16'b11010111_00001010 : OUT <= 21;  //215 / 10 = 21
    16'b11010111_00001011 : OUT <= 19;  //215 / 11 = 19
    16'b11010111_00001100 : OUT <= 17;  //215 / 12 = 17
    16'b11010111_00001101 : OUT <= 16;  //215 / 13 = 16
    16'b11010111_00001110 : OUT <= 15;  //215 / 14 = 15
    16'b11010111_00001111 : OUT <= 14;  //215 / 15 = 14
    16'b11010111_00010000 : OUT <= 13;  //215 / 16 = 13
    16'b11010111_00010001 : OUT <= 12;  //215 / 17 = 12
    16'b11010111_00010010 : OUT <= 11;  //215 / 18 = 11
    16'b11010111_00010011 : OUT <= 11;  //215 / 19 = 11
    16'b11010111_00010100 : OUT <= 10;  //215 / 20 = 10
    16'b11010111_00010101 : OUT <= 10;  //215 / 21 = 10
    16'b11010111_00010110 : OUT <= 9;  //215 / 22 = 9
    16'b11010111_00010111 : OUT <= 9;  //215 / 23 = 9
    16'b11010111_00011000 : OUT <= 8;  //215 / 24 = 8
    16'b11010111_00011001 : OUT <= 8;  //215 / 25 = 8
    16'b11010111_00011010 : OUT <= 8;  //215 / 26 = 8
    16'b11010111_00011011 : OUT <= 7;  //215 / 27 = 7
    16'b11010111_00011100 : OUT <= 7;  //215 / 28 = 7
    16'b11010111_00011101 : OUT <= 7;  //215 / 29 = 7
    16'b11010111_00011110 : OUT <= 7;  //215 / 30 = 7
    16'b11010111_00011111 : OUT <= 6;  //215 / 31 = 6
    16'b11010111_00100000 : OUT <= 6;  //215 / 32 = 6
    16'b11010111_00100001 : OUT <= 6;  //215 / 33 = 6
    16'b11010111_00100010 : OUT <= 6;  //215 / 34 = 6
    16'b11010111_00100011 : OUT <= 6;  //215 / 35 = 6
    16'b11010111_00100100 : OUT <= 5;  //215 / 36 = 5
    16'b11010111_00100101 : OUT <= 5;  //215 / 37 = 5
    16'b11010111_00100110 : OUT <= 5;  //215 / 38 = 5
    16'b11010111_00100111 : OUT <= 5;  //215 / 39 = 5
    16'b11010111_00101000 : OUT <= 5;  //215 / 40 = 5
    16'b11010111_00101001 : OUT <= 5;  //215 / 41 = 5
    16'b11010111_00101010 : OUT <= 5;  //215 / 42 = 5
    16'b11010111_00101011 : OUT <= 5;  //215 / 43 = 5
    16'b11010111_00101100 : OUT <= 4;  //215 / 44 = 4
    16'b11010111_00101101 : OUT <= 4;  //215 / 45 = 4
    16'b11010111_00101110 : OUT <= 4;  //215 / 46 = 4
    16'b11010111_00101111 : OUT <= 4;  //215 / 47 = 4
    16'b11010111_00110000 : OUT <= 4;  //215 / 48 = 4
    16'b11010111_00110001 : OUT <= 4;  //215 / 49 = 4
    16'b11010111_00110010 : OUT <= 4;  //215 / 50 = 4
    16'b11010111_00110011 : OUT <= 4;  //215 / 51 = 4
    16'b11010111_00110100 : OUT <= 4;  //215 / 52 = 4
    16'b11010111_00110101 : OUT <= 4;  //215 / 53 = 4
    16'b11010111_00110110 : OUT <= 3;  //215 / 54 = 3
    16'b11010111_00110111 : OUT <= 3;  //215 / 55 = 3
    16'b11010111_00111000 : OUT <= 3;  //215 / 56 = 3
    16'b11010111_00111001 : OUT <= 3;  //215 / 57 = 3
    16'b11010111_00111010 : OUT <= 3;  //215 / 58 = 3
    16'b11010111_00111011 : OUT <= 3;  //215 / 59 = 3
    16'b11010111_00111100 : OUT <= 3;  //215 / 60 = 3
    16'b11010111_00111101 : OUT <= 3;  //215 / 61 = 3
    16'b11010111_00111110 : OUT <= 3;  //215 / 62 = 3
    16'b11010111_00111111 : OUT <= 3;  //215 / 63 = 3
    16'b11010111_01000000 : OUT <= 3;  //215 / 64 = 3
    16'b11010111_01000001 : OUT <= 3;  //215 / 65 = 3
    16'b11010111_01000010 : OUT <= 3;  //215 / 66 = 3
    16'b11010111_01000011 : OUT <= 3;  //215 / 67 = 3
    16'b11010111_01000100 : OUT <= 3;  //215 / 68 = 3
    16'b11010111_01000101 : OUT <= 3;  //215 / 69 = 3
    16'b11010111_01000110 : OUT <= 3;  //215 / 70 = 3
    16'b11010111_01000111 : OUT <= 3;  //215 / 71 = 3
    16'b11010111_01001000 : OUT <= 2;  //215 / 72 = 2
    16'b11010111_01001001 : OUT <= 2;  //215 / 73 = 2
    16'b11010111_01001010 : OUT <= 2;  //215 / 74 = 2
    16'b11010111_01001011 : OUT <= 2;  //215 / 75 = 2
    16'b11010111_01001100 : OUT <= 2;  //215 / 76 = 2
    16'b11010111_01001101 : OUT <= 2;  //215 / 77 = 2
    16'b11010111_01001110 : OUT <= 2;  //215 / 78 = 2
    16'b11010111_01001111 : OUT <= 2;  //215 / 79 = 2
    16'b11010111_01010000 : OUT <= 2;  //215 / 80 = 2
    16'b11010111_01010001 : OUT <= 2;  //215 / 81 = 2
    16'b11010111_01010010 : OUT <= 2;  //215 / 82 = 2
    16'b11010111_01010011 : OUT <= 2;  //215 / 83 = 2
    16'b11010111_01010100 : OUT <= 2;  //215 / 84 = 2
    16'b11010111_01010101 : OUT <= 2;  //215 / 85 = 2
    16'b11010111_01010110 : OUT <= 2;  //215 / 86 = 2
    16'b11010111_01010111 : OUT <= 2;  //215 / 87 = 2
    16'b11010111_01011000 : OUT <= 2;  //215 / 88 = 2
    16'b11010111_01011001 : OUT <= 2;  //215 / 89 = 2
    16'b11010111_01011010 : OUT <= 2;  //215 / 90 = 2
    16'b11010111_01011011 : OUT <= 2;  //215 / 91 = 2
    16'b11010111_01011100 : OUT <= 2;  //215 / 92 = 2
    16'b11010111_01011101 : OUT <= 2;  //215 / 93 = 2
    16'b11010111_01011110 : OUT <= 2;  //215 / 94 = 2
    16'b11010111_01011111 : OUT <= 2;  //215 / 95 = 2
    16'b11010111_01100000 : OUT <= 2;  //215 / 96 = 2
    16'b11010111_01100001 : OUT <= 2;  //215 / 97 = 2
    16'b11010111_01100010 : OUT <= 2;  //215 / 98 = 2
    16'b11010111_01100011 : OUT <= 2;  //215 / 99 = 2
    16'b11010111_01100100 : OUT <= 2;  //215 / 100 = 2
    16'b11010111_01100101 : OUT <= 2;  //215 / 101 = 2
    16'b11010111_01100110 : OUT <= 2;  //215 / 102 = 2
    16'b11010111_01100111 : OUT <= 2;  //215 / 103 = 2
    16'b11010111_01101000 : OUT <= 2;  //215 / 104 = 2
    16'b11010111_01101001 : OUT <= 2;  //215 / 105 = 2
    16'b11010111_01101010 : OUT <= 2;  //215 / 106 = 2
    16'b11010111_01101011 : OUT <= 2;  //215 / 107 = 2
    16'b11010111_01101100 : OUT <= 1;  //215 / 108 = 1
    16'b11010111_01101101 : OUT <= 1;  //215 / 109 = 1
    16'b11010111_01101110 : OUT <= 1;  //215 / 110 = 1
    16'b11010111_01101111 : OUT <= 1;  //215 / 111 = 1
    16'b11010111_01110000 : OUT <= 1;  //215 / 112 = 1
    16'b11010111_01110001 : OUT <= 1;  //215 / 113 = 1
    16'b11010111_01110010 : OUT <= 1;  //215 / 114 = 1
    16'b11010111_01110011 : OUT <= 1;  //215 / 115 = 1
    16'b11010111_01110100 : OUT <= 1;  //215 / 116 = 1
    16'b11010111_01110101 : OUT <= 1;  //215 / 117 = 1
    16'b11010111_01110110 : OUT <= 1;  //215 / 118 = 1
    16'b11010111_01110111 : OUT <= 1;  //215 / 119 = 1
    16'b11010111_01111000 : OUT <= 1;  //215 / 120 = 1
    16'b11010111_01111001 : OUT <= 1;  //215 / 121 = 1
    16'b11010111_01111010 : OUT <= 1;  //215 / 122 = 1
    16'b11010111_01111011 : OUT <= 1;  //215 / 123 = 1
    16'b11010111_01111100 : OUT <= 1;  //215 / 124 = 1
    16'b11010111_01111101 : OUT <= 1;  //215 / 125 = 1
    16'b11010111_01111110 : OUT <= 1;  //215 / 126 = 1
    16'b11010111_01111111 : OUT <= 1;  //215 / 127 = 1
    16'b11010111_10000000 : OUT <= 1;  //215 / 128 = 1
    16'b11010111_10000001 : OUT <= 1;  //215 / 129 = 1
    16'b11010111_10000010 : OUT <= 1;  //215 / 130 = 1
    16'b11010111_10000011 : OUT <= 1;  //215 / 131 = 1
    16'b11010111_10000100 : OUT <= 1;  //215 / 132 = 1
    16'b11010111_10000101 : OUT <= 1;  //215 / 133 = 1
    16'b11010111_10000110 : OUT <= 1;  //215 / 134 = 1
    16'b11010111_10000111 : OUT <= 1;  //215 / 135 = 1
    16'b11010111_10001000 : OUT <= 1;  //215 / 136 = 1
    16'b11010111_10001001 : OUT <= 1;  //215 / 137 = 1
    16'b11010111_10001010 : OUT <= 1;  //215 / 138 = 1
    16'b11010111_10001011 : OUT <= 1;  //215 / 139 = 1
    16'b11010111_10001100 : OUT <= 1;  //215 / 140 = 1
    16'b11010111_10001101 : OUT <= 1;  //215 / 141 = 1
    16'b11010111_10001110 : OUT <= 1;  //215 / 142 = 1
    16'b11010111_10001111 : OUT <= 1;  //215 / 143 = 1
    16'b11010111_10010000 : OUT <= 1;  //215 / 144 = 1
    16'b11010111_10010001 : OUT <= 1;  //215 / 145 = 1
    16'b11010111_10010010 : OUT <= 1;  //215 / 146 = 1
    16'b11010111_10010011 : OUT <= 1;  //215 / 147 = 1
    16'b11010111_10010100 : OUT <= 1;  //215 / 148 = 1
    16'b11010111_10010101 : OUT <= 1;  //215 / 149 = 1
    16'b11010111_10010110 : OUT <= 1;  //215 / 150 = 1
    16'b11010111_10010111 : OUT <= 1;  //215 / 151 = 1
    16'b11010111_10011000 : OUT <= 1;  //215 / 152 = 1
    16'b11010111_10011001 : OUT <= 1;  //215 / 153 = 1
    16'b11010111_10011010 : OUT <= 1;  //215 / 154 = 1
    16'b11010111_10011011 : OUT <= 1;  //215 / 155 = 1
    16'b11010111_10011100 : OUT <= 1;  //215 / 156 = 1
    16'b11010111_10011101 : OUT <= 1;  //215 / 157 = 1
    16'b11010111_10011110 : OUT <= 1;  //215 / 158 = 1
    16'b11010111_10011111 : OUT <= 1;  //215 / 159 = 1
    16'b11010111_10100000 : OUT <= 1;  //215 / 160 = 1
    16'b11010111_10100001 : OUT <= 1;  //215 / 161 = 1
    16'b11010111_10100010 : OUT <= 1;  //215 / 162 = 1
    16'b11010111_10100011 : OUT <= 1;  //215 / 163 = 1
    16'b11010111_10100100 : OUT <= 1;  //215 / 164 = 1
    16'b11010111_10100101 : OUT <= 1;  //215 / 165 = 1
    16'b11010111_10100110 : OUT <= 1;  //215 / 166 = 1
    16'b11010111_10100111 : OUT <= 1;  //215 / 167 = 1
    16'b11010111_10101000 : OUT <= 1;  //215 / 168 = 1
    16'b11010111_10101001 : OUT <= 1;  //215 / 169 = 1
    16'b11010111_10101010 : OUT <= 1;  //215 / 170 = 1
    16'b11010111_10101011 : OUT <= 1;  //215 / 171 = 1
    16'b11010111_10101100 : OUT <= 1;  //215 / 172 = 1
    16'b11010111_10101101 : OUT <= 1;  //215 / 173 = 1
    16'b11010111_10101110 : OUT <= 1;  //215 / 174 = 1
    16'b11010111_10101111 : OUT <= 1;  //215 / 175 = 1
    16'b11010111_10110000 : OUT <= 1;  //215 / 176 = 1
    16'b11010111_10110001 : OUT <= 1;  //215 / 177 = 1
    16'b11010111_10110010 : OUT <= 1;  //215 / 178 = 1
    16'b11010111_10110011 : OUT <= 1;  //215 / 179 = 1
    16'b11010111_10110100 : OUT <= 1;  //215 / 180 = 1
    16'b11010111_10110101 : OUT <= 1;  //215 / 181 = 1
    16'b11010111_10110110 : OUT <= 1;  //215 / 182 = 1
    16'b11010111_10110111 : OUT <= 1;  //215 / 183 = 1
    16'b11010111_10111000 : OUT <= 1;  //215 / 184 = 1
    16'b11010111_10111001 : OUT <= 1;  //215 / 185 = 1
    16'b11010111_10111010 : OUT <= 1;  //215 / 186 = 1
    16'b11010111_10111011 : OUT <= 1;  //215 / 187 = 1
    16'b11010111_10111100 : OUT <= 1;  //215 / 188 = 1
    16'b11010111_10111101 : OUT <= 1;  //215 / 189 = 1
    16'b11010111_10111110 : OUT <= 1;  //215 / 190 = 1
    16'b11010111_10111111 : OUT <= 1;  //215 / 191 = 1
    16'b11010111_11000000 : OUT <= 1;  //215 / 192 = 1
    16'b11010111_11000001 : OUT <= 1;  //215 / 193 = 1
    16'b11010111_11000010 : OUT <= 1;  //215 / 194 = 1
    16'b11010111_11000011 : OUT <= 1;  //215 / 195 = 1
    16'b11010111_11000100 : OUT <= 1;  //215 / 196 = 1
    16'b11010111_11000101 : OUT <= 1;  //215 / 197 = 1
    16'b11010111_11000110 : OUT <= 1;  //215 / 198 = 1
    16'b11010111_11000111 : OUT <= 1;  //215 / 199 = 1
    16'b11010111_11001000 : OUT <= 1;  //215 / 200 = 1
    16'b11010111_11001001 : OUT <= 1;  //215 / 201 = 1
    16'b11010111_11001010 : OUT <= 1;  //215 / 202 = 1
    16'b11010111_11001011 : OUT <= 1;  //215 / 203 = 1
    16'b11010111_11001100 : OUT <= 1;  //215 / 204 = 1
    16'b11010111_11001101 : OUT <= 1;  //215 / 205 = 1
    16'b11010111_11001110 : OUT <= 1;  //215 / 206 = 1
    16'b11010111_11001111 : OUT <= 1;  //215 / 207 = 1
    16'b11010111_11010000 : OUT <= 1;  //215 / 208 = 1
    16'b11010111_11010001 : OUT <= 1;  //215 / 209 = 1
    16'b11010111_11010010 : OUT <= 1;  //215 / 210 = 1
    16'b11010111_11010011 : OUT <= 1;  //215 / 211 = 1
    16'b11010111_11010100 : OUT <= 1;  //215 / 212 = 1
    16'b11010111_11010101 : OUT <= 1;  //215 / 213 = 1
    16'b11010111_11010110 : OUT <= 1;  //215 / 214 = 1
    16'b11010111_11010111 : OUT <= 1;  //215 / 215 = 1
    16'b11010111_11011000 : OUT <= 0;  //215 / 216 = 0
    16'b11010111_11011001 : OUT <= 0;  //215 / 217 = 0
    16'b11010111_11011010 : OUT <= 0;  //215 / 218 = 0
    16'b11010111_11011011 : OUT <= 0;  //215 / 219 = 0
    16'b11010111_11011100 : OUT <= 0;  //215 / 220 = 0
    16'b11010111_11011101 : OUT <= 0;  //215 / 221 = 0
    16'b11010111_11011110 : OUT <= 0;  //215 / 222 = 0
    16'b11010111_11011111 : OUT <= 0;  //215 / 223 = 0
    16'b11010111_11100000 : OUT <= 0;  //215 / 224 = 0
    16'b11010111_11100001 : OUT <= 0;  //215 / 225 = 0
    16'b11010111_11100010 : OUT <= 0;  //215 / 226 = 0
    16'b11010111_11100011 : OUT <= 0;  //215 / 227 = 0
    16'b11010111_11100100 : OUT <= 0;  //215 / 228 = 0
    16'b11010111_11100101 : OUT <= 0;  //215 / 229 = 0
    16'b11010111_11100110 : OUT <= 0;  //215 / 230 = 0
    16'b11010111_11100111 : OUT <= 0;  //215 / 231 = 0
    16'b11010111_11101000 : OUT <= 0;  //215 / 232 = 0
    16'b11010111_11101001 : OUT <= 0;  //215 / 233 = 0
    16'b11010111_11101010 : OUT <= 0;  //215 / 234 = 0
    16'b11010111_11101011 : OUT <= 0;  //215 / 235 = 0
    16'b11010111_11101100 : OUT <= 0;  //215 / 236 = 0
    16'b11010111_11101101 : OUT <= 0;  //215 / 237 = 0
    16'b11010111_11101110 : OUT <= 0;  //215 / 238 = 0
    16'b11010111_11101111 : OUT <= 0;  //215 / 239 = 0
    16'b11010111_11110000 : OUT <= 0;  //215 / 240 = 0
    16'b11010111_11110001 : OUT <= 0;  //215 / 241 = 0
    16'b11010111_11110010 : OUT <= 0;  //215 / 242 = 0
    16'b11010111_11110011 : OUT <= 0;  //215 / 243 = 0
    16'b11010111_11110100 : OUT <= 0;  //215 / 244 = 0
    16'b11010111_11110101 : OUT <= 0;  //215 / 245 = 0
    16'b11010111_11110110 : OUT <= 0;  //215 / 246 = 0
    16'b11010111_11110111 : OUT <= 0;  //215 / 247 = 0
    16'b11010111_11111000 : OUT <= 0;  //215 / 248 = 0
    16'b11010111_11111001 : OUT <= 0;  //215 / 249 = 0
    16'b11010111_11111010 : OUT <= 0;  //215 / 250 = 0
    16'b11010111_11111011 : OUT <= 0;  //215 / 251 = 0
    16'b11010111_11111100 : OUT <= 0;  //215 / 252 = 0
    16'b11010111_11111101 : OUT <= 0;  //215 / 253 = 0
    16'b11010111_11111110 : OUT <= 0;  //215 / 254 = 0
    16'b11010111_11111111 : OUT <= 0;  //215 / 255 = 0
    16'b11011000_00000000 : OUT <= 0;  //216 / 0 = 0
    16'b11011000_00000001 : OUT <= 216;  //216 / 1 = 216
    16'b11011000_00000010 : OUT <= 108;  //216 / 2 = 108
    16'b11011000_00000011 : OUT <= 72;  //216 / 3 = 72
    16'b11011000_00000100 : OUT <= 54;  //216 / 4 = 54
    16'b11011000_00000101 : OUT <= 43;  //216 / 5 = 43
    16'b11011000_00000110 : OUT <= 36;  //216 / 6 = 36
    16'b11011000_00000111 : OUT <= 30;  //216 / 7 = 30
    16'b11011000_00001000 : OUT <= 27;  //216 / 8 = 27
    16'b11011000_00001001 : OUT <= 24;  //216 / 9 = 24
    16'b11011000_00001010 : OUT <= 21;  //216 / 10 = 21
    16'b11011000_00001011 : OUT <= 19;  //216 / 11 = 19
    16'b11011000_00001100 : OUT <= 18;  //216 / 12 = 18
    16'b11011000_00001101 : OUT <= 16;  //216 / 13 = 16
    16'b11011000_00001110 : OUT <= 15;  //216 / 14 = 15
    16'b11011000_00001111 : OUT <= 14;  //216 / 15 = 14
    16'b11011000_00010000 : OUT <= 13;  //216 / 16 = 13
    16'b11011000_00010001 : OUT <= 12;  //216 / 17 = 12
    16'b11011000_00010010 : OUT <= 12;  //216 / 18 = 12
    16'b11011000_00010011 : OUT <= 11;  //216 / 19 = 11
    16'b11011000_00010100 : OUT <= 10;  //216 / 20 = 10
    16'b11011000_00010101 : OUT <= 10;  //216 / 21 = 10
    16'b11011000_00010110 : OUT <= 9;  //216 / 22 = 9
    16'b11011000_00010111 : OUT <= 9;  //216 / 23 = 9
    16'b11011000_00011000 : OUT <= 9;  //216 / 24 = 9
    16'b11011000_00011001 : OUT <= 8;  //216 / 25 = 8
    16'b11011000_00011010 : OUT <= 8;  //216 / 26 = 8
    16'b11011000_00011011 : OUT <= 8;  //216 / 27 = 8
    16'b11011000_00011100 : OUT <= 7;  //216 / 28 = 7
    16'b11011000_00011101 : OUT <= 7;  //216 / 29 = 7
    16'b11011000_00011110 : OUT <= 7;  //216 / 30 = 7
    16'b11011000_00011111 : OUT <= 6;  //216 / 31 = 6
    16'b11011000_00100000 : OUT <= 6;  //216 / 32 = 6
    16'b11011000_00100001 : OUT <= 6;  //216 / 33 = 6
    16'b11011000_00100010 : OUT <= 6;  //216 / 34 = 6
    16'b11011000_00100011 : OUT <= 6;  //216 / 35 = 6
    16'b11011000_00100100 : OUT <= 6;  //216 / 36 = 6
    16'b11011000_00100101 : OUT <= 5;  //216 / 37 = 5
    16'b11011000_00100110 : OUT <= 5;  //216 / 38 = 5
    16'b11011000_00100111 : OUT <= 5;  //216 / 39 = 5
    16'b11011000_00101000 : OUT <= 5;  //216 / 40 = 5
    16'b11011000_00101001 : OUT <= 5;  //216 / 41 = 5
    16'b11011000_00101010 : OUT <= 5;  //216 / 42 = 5
    16'b11011000_00101011 : OUT <= 5;  //216 / 43 = 5
    16'b11011000_00101100 : OUT <= 4;  //216 / 44 = 4
    16'b11011000_00101101 : OUT <= 4;  //216 / 45 = 4
    16'b11011000_00101110 : OUT <= 4;  //216 / 46 = 4
    16'b11011000_00101111 : OUT <= 4;  //216 / 47 = 4
    16'b11011000_00110000 : OUT <= 4;  //216 / 48 = 4
    16'b11011000_00110001 : OUT <= 4;  //216 / 49 = 4
    16'b11011000_00110010 : OUT <= 4;  //216 / 50 = 4
    16'b11011000_00110011 : OUT <= 4;  //216 / 51 = 4
    16'b11011000_00110100 : OUT <= 4;  //216 / 52 = 4
    16'b11011000_00110101 : OUT <= 4;  //216 / 53 = 4
    16'b11011000_00110110 : OUT <= 4;  //216 / 54 = 4
    16'b11011000_00110111 : OUT <= 3;  //216 / 55 = 3
    16'b11011000_00111000 : OUT <= 3;  //216 / 56 = 3
    16'b11011000_00111001 : OUT <= 3;  //216 / 57 = 3
    16'b11011000_00111010 : OUT <= 3;  //216 / 58 = 3
    16'b11011000_00111011 : OUT <= 3;  //216 / 59 = 3
    16'b11011000_00111100 : OUT <= 3;  //216 / 60 = 3
    16'b11011000_00111101 : OUT <= 3;  //216 / 61 = 3
    16'b11011000_00111110 : OUT <= 3;  //216 / 62 = 3
    16'b11011000_00111111 : OUT <= 3;  //216 / 63 = 3
    16'b11011000_01000000 : OUT <= 3;  //216 / 64 = 3
    16'b11011000_01000001 : OUT <= 3;  //216 / 65 = 3
    16'b11011000_01000010 : OUT <= 3;  //216 / 66 = 3
    16'b11011000_01000011 : OUT <= 3;  //216 / 67 = 3
    16'b11011000_01000100 : OUT <= 3;  //216 / 68 = 3
    16'b11011000_01000101 : OUT <= 3;  //216 / 69 = 3
    16'b11011000_01000110 : OUT <= 3;  //216 / 70 = 3
    16'b11011000_01000111 : OUT <= 3;  //216 / 71 = 3
    16'b11011000_01001000 : OUT <= 3;  //216 / 72 = 3
    16'b11011000_01001001 : OUT <= 2;  //216 / 73 = 2
    16'b11011000_01001010 : OUT <= 2;  //216 / 74 = 2
    16'b11011000_01001011 : OUT <= 2;  //216 / 75 = 2
    16'b11011000_01001100 : OUT <= 2;  //216 / 76 = 2
    16'b11011000_01001101 : OUT <= 2;  //216 / 77 = 2
    16'b11011000_01001110 : OUT <= 2;  //216 / 78 = 2
    16'b11011000_01001111 : OUT <= 2;  //216 / 79 = 2
    16'b11011000_01010000 : OUT <= 2;  //216 / 80 = 2
    16'b11011000_01010001 : OUT <= 2;  //216 / 81 = 2
    16'b11011000_01010010 : OUT <= 2;  //216 / 82 = 2
    16'b11011000_01010011 : OUT <= 2;  //216 / 83 = 2
    16'b11011000_01010100 : OUT <= 2;  //216 / 84 = 2
    16'b11011000_01010101 : OUT <= 2;  //216 / 85 = 2
    16'b11011000_01010110 : OUT <= 2;  //216 / 86 = 2
    16'b11011000_01010111 : OUT <= 2;  //216 / 87 = 2
    16'b11011000_01011000 : OUT <= 2;  //216 / 88 = 2
    16'b11011000_01011001 : OUT <= 2;  //216 / 89 = 2
    16'b11011000_01011010 : OUT <= 2;  //216 / 90 = 2
    16'b11011000_01011011 : OUT <= 2;  //216 / 91 = 2
    16'b11011000_01011100 : OUT <= 2;  //216 / 92 = 2
    16'b11011000_01011101 : OUT <= 2;  //216 / 93 = 2
    16'b11011000_01011110 : OUT <= 2;  //216 / 94 = 2
    16'b11011000_01011111 : OUT <= 2;  //216 / 95 = 2
    16'b11011000_01100000 : OUT <= 2;  //216 / 96 = 2
    16'b11011000_01100001 : OUT <= 2;  //216 / 97 = 2
    16'b11011000_01100010 : OUT <= 2;  //216 / 98 = 2
    16'b11011000_01100011 : OUT <= 2;  //216 / 99 = 2
    16'b11011000_01100100 : OUT <= 2;  //216 / 100 = 2
    16'b11011000_01100101 : OUT <= 2;  //216 / 101 = 2
    16'b11011000_01100110 : OUT <= 2;  //216 / 102 = 2
    16'b11011000_01100111 : OUT <= 2;  //216 / 103 = 2
    16'b11011000_01101000 : OUT <= 2;  //216 / 104 = 2
    16'b11011000_01101001 : OUT <= 2;  //216 / 105 = 2
    16'b11011000_01101010 : OUT <= 2;  //216 / 106 = 2
    16'b11011000_01101011 : OUT <= 2;  //216 / 107 = 2
    16'b11011000_01101100 : OUT <= 2;  //216 / 108 = 2
    16'b11011000_01101101 : OUT <= 1;  //216 / 109 = 1
    16'b11011000_01101110 : OUT <= 1;  //216 / 110 = 1
    16'b11011000_01101111 : OUT <= 1;  //216 / 111 = 1
    16'b11011000_01110000 : OUT <= 1;  //216 / 112 = 1
    16'b11011000_01110001 : OUT <= 1;  //216 / 113 = 1
    16'b11011000_01110010 : OUT <= 1;  //216 / 114 = 1
    16'b11011000_01110011 : OUT <= 1;  //216 / 115 = 1
    16'b11011000_01110100 : OUT <= 1;  //216 / 116 = 1
    16'b11011000_01110101 : OUT <= 1;  //216 / 117 = 1
    16'b11011000_01110110 : OUT <= 1;  //216 / 118 = 1
    16'b11011000_01110111 : OUT <= 1;  //216 / 119 = 1
    16'b11011000_01111000 : OUT <= 1;  //216 / 120 = 1
    16'b11011000_01111001 : OUT <= 1;  //216 / 121 = 1
    16'b11011000_01111010 : OUT <= 1;  //216 / 122 = 1
    16'b11011000_01111011 : OUT <= 1;  //216 / 123 = 1
    16'b11011000_01111100 : OUT <= 1;  //216 / 124 = 1
    16'b11011000_01111101 : OUT <= 1;  //216 / 125 = 1
    16'b11011000_01111110 : OUT <= 1;  //216 / 126 = 1
    16'b11011000_01111111 : OUT <= 1;  //216 / 127 = 1
    16'b11011000_10000000 : OUT <= 1;  //216 / 128 = 1
    16'b11011000_10000001 : OUT <= 1;  //216 / 129 = 1
    16'b11011000_10000010 : OUT <= 1;  //216 / 130 = 1
    16'b11011000_10000011 : OUT <= 1;  //216 / 131 = 1
    16'b11011000_10000100 : OUT <= 1;  //216 / 132 = 1
    16'b11011000_10000101 : OUT <= 1;  //216 / 133 = 1
    16'b11011000_10000110 : OUT <= 1;  //216 / 134 = 1
    16'b11011000_10000111 : OUT <= 1;  //216 / 135 = 1
    16'b11011000_10001000 : OUT <= 1;  //216 / 136 = 1
    16'b11011000_10001001 : OUT <= 1;  //216 / 137 = 1
    16'b11011000_10001010 : OUT <= 1;  //216 / 138 = 1
    16'b11011000_10001011 : OUT <= 1;  //216 / 139 = 1
    16'b11011000_10001100 : OUT <= 1;  //216 / 140 = 1
    16'b11011000_10001101 : OUT <= 1;  //216 / 141 = 1
    16'b11011000_10001110 : OUT <= 1;  //216 / 142 = 1
    16'b11011000_10001111 : OUT <= 1;  //216 / 143 = 1
    16'b11011000_10010000 : OUT <= 1;  //216 / 144 = 1
    16'b11011000_10010001 : OUT <= 1;  //216 / 145 = 1
    16'b11011000_10010010 : OUT <= 1;  //216 / 146 = 1
    16'b11011000_10010011 : OUT <= 1;  //216 / 147 = 1
    16'b11011000_10010100 : OUT <= 1;  //216 / 148 = 1
    16'b11011000_10010101 : OUT <= 1;  //216 / 149 = 1
    16'b11011000_10010110 : OUT <= 1;  //216 / 150 = 1
    16'b11011000_10010111 : OUT <= 1;  //216 / 151 = 1
    16'b11011000_10011000 : OUT <= 1;  //216 / 152 = 1
    16'b11011000_10011001 : OUT <= 1;  //216 / 153 = 1
    16'b11011000_10011010 : OUT <= 1;  //216 / 154 = 1
    16'b11011000_10011011 : OUT <= 1;  //216 / 155 = 1
    16'b11011000_10011100 : OUT <= 1;  //216 / 156 = 1
    16'b11011000_10011101 : OUT <= 1;  //216 / 157 = 1
    16'b11011000_10011110 : OUT <= 1;  //216 / 158 = 1
    16'b11011000_10011111 : OUT <= 1;  //216 / 159 = 1
    16'b11011000_10100000 : OUT <= 1;  //216 / 160 = 1
    16'b11011000_10100001 : OUT <= 1;  //216 / 161 = 1
    16'b11011000_10100010 : OUT <= 1;  //216 / 162 = 1
    16'b11011000_10100011 : OUT <= 1;  //216 / 163 = 1
    16'b11011000_10100100 : OUT <= 1;  //216 / 164 = 1
    16'b11011000_10100101 : OUT <= 1;  //216 / 165 = 1
    16'b11011000_10100110 : OUT <= 1;  //216 / 166 = 1
    16'b11011000_10100111 : OUT <= 1;  //216 / 167 = 1
    16'b11011000_10101000 : OUT <= 1;  //216 / 168 = 1
    16'b11011000_10101001 : OUT <= 1;  //216 / 169 = 1
    16'b11011000_10101010 : OUT <= 1;  //216 / 170 = 1
    16'b11011000_10101011 : OUT <= 1;  //216 / 171 = 1
    16'b11011000_10101100 : OUT <= 1;  //216 / 172 = 1
    16'b11011000_10101101 : OUT <= 1;  //216 / 173 = 1
    16'b11011000_10101110 : OUT <= 1;  //216 / 174 = 1
    16'b11011000_10101111 : OUT <= 1;  //216 / 175 = 1
    16'b11011000_10110000 : OUT <= 1;  //216 / 176 = 1
    16'b11011000_10110001 : OUT <= 1;  //216 / 177 = 1
    16'b11011000_10110010 : OUT <= 1;  //216 / 178 = 1
    16'b11011000_10110011 : OUT <= 1;  //216 / 179 = 1
    16'b11011000_10110100 : OUT <= 1;  //216 / 180 = 1
    16'b11011000_10110101 : OUT <= 1;  //216 / 181 = 1
    16'b11011000_10110110 : OUT <= 1;  //216 / 182 = 1
    16'b11011000_10110111 : OUT <= 1;  //216 / 183 = 1
    16'b11011000_10111000 : OUT <= 1;  //216 / 184 = 1
    16'b11011000_10111001 : OUT <= 1;  //216 / 185 = 1
    16'b11011000_10111010 : OUT <= 1;  //216 / 186 = 1
    16'b11011000_10111011 : OUT <= 1;  //216 / 187 = 1
    16'b11011000_10111100 : OUT <= 1;  //216 / 188 = 1
    16'b11011000_10111101 : OUT <= 1;  //216 / 189 = 1
    16'b11011000_10111110 : OUT <= 1;  //216 / 190 = 1
    16'b11011000_10111111 : OUT <= 1;  //216 / 191 = 1
    16'b11011000_11000000 : OUT <= 1;  //216 / 192 = 1
    16'b11011000_11000001 : OUT <= 1;  //216 / 193 = 1
    16'b11011000_11000010 : OUT <= 1;  //216 / 194 = 1
    16'b11011000_11000011 : OUT <= 1;  //216 / 195 = 1
    16'b11011000_11000100 : OUT <= 1;  //216 / 196 = 1
    16'b11011000_11000101 : OUT <= 1;  //216 / 197 = 1
    16'b11011000_11000110 : OUT <= 1;  //216 / 198 = 1
    16'b11011000_11000111 : OUT <= 1;  //216 / 199 = 1
    16'b11011000_11001000 : OUT <= 1;  //216 / 200 = 1
    16'b11011000_11001001 : OUT <= 1;  //216 / 201 = 1
    16'b11011000_11001010 : OUT <= 1;  //216 / 202 = 1
    16'b11011000_11001011 : OUT <= 1;  //216 / 203 = 1
    16'b11011000_11001100 : OUT <= 1;  //216 / 204 = 1
    16'b11011000_11001101 : OUT <= 1;  //216 / 205 = 1
    16'b11011000_11001110 : OUT <= 1;  //216 / 206 = 1
    16'b11011000_11001111 : OUT <= 1;  //216 / 207 = 1
    16'b11011000_11010000 : OUT <= 1;  //216 / 208 = 1
    16'b11011000_11010001 : OUT <= 1;  //216 / 209 = 1
    16'b11011000_11010010 : OUT <= 1;  //216 / 210 = 1
    16'b11011000_11010011 : OUT <= 1;  //216 / 211 = 1
    16'b11011000_11010100 : OUT <= 1;  //216 / 212 = 1
    16'b11011000_11010101 : OUT <= 1;  //216 / 213 = 1
    16'b11011000_11010110 : OUT <= 1;  //216 / 214 = 1
    16'b11011000_11010111 : OUT <= 1;  //216 / 215 = 1
    16'b11011000_11011000 : OUT <= 1;  //216 / 216 = 1
    16'b11011000_11011001 : OUT <= 0;  //216 / 217 = 0
    16'b11011000_11011010 : OUT <= 0;  //216 / 218 = 0
    16'b11011000_11011011 : OUT <= 0;  //216 / 219 = 0
    16'b11011000_11011100 : OUT <= 0;  //216 / 220 = 0
    16'b11011000_11011101 : OUT <= 0;  //216 / 221 = 0
    16'b11011000_11011110 : OUT <= 0;  //216 / 222 = 0
    16'b11011000_11011111 : OUT <= 0;  //216 / 223 = 0
    16'b11011000_11100000 : OUT <= 0;  //216 / 224 = 0
    16'b11011000_11100001 : OUT <= 0;  //216 / 225 = 0
    16'b11011000_11100010 : OUT <= 0;  //216 / 226 = 0
    16'b11011000_11100011 : OUT <= 0;  //216 / 227 = 0
    16'b11011000_11100100 : OUT <= 0;  //216 / 228 = 0
    16'b11011000_11100101 : OUT <= 0;  //216 / 229 = 0
    16'b11011000_11100110 : OUT <= 0;  //216 / 230 = 0
    16'b11011000_11100111 : OUT <= 0;  //216 / 231 = 0
    16'b11011000_11101000 : OUT <= 0;  //216 / 232 = 0
    16'b11011000_11101001 : OUT <= 0;  //216 / 233 = 0
    16'b11011000_11101010 : OUT <= 0;  //216 / 234 = 0
    16'b11011000_11101011 : OUT <= 0;  //216 / 235 = 0
    16'b11011000_11101100 : OUT <= 0;  //216 / 236 = 0
    16'b11011000_11101101 : OUT <= 0;  //216 / 237 = 0
    16'b11011000_11101110 : OUT <= 0;  //216 / 238 = 0
    16'b11011000_11101111 : OUT <= 0;  //216 / 239 = 0
    16'b11011000_11110000 : OUT <= 0;  //216 / 240 = 0
    16'b11011000_11110001 : OUT <= 0;  //216 / 241 = 0
    16'b11011000_11110010 : OUT <= 0;  //216 / 242 = 0
    16'b11011000_11110011 : OUT <= 0;  //216 / 243 = 0
    16'b11011000_11110100 : OUT <= 0;  //216 / 244 = 0
    16'b11011000_11110101 : OUT <= 0;  //216 / 245 = 0
    16'b11011000_11110110 : OUT <= 0;  //216 / 246 = 0
    16'b11011000_11110111 : OUT <= 0;  //216 / 247 = 0
    16'b11011000_11111000 : OUT <= 0;  //216 / 248 = 0
    16'b11011000_11111001 : OUT <= 0;  //216 / 249 = 0
    16'b11011000_11111010 : OUT <= 0;  //216 / 250 = 0
    16'b11011000_11111011 : OUT <= 0;  //216 / 251 = 0
    16'b11011000_11111100 : OUT <= 0;  //216 / 252 = 0
    16'b11011000_11111101 : OUT <= 0;  //216 / 253 = 0
    16'b11011000_11111110 : OUT <= 0;  //216 / 254 = 0
    16'b11011000_11111111 : OUT <= 0;  //216 / 255 = 0
    16'b11011001_00000000 : OUT <= 0;  //217 / 0 = 0
    16'b11011001_00000001 : OUT <= 217;  //217 / 1 = 217
    16'b11011001_00000010 : OUT <= 108;  //217 / 2 = 108
    16'b11011001_00000011 : OUT <= 72;  //217 / 3 = 72
    16'b11011001_00000100 : OUT <= 54;  //217 / 4 = 54
    16'b11011001_00000101 : OUT <= 43;  //217 / 5 = 43
    16'b11011001_00000110 : OUT <= 36;  //217 / 6 = 36
    16'b11011001_00000111 : OUT <= 31;  //217 / 7 = 31
    16'b11011001_00001000 : OUT <= 27;  //217 / 8 = 27
    16'b11011001_00001001 : OUT <= 24;  //217 / 9 = 24
    16'b11011001_00001010 : OUT <= 21;  //217 / 10 = 21
    16'b11011001_00001011 : OUT <= 19;  //217 / 11 = 19
    16'b11011001_00001100 : OUT <= 18;  //217 / 12 = 18
    16'b11011001_00001101 : OUT <= 16;  //217 / 13 = 16
    16'b11011001_00001110 : OUT <= 15;  //217 / 14 = 15
    16'b11011001_00001111 : OUT <= 14;  //217 / 15 = 14
    16'b11011001_00010000 : OUT <= 13;  //217 / 16 = 13
    16'b11011001_00010001 : OUT <= 12;  //217 / 17 = 12
    16'b11011001_00010010 : OUT <= 12;  //217 / 18 = 12
    16'b11011001_00010011 : OUT <= 11;  //217 / 19 = 11
    16'b11011001_00010100 : OUT <= 10;  //217 / 20 = 10
    16'b11011001_00010101 : OUT <= 10;  //217 / 21 = 10
    16'b11011001_00010110 : OUT <= 9;  //217 / 22 = 9
    16'b11011001_00010111 : OUT <= 9;  //217 / 23 = 9
    16'b11011001_00011000 : OUT <= 9;  //217 / 24 = 9
    16'b11011001_00011001 : OUT <= 8;  //217 / 25 = 8
    16'b11011001_00011010 : OUT <= 8;  //217 / 26 = 8
    16'b11011001_00011011 : OUT <= 8;  //217 / 27 = 8
    16'b11011001_00011100 : OUT <= 7;  //217 / 28 = 7
    16'b11011001_00011101 : OUT <= 7;  //217 / 29 = 7
    16'b11011001_00011110 : OUT <= 7;  //217 / 30 = 7
    16'b11011001_00011111 : OUT <= 7;  //217 / 31 = 7
    16'b11011001_00100000 : OUT <= 6;  //217 / 32 = 6
    16'b11011001_00100001 : OUT <= 6;  //217 / 33 = 6
    16'b11011001_00100010 : OUT <= 6;  //217 / 34 = 6
    16'b11011001_00100011 : OUT <= 6;  //217 / 35 = 6
    16'b11011001_00100100 : OUT <= 6;  //217 / 36 = 6
    16'b11011001_00100101 : OUT <= 5;  //217 / 37 = 5
    16'b11011001_00100110 : OUT <= 5;  //217 / 38 = 5
    16'b11011001_00100111 : OUT <= 5;  //217 / 39 = 5
    16'b11011001_00101000 : OUT <= 5;  //217 / 40 = 5
    16'b11011001_00101001 : OUT <= 5;  //217 / 41 = 5
    16'b11011001_00101010 : OUT <= 5;  //217 / 42 = 5
    16'b11011001_00101011 : OUT <= 5;  //217 / 43 = 5
    16'b11011001_00101100 : OUT <= 4;  //217 / 44 = 4
    16'b11011001_00101101 : OUT <= 4;  //217 / 45 = 4
    16'b11011001_00101110 : OUT <= 4;  //217 / 46 = 4
    16'b11011001_00101111 : OUT <= 4;  //217 / 47 = 4
    16'b11011001_00110000 : OUT <= 4;  //217 / 48 = 4
    16'b11011001_00110001 : OUT <= 4;  //217 / 49 = 4
    16'b11011001_00110010 : OUT <= 4;  //217 / 50 = 4
    16'b11011001_00110011 : OUT <= 4;  //217 / 51 = 4
    16'b11011001_00110100 : OUT <= 4;  //217 / 52 = 4
    16'b11011001_00110101 : OUT <= 4;  //217 / 53 = 4
    16'b11011001_00110110 : OUT <= 4;  //217 / 54 = 4
    16'b11011001_00110111 : OUT <= 3;  //217 / 55 = 3
    16'b11011001_00111000 : OUT <= 3;  //217 / 56 = 3
    16'b11011001_00111001 : OUT <= 3;  //217 / 57 = 3
    16'b11011001_00111010 : OUT <= 3;  //217 / 58 = 3
    16'b11011001_00111011 : OUT <= 3;  //217 / 59 = 3
    16'b11011001_00111100 : OUT <= 3;  //217 / 60 = 3
    16'b11011001_00111101 : OUT <= 3;  //217 / 61 = 3
    16'b11011001_00111110 : OUT <= 3;  //217 / 62 = 3
    16'b11011001_00111111 : OUT <= 3;  //217 / 63 = 3
    16'b11011001_01000000 : OUT <= 3;  //217 / 64 = 3
    16'b11011001_01000001 : OUT <= 3;  //217 / 65 = 3
    16'b11011001_01000010 : OUT <= 3;  //217 / 66 = 3
    16'b11011001_01000011 : OUT <= 3;  //217 / 67 = 3
    16'b11011001_01000100 : OUT <= 3;  //217 / 68 = 3
    16'b11011001_01000101 : OUT <= 3;  //217 / 69 = 3
    16'b11011001_01000110 : OUT <= 3;  //217 / 70 = 3
    16'b11011001_01000111 : OUT <= 3;  //217 / 71 = 3
    16'b11011001_01001000 : OUT <= 3;  //217 / 72 = 3
    16'b11011001_01001001 : OUT <= 2;  //217 / 73 = 2
    16'b11011001_01001010 : OUT <= 2;  //217 / 74 = 2
    16'b11011001_01001011 : OUT <= 2;  //217 / 75 = 2
    16'b11011001_01001100 : OUT <= 2;  //217 / 76 = 2
    16'b11011001_01001101 : OUT <= 2;  //217 / 77 = 2
    16'b11011001_01001110 : OUT <= 2;  //217 / 78 = 2
    16'b11011001_01001111 : OUT <= 2;  //217 / 79 = 2
    16'b11011001_01010000 : OUT <= 2;  //217 / 80 = 2
    16'b11011001_01010001 : OUT <= 2;  //217 / 81 = 2
    16'b11011001_01010010 : OUT <= 2;  //217 / 82 = 2
    16'b11011001_01010011 : OUT <= 2;  //217 / 83 = 2
    16'b11011001_01010100 : OUT <= 2;  //217 / 84 = 2
    16'b11011001_01010101 : OUT <= 2;  //217 / 85 = 2
    16'b11011001_01010110 : OUT <= 2;  //217 / 86 = 2
    16'b11011001_01010111 : OUT <= 2;  //217 / 87 = 2
    16'b11011001_01011000 : OUT <= 2;  //217 / 88 = 2
    16'b11011001_01011001 : OUT <= 2;  //217 / 89 = 2
    16'b11011001_01011010 : OUT <= 2;  //217 / 90 = 2
    16'b11011001_01011011 : OUT <= 2;  //217 / 91 = 2
    16'b11011001_01011100 : OUT <= 2;  //217 / 92 = 2
    16'b11011001_01011101 : OUT <= 2;  //217 / 93 = 2
    16'b11011001_01011110 : OUT <= 2;  //217 / 94 = 2
    16'b11011001_01011111 : OUT <= 2;  //217 / 95 = 2
    16'b11011001_01100000 : OUT <= 2;  //217 / 96 = 2
    16'b11011001_01100001 : OUT <= 2;  //217 / 97 = 2
    16'b11011001_01100010 : OUT <= 2;  //217 / 98 = 2
    16'b11011001_01100011 : OUT <= 2;  //217 / 99 = 2
    16'b11011001_01100100 : OUT <= 2;  //217 / 100 = 2
    16'b11011001_01100101 : OUT <= 2;  //217 / 101 = 2
    16'b11011001_01100110 : OUT <= 2;  //217 / 102 = 2
    16'b11011001_01100111 : OUT <= 2;  //217 / 103 = 2
    16'b11011001_01101000 : OUT <= 2;  //217 / 104 = 2
    16'b11011001_01101001 : OUT <= 2;  //217 / 105 = 2
    16'b11011001_01101010 : OUT <= 2;  //217 / 106 = 2
    16'b11011001_01101011 : OUT <= 2;  //217 / 107 = 2
    16'b11011001_01101100 : OUT <= 2;  //217 / 108 = 2
    16'b11011001_01101101 : OUT <= 1;  //217 / 109 = 1
    16'b11011001_01101110 : OUT <= 1;  //217 / 110 = 1
    16'b11011001_01101111 : OUT <= 1;  //217 / 111 = 1
    16'b11011001_01110000 : OUT <= 1;  //217 / 112 = 1
    16'b11011001_01110001 : OUT <= 1;  //217 / 113 = 1
    16'b11011001_01110010 : OUT <= 1;  //217 / 114 = 1
    16'b11011001_01110011 : OUT <= 1;  //217 / 115 = 1
    16'b11011001_01110100 : OUT <= 1;  //217 / 116 = 1
    16'b11011001_01110101 : OUT <= 1;  //217 / 117 = 1
    16'b11011001_01110110 : OUT <= 1;  //217 / 118 = 1
    16'b11011001_01110111 : OUT <= 1;  //217 / 119 = 1
    16'b11011001_01111000 : OUT <= 1;  //217 / 120 = 1
    16'b11011001_01111001 : OUT <= 1;  //217 / 121 = 1
    16'b11011001_01111010 : OUT <= 1;  //217 / 122 = 1
    16'b11011001_01111011 : OUT <= 1;  //217 / 123 = 1
    16'b11011001_01111100 : OUT <= 1;  //217 / 124 = 1
    16'b11011001_01111101 : OUT <= 1;  //217 / 125 = 1
    16'b11011001_01111110 : OUT <= 1;  //217 / 126 = 1
    16'b11011001_01111111 : OUT <= 1;  //217 / 127 = 1
    16'b11011001_10000000 : OUT <= 1;  //217 / 128 = 1
    16'b11011001_10000001 : OUT <= 1;  //217 / 129 = 1
    16'b11011001_10000010 : OUT <= 1;  //217 / 130 = 1
    16'b11011001_10000011 : OUT <= 1;  //217 / 131 = 1
    16'b11011001_10000100 : OUT <= 1;  //217 / 132 = 1
    16'b11011001_10000101 : OUT <= 1;  //217 / 133 = 1
    16'b11011001_10000110 : OUT <= 1;  //217 / 134 = 1
    16'b11011001_10000111 : OUT <= 1;  //217 / 135 = 1
    16'b11011001_10001000 : OUT <= 1;  //217 / 136 = 1
    16'b11011001_10001001 : OUT <= 1;  //217 / 137 = 1
    16'b11011001_10001010 : OUT <= 1;  //217 / 138 = 1
    16'b11011001_10001011 : OUT <= 1;  //217 / 139 = 1
    16'b11011001_10001100 : OUT <= 1;  //217 / 140 = 1
    16'b11011001_10001101 : OUT <= 1;  //217 / 141 = 1
    16'b11011001_10001110 : OUT <= 1;  //217 / 142 = 1
    16'b11011001_10001111 : OUT <= 1;  //217 / 143 = 1
    16'b11011001_10010000 : OUT <= 1;  //217 / 144 = 1
    16'b11011001_10010001 : OUT <= 1;  //217 / 145 = 1
    16'b11011001_10010010 : OUT <= 1;  //217 / 146 = 1
    16'b11011001_10010011 : OUT <= 1;  //217 / 147 = 1
    16'b11011001_10010100 : OUT <= 1;  //217 / 148 = 1
    16'b11011001_10010101 : OUT <= 1;  //217 / 149 = 1
    16'b11011001_10010110 : OUT <= 1;  //217 / 150 = 1
    16'b11011001_10010111 : OUT <= 1;  //217 / 151 = 1
    16'b11011001_10011000 : OUT <= 1;  //217 / 152 = 1
    16'b11011001_10011001 : OUT <= 1;  //217 / 153 = 1
    16'b11011001_10011010 : OUT <= 1;  //217 / 154 = 1
    16'b11011001_10011011 : OUT <= 1;  //217 / 155 = 1
    16'b11011001_10011100 : OUT <= 1;  //217 / 156 = 1
    16'b11011001_10011101 : OUT <= 1;  //217 / 157 = 1
    16'b11011001_10011110 : OUT <= 1;  //217 / 158 = 1
    16'b11011001_10011111 : OUT <= 1;  //217 / 159 = 1
    16'b11011001_10100000 : OUT <= 1;  //217 / 160 = 1
    16'b11011001_10100001 : OUT <= 1;  //217 / 161 = 1
    16'b11011001_10100010 : OUT <= 1;  //217 / 162 = 1
    16'b11011001_10100011 : OUT <= 1;  //217 / 163 = 1
    16'b11011001_10100100 : OUT <= 1;  //217 / 164 = 1
    16'b11011001_10100101 : OUT <= 1;  //217 / 165 = 1
    16'b11011001_10100110 : OUT <= 1;  //217 / 166 = 1
    16'b11011001_10100111 : OUT <= 1;  //217 / 167 = 1
    16'b11011001_10101000 : OUT <= 1;  //217 / 168 = 1
    16'b11011001_10101001 : OUT <= 1;  //217 / 169 = 1
    16'b11011001_10101010 : OUT <= 1;  //217 / 170 = 1
    16'b11011001_10101011 : OUT <= 1;  //217 / 171 = 1
    16'b11011001_10101100 : OUT <= 1;  //217 / 172 = 1
    16'b11011001_10101101 : OUT <= 1;  //217 / 173 = 1
    16'b11011001_10101110 : OUT <= 1;  //217 / 174 = 1
    16'b11011001_10101111 : OUT <= 1;  //217 / 175 = 1
    16'b11011001_10110000 : OUT <= 1;  //217 / 176 = 1
    16'b11011001_10110001 : OUT <= 1;  //217 / 177 = 1
    16'b11011001_10110010 : OUT <= 1;  //217 / 178 = 1
    16'b11011001_10110011 : OUT <= 1;  //217 / 179 = 1
    16'b11011001_10110100 : OUT <= 1;  //217 / 180 = 1
    16'b11011001_10110101 : OUT <= 1;  //217 / 181 = 1
    16'b11011001_10110110 : OUT <= 1;  //217 / 182 = 1
    16'b11011001_10110111 : OUT <= 1;  //217 / 183 = 1
    16'b11011001_10111000 : OUT <= 1;  //217 / 184 = 1
    16'b11011001_10111001 : OUT <= 1;  //217 / 185 = 1
    16'b11011001_10111010 : OUT <= 1;  //217 / 186 = 1
    16'b11011001_10111011 : OUT <= 1;  //217 / 187 = 1
    16'b11011001_10111100 : OUT <= 1;  //217 / 188 = 1
    16'b11011001_10111101 : OUT <= 1;  //217 / 189 = 1
    16'b11011001_10111110 : OUT <= 1;  //217 / 190 = 1
    16'b11011001_10111111 : OUT <= 1;  //217 / 191 = 1
    16'b11011001_11000000 : OUT <= 1;  //217 / 192 = 1
    16'b11011001_11000001 : OUT <= 1;  //217 / 193 = 1
    16'b11011001_11000010 : OUT <= 1;  //217 / 194 = 1
    16'b11011001_11000011 : OUT <= 1;  //217 / 195 = 1
    16'b11011001_11000100 : OUT <= 1;  //217 / 196 = 1
    16'b11011001_11000101 : OUT <= 1;  //217 / 197 = 1
    16'b11011001_11000110 : OUT <= 1;  //217 / 198 = 1
    16'b11011001_11000111 : OUT <= 1;  //217 / 199 = 1
    16'b11011001_11001000 : OUT <= 1;  //217 / 200 = 1
    16'b11011001_11001001 : OUT <= 1;  //217 / 201 = 1
    16'b11011001_11001010 : OUT <= 1;  //217 / 202 = 1
    16'b11011001_11001011 : OUT <= 1;  //217 / 203 = 1
    16'b11011001_11001100 : OUT <= 1;  //217 / 204 = 1
    16'b11011001_11001101 : OUT <= 1;  //217 / 205 = 1
    16'b11011001_11001110 : OUT <= 1;  //217 / 206 = 1
    16'b11011001_11001111 : OUT <= 1;  //217 / 207 = 1
    16'b11011001_11010000 : OUT <= 1;  //217 / 208 = 1
    16'b11011001_11010001 : OUT <= 1;  //217 / 209 = 1
    16'b11011001_11010010 : OUT <= 1;  //217 / 210 = 1
    16'b11011001_11010011 : OUT <= 1;  //217 / 211 = 1
    16'b11011001_11010100 : OUT <= 1;  //217 / 212 = 1
    16'b11011001_11010101 : OUT <= 1;  //217 / 213 = 1
    16'b11011001_11010110 : OUT <= 1;  //217 / 214 = 1
    16'b11011001_11010111 : OUT <= 1;  //217 / 215 = 1
    16'b11011001_11011000 : OUT <= 1;  //217 / 216 = 1
    16'b11011001_11011001 : OUT <= 1;  //217 / 217 = 1
    16'b11011001_11011010 : OUT <= 0;  //217 / 218 = 0
    16'b11011001_11011011 : OUT <= 0;  //217 / 219 = 0
    16'b11011001_11011100 : OUT <= 0;  //217 / 220 = 0
    16'b11011001_11011101 : OUT <= 0;  //217 / 221 = 0
    16'b11011001_11011110 : OUT <= 0;  //217 / 222 = 0
    16'b11011001_11011111 : OUT <= 0;  //217 / 223 = 0
    16'b11011001_11100000 : OUT <= 0;  //217 / 224 = 0
    16'b11011001_11100001 : OUT <= 0;  //217 / 225 = 0
    16'b11011001_11100010 : OUT <= 0;  //217 / 226 = 0
    16'b11011001_11100011 : OUT <= 0;  //217 / 227 = 0
    16'b11011001_11100100 : OUT <= 0;  //217 / 228 = 0
    16'b11011001_11100101 : OUT <= 0;  //217 / 229 = 0
    16'b11011001_11100110 : OUT <= 0;  //217 / 230 = 0
    16'b11011001_11100111 : OUT <= 0;  //217 / 231 = 0
    16'b11011001_11101000 : OUT <= 0;  //217 / 232 = 0
    16'b11011001_11101001 : OUT <= 0;  //217 / 233 = 0
    16'b11011001_11101010 : OUT <= 0;  //217 / 234 = 0
    16'b11011001_11101011 : OUT <= 0;  //217 / 235 = 0
    16'b11011001_11101100 : OUT <= 0;  //217 / 236 = 0
    16'b11011001_11101101 : OUT <= 0;  //217 / 237 = 0
    16'b11011001_11101110 : OUT <= 0;  //217 / 238 = 0
    16'b11011001_11101111 : OUT <= 0;  //217 / 239 = 0
    16'b11011001_11110000 : OUT <= 0;  //217 / 240 = 0
    16'b11011001_11110001 : OUT <= 0;  //217 / 241 = 0
    16'b11011001_11110010 : OUT <= 0;  //217 / 242 = 0
    16'b11011001_11110011 : OUT <= 0;  //217 / 243 = 0
    16'b11011001_11110100 : OUT <= 0;  //217 / 244 = 0
    16'b11011001_11110101 : OUT <= 0;  //217 / 245 = 0
    16'b11011001_11110110 : OUT <= 0;  //217 / 246 = 0
    16'b11011001_11110111 : OUT <= 0;  //217 / 247 = 0
    16'b11011001_11111000 : OUT <= 0;  //217 / 248 = 0
    16'b11011001_11111001 : OUT <= 0;  //217 / 249 = 0
    16'b11011001_11111010 : OUT <= 0;  //217 / 250 = 0
    16'b11011001_11111011 : OUT <= 0;  //217 / 251 = 0
    16'b11011001_11111100 : OUT <= 0;  //217 / 252 = 0
    16'b11011001_11111101 : OUT <= 0;  //217 / 253 = 0
    16'b11011001_11111110 : OUT <= 0;  //217 / 254 = 0
    16'b11011001_11111111 : OUT <= 0;  //217 / 255 = 0
    16'b11011010_00000000 : OUT <= 0;  //218 / 0 = 0
    16'b11011010_00000001 : OUT <= 218;  //218 / 1 = 218
    16'b11011010_00000010 : OUT <= 109;  //218 / 2 = 109
    16'b11011010_00000011 : OUT <= 72;  //218 / 3 = 72
    16'b11011010_00000100 : OUT <= 54;  //218 / 4 = 54
    16'b11011010_00000101 : OUT <= 43;  //218 / 5 = 43
    16'b11011010_00000110 : OUT <= 36;  //218 / 6 = 36
    16'b11011010_00000111 : OUT <= 31;  //218 / 7 = 31
    16'b11011010_00001000 : OUT <= 27;  //218 / 8 = 27
    16'b11011010_00001001 : OUT <= 24;  //218 / 9 = 24
    16'b11011010_00001010 : OUT <= 21;  //218 / 10 = 21
    16'b11011010_00001011 : OUT <= 19;  //218 / 11 = 19
    16'b11011010_00001100 : OUT <= 18;  //218 / 12 = 18
    16'b11011010_00001101 : OUT <= 16;  //218 / 13 = 16
    16'b11011010_00001110 : OUT <= 15;  //218 / 14 = 15
    16'b11011010_00001111 : OUT <= 14;  //218 / 15 = 14
    16'b11011010_00010000 : OUT <= 13;  //218 / 16 = 13
    16'b11011010_00010001 : OUT <= 12;  //218 / 17 = 12
    16'b11011010_00010010 : OUT <= 12;  //218 / 18 = 12
    16'b11011010_00010011 : OUT <= 11;  //218 / 19 = 11
    16'b11011010_00010100 : OUT <= 10;  //218 / 20 = 10
    16'b11011010_00010101 : OUT <= 10;  //218 / 21 = 10
    16'b11011010_00010110 : OUT <= 9;  //218 / 22 = 9
    16'b11011010_00010111 : OUT <= 9;  //218 / 23 = 9
    16'b11011010_00011000 : OUT <= 9;  //218 / 24 = 9
    16'b11011010_00011001 : OUT <= 8;  //218 / 25 = 8
    16'b11011010_00011010 : OUT <= 8;  //218 / 26 = 8
    16'b11011010_00011011 : OUT <= 8;  //218 / 27 = 8
    16'b11011010_00011100 : OUT <= 7;  //218 / 28 = 7
    16'b11011010_00011101 : OUT <= 7;  //218 / 29 = 7
    16'b11011010_00011110 : OUT <= 7;  //218 / 30 = 7
    16'b11011010_00011111 : OUT <= 7;  //218 / 31 = 7
    16'b11011010_00100000 : OUT <= 6;  //218 / 32 = 6
    16'b11011010_00100001 : OUT <= 6;  //218 / 33 = 6
    16'b11011010_00100010 : OUT <= 6;  //218 / 34 = 6
    16'b11011010_00100011 : OUT <= 6;  //218 / 35 = 6
    16'b11011010_00100100 : OUT <= 6;  //218 / 36 = 6
    16'b11011010_00100101 : OUT <= 5;  //218 / 37 = 5
    16'b11011010_00100110 : OUT <= 5;  //218 / 38 = 5
    16'b11011010_00100111 : OUT <= 5;  //218 / 39 = 5
    16'b11011010_00101000 : OUT <= 5;  //218 / 40 = 5
    16'b11011010_00101001 : OUT <= 5;  //218 / 41 = 5
    16'b11011010_00101010 : OUT <= 5;  //218 / 42 = 5
    16'b11011010_00101011 : OUT <= 5;  //218 / 43 = 5
    16'b11011010_00101100 : OUT <= 4;  //218 / 44 = 4
    16'b11011010_00101101 : OUT <= 4;  //218 / 45 = 4
    16'b11011010_00101110 : OUT <= 4;  //218 / 46 = 4
    16'b11011010_00101111 : OUT <= 4;  //218 / 47 = 4
    16'b11011010_00110000 : OUT <= 4;  //218 / 48 = 4
    16'b11011010_00110001 : OUT <= 4;  //218 / 49 = 4
    16'b11011010_00110010 : OUT <= 4;  //218 / 50 = 4
    16'b11011010_00110011 : OUT <= 4;  //218 / 51 = 4
    16'b11011010_00110100 : OUT <= 4;  //218 / 52 = 4
    16'b11011010_00110101 : OUT <= 4;  //218 / 53 = 4
    16'b11011010_00110110 : OUT <= 4;  //218 / 54 = 4
    16'b11011010_00110111 : OUT <= 3;  //218 / 55 = 3
    16'b11011010_00111000 : OUT <= 3;  //218 / 56 = 3
    16'b11011010_00111001 : OUT <= 3;  //218 / 57 = 3
    16'b11011010_00111010 : OUT <= 3;  //218 / 58 = 3
    16'b11011010_00111011 : OUT <= 3;  //218 / 59 = 3
    16'b11011010_00111100 : OUT <= 3;  //218 / 60 = 3
    16'b11011010_00111101 : OUT <= 3;  //218 / 61 = 3
    16'b11011010_00111110 : OUT <= 3;  //218 / 62 = 3
    16'b11011010_00111111 : OUT <= 3;  //218 / 63 = 3
    16'b11011010_01000000 : OUT <= 3;  //218 / 64 = 3
    16'b11011010_01000001 : OUT <= 3;  //218 / 65 = 3
    16'b11011010_01000010 : OUT <= 3;  //218 / 66 = 3
    16'b11011010_01000011 : OUT <= 3;  //218 / 67 = 3
    16'b11011010_01000100 : OUT <= 3;  //218 / 68 = 3
    16'b11011010_01000101 : OUT <= 3;  //218 / 69 = 3
    16'b11011010_01000110 : OUT <= 3;  //218 / 70 = 3
    16'b11011010_01000111 : OUT <= 3;  //218 / 71 = 3
    16'b11011010_01001000 : OUT <= 3;  //218 / 72 = 3
    16'b11011010_01001001 : OUT <= 2;  //218 / 73 = 2
    16'b11011010_01001010 : OUT <= 2;  //218 / 74 = 2
    16'b11011010_01001011 : OUT <= 2;  //218 / 75 = 2
    16'b11011010_01001100 : OUT <= 2;  //218 / 76 = 2
    16'b11011010_01001101 : OUT <= 2;  //218 / 77 = 2
    16'b11011010_01001110 : OUT <= 2;  //218 / 78 = 2
    16'b11011010_01001111 : OUT <= 2;  //218 / 79 = 2
    16'b11011010_01010000 : OUT <= 2;  //218 / 80 = 2
    16'b11011010_01010001 : OUT <= 2;  //218 / 81 = 2
    16'b11011010_01010010 : OUT <= 2;  //218 / 82 = 2
    16'b11011010_01010011 : OUT <= 2;  //218 / 83 = 2
    16'b11011010_01010100 : OUT <= 2;  //218 / 84 = 2
    16'b11011010_01010101 : OUT <= 2;  //218 / 85 = 2
    16'b11011010_01010110 : OUT <= 2;  //218 / 86 = 2
    16'b11011010_01010111 : OUT <= 2;  //218 / 87 = 2
    16'b11011010_01011000 : OUT <= 2;  //218 / 88 = 2
    16'b11011010_01011001 : OUT <= 2;  //218 / 89 = 2
    16'b11011010_01011010 : OUT <= 2;  //218 / 90 = 2
    16'b11011010_01011011 : OUT <= 2;  //218 / 91 = 2
    16'b11011010_01011100 : OUT <= 2;  //218 / 92 = 2
    16'b11011010_01011101 : OUT <= 2;  //218 / 93 = 2
    16'b11011010_01011110 : OUT <= 2;  //218 / 94 = 2
    16'b11011010_01011111 : OUT <= 2;  //218 / 95 = 2
    16'b11011010_01100000 : OUT <= 2;  //218 / 96 = 2
    16'b11011010_01100001 : OUT <= 2;  //218 / 97 = 2
    16'b11011010_01100010 : OUT <= 2;  //218 / 98 = 2
    16'b11011010_01100011 : OUT <= 2;  //218 / 99 = 2
    16'b11011010_01100100 : OUT <= 2;  //218 / 100 = 2
    16'b11011010_01100101 : OUT <= 2;  //218 / 101 = 2
    16'b11011010_01100110 : OUT <= 2;  //218 / 102 = 2
    16'b11011010_01100111 : OUT <= 2;  //218 / 103 = 2
    16'b11011010_01101000 : OUT <= 2;  //218 / 104 = 2
    16'b11011010_01101001 : OUT <= 2;  //218 / 105 = 2
    16'b11011010_01101010 : OUT <= 2;  //218 / 106 = 2
    16'b11011010_01101011 : OUT <= 2;  //218 / 107 = 2
    16'b11011010_01101100 : OUT <= 2;  //218 / 108 = 2
    16'b11011010_01101101 : OUT <= 2;  //218 / 109 = 2
    16'b11011010_01101110 : OUT <= 1;  //218 / 110 = 1
    16'b11011010_01101111 : OUT <= 1;  //218 / 111 = 1
    16'b11011010_01110000 : OUT <= 1;  //218 / 112 = 1
    16'b11011010_01110001 : OUT <= 1;  //218 / 113 = 1
    16'b11011010_01110010 : OUT <= 1;  //218 / 114 = 1
    16'b11011010_01110011 : OUT <= 1;  //218 / 115 = 1
    16'b11011010_01110100 : OUT <= 1;  //218 / 116 = 1
    16'b11011010_01110101 : OUT <= 1;  //218 / 117 = 1
    16'b11011010_01110110 : OUT <= 1;  //218 / 118 = 1
    16'b11011010_01110111 : OUT <= 1;  //218 / 119 = 1
    16'b11011010_01111000 : OUT <= 1;  //218 / 120 = 1
    16'b11011010_01111001 : OUT <= 1;  //218 / 121 = 1
    16'b11011010_01111010 : OUT <= 1;  //218 / 122 = 1
    16'b11011010_01111011 : OUT <= 1;  //218 / 123 = 1
    16'b11011010_01111100 : OUT <= 1;  //218 / 124 = 1
    16'b11011010_01111101 : OUT <= 1;  //218 / 125 = 1
    16'b11011010_01111110 : OUT <= 1;  //218 / 126 = 1
    16'b11011010_01111111 : OUT <= 1;  //218 / 127 = 1
    16'b11011010_10000000 : OUT <= 1;  //218 / 128 = 1
    16'b11011010_10000001 : OUT <= 1;  //218 / 129 = 1
    16'b11011010_10000010 : OUT <= 1;  //218 / 130 = 1
    16'b11011010_10000011 : OUT <= 1;  //218 / 131 = 1
    16'b11011010_10000100 : OUT <= 1;  //218 / 132 = 1
    16'b11011010_10000101 : OUT <= 1;  //218 / 133 = 1
    16'b11011010_10000110 : OUT <= 1;  //218 / 134 = 1
    16'b11011010_10000111 : OUT <= 1;  //218 / 135 = 1
    16'b11011010_10001000 : OUT <= 1;  //218 / 136 = 1
    16'b11011010_10001001 : OUT <= 1;  //218 / 137 = 1
    16'b11011010_10001010 : OUT <= 1;  //218 / 138 = 1
    16'b11011010_10001011 : OUT <= 1;  //218 / 139 = 1
    16'b11011010_10001100 : OUT <= 1;  //218 / 140 = 1
    16'b11011010_10001101 : OUT <= 1;  //218 / 141 = 1
    16'b11011010_10001110 : OUT <= 1;  //218 / 142 = 1
    16'b11011010_10001111 : OUT <= 1;  //218 / 143 = 1
    16'b11011010_10010000 : OUT <= 1;  //218 / 144 = 1
    16'b11011010_10010001 : OUT <= 1;  //218 / 145 = 1
    16'b11011010_10010010 : OUT <= 1;  //218 / 146 = 1
    16'b11011010_10010011 : OUT <= 1;  //218 / 147 = 1
    16'b11011010_10010100 : OUT <= 1;  //218 / 148 = 1
    16'b11011010_10010101 : OUT <= 1;  //218 / 149 = 1
    16'b11011010_10010110 : OUT <= 1;  //218 / 150 = 1
    16'b11011010_10010111 : OUT <= 1;  //218 / 151 = 1
    16'b11011010_10011000 : OUT <= 1;  //218 / 152 = 1
    16'b11011010_10011001 : OUT <= 1;  //218 / 153 = 1
    16'b11011010_10011010 : OUT <= 1;  //218 / 154 = 1
    16'b11011010_10011011 : OUT <= 1;  //218 / 155 = 1
    16'b11011010_10011100 : OUT <= 1;  //218 / 156 = 1
    16'b11011010_10011101 : OUT <= 1;  //218 / 157 = 1
    16'b11011010_10011110 : OUT <= 1;  //218 / 158 = 1
    16'b11011010_10011111 : OUT <= 1;  //218 / 159 = 1
    16'b11011010_10100000 : OUT <= 1;  //218 / 160 = 1
    16'b11011010_10100001 : OUT <= 1;  //218 / 161 = 1
    16'b11011010_10100010 : OUT <= 1;  //218 / 162 = 1
    16'b11011010_10100011 : OUT <= 1;  //218 / 163 = 1
    16'b11011010_10100100 : OUT <= 1;  //218 / 164 = 1
    16'b11011010_10100101 : OUT <= 1;  //218 / 165 = 1
    16'b11011010_10100110 : OUT <= 1;  //218 / 166 = 1
    16'b11011010_10100111 : OUT <= 1;  //218 / 167 = 1
    16'b11011010_10101000 : OUT <= 1;  //218 / 168 = 1
    16'b11011010_10101001 : OUT <= 1;  //218 / 169 = 1
    16'b11011010_10101010 : OUT <= 1;  //218 / 170 = 1
    16'b11011010_10101011 : OUT <= 1;  //218 / 171 = 1
    16'b11011010_10101100 : OUT <= 1;  //218 / 172 = 1
    16'b11011010_10101101 : OUT <= 1;  //218 / 173 = 1
    16'b11011010_10101110 : OUT <= 1;  //218 / 174 = 1
    16'b11011010_10101111 : OUT <= 1;  //218 / 175 = 1
    16'b11011010_10110000 : OUT <= 1;  //218 / 176 = 1
    16'b11011010_10110001 : OUT <= 1;  //218 / 177 = 1
    16'b11011010_10110010 : OUT <= 1;  //218 / 178 = 1
    16'b11011010_10110011 : OUT <= 1;  //218 / 179 = 1
    16'b11011010_10110100 : OUT <= 1;  //218 / 180 = 1
    16'b11011010_10110101 : OUT <= 1;  //218 / 181 = 1
    16'b11011010_10110110 : OUT <= 1;  //218 / 182 = 1
    16'b11011010_10110111 : OUT <= 1;  //218 / 183 = 1
    16'b11011010_10111000 : OUT <= 1;  //218 / 184 = 1
    16'b11011010_10111001 : OUT <= 1;  //218 / 185 = 1
    16'b11011010_10111010 : OUT <= 1;  //218 / 186 = 1
    16'b11011010_10111011 : OUT <= 1;  //218 / 187 = 1
    16'b11011010_10111100 : OUT <= 1;  //218 / 188 = 1
    16'b11011010_10111101 : OUT <= 1;  //218 / 189 = 1
    16'b11011010_10111110 : OUT <= 1;  //218 / 190 = 1
    16'b11011010_10111111 : OUT <= 1;  //218 / 191 = 1
    16'b11011010_11000000 : OUT <= 1;  //218 / 192 = 1
    16'b11011010_11000001 : OUT <= 1;  //218 / 193 = 1
    16'b11011010_11000010 : OUT <= 1;  //218 / 194 = 1
    16'b11011010_11000011 : OUT <= 1;  //218 / 195 = 1
    16'b11011010_11000100 : OUT <= 1;  //218 / 196 = 1
    16'b11011010_11000101 : OUT <= 1;  //218 / 197 = 1
    16'b11011010_11000110 : OUT <= 1;  //218 / 198 = 1
    16'b11011010_11000111 : OUT <= 1;  //218 / 199 = 1
    16'b11011010_11001000 : OUT <= 1;  //218 / 200 = 1
    16'b11011010_11001001 : OUT <= 1;  //218 / 201 = 1
    16'b11011010_11001010 : OUT <= 1;  //218 / 202 = 1
    16'b11011010_11001011 : OUT <= 1;  //218 / 203 = 1
    16'b11011010_11001100 : OUT <= 1;  //218 / 204 = 1
    16'b11011010_11001101 : OUT <= 1;  //218 / 205 = 1
    16'b11011010_11001110 : OUT <= 1;  //218 / 206 = 1
    16'b11011010_11001111 : OUT <= 1;  //218 / 207 = 1
    16'b11011010_11010000 : OUT <= 1;  //218 / 208 = 1
    16'b11011010_11010001 : OUT <= 1;  //218 / 209 = 1
    16'b11011010_11010010 : OUT <= 1;  //218 / 210 = 1
    16'b11011010_11010011 : OUT <= 1;  //218 / 211 = 1
    16'b11011010_11010100 : OUT <= 1;  //218 / 212 = 1
    16'b11011010_11010101 : OUT <= 1;  //218 / 213 = 1
    16'b11011010_11010110 : OUT <= 1;  //218 / 214 = 1
    16'b11011010_11010111 : OUT <= 1;  //218 / 215 = 1
    16'b11011010_11011000 : OUT <= 1;  //218 / 216 = 1
    16'b11011010_11011001 : OUT <= 1;  //218 / 217 = 1
    16'b11011010_11011010 : OUT <= 1;  //218 / 218 = 1
    16'b11011010_11011011 : OUT <= 0;  //218 / 219 = 0
    16'b11011010_11011100 : OUT <= 0;  //218 / 220 = 0
    16'b11011010_11011101 : OUT <= 0;  //218 / 221 = 0
    16'b11011010_11011110 : OUT <= 0;  //218 / 222 = 0
    16'b11011010_11011111 : OUT <= 0;  //218 / 223 = 0
    16'b11011010_11100000 : OUT <= 0;  //218 / 224 = 0
    16'b11011010_11100001 : OUT <= 0;  //218 / 225 = 0
    16'b11011010_11100010 : OUT <= 0;  //218 / 226 = 0
    16'b11011010_11100011 : OUT <= 0;  //218 / 227 = 0
    16'b11011010_11100100 : OUT <= 0;  //218 / 228 = 0
    16'b11011010_11100101 : OUT <= 0;  //218 / 229 = 0
    16'b11011010_11100110 : OUT <= 0;  //218 / 230 = 0
    16'b11011010_11100111 : OUT <= 0;  //218 / 231 = 0
    16'b11011010_11101000 : OUT <= 0;  //218 / 232 = 0
    16'b11011010_11101001 : OUT <= 0;  //218 / 233 = 0
    16'b11011010_11101010 : OUT <= 0;  //218 / 234 = 0
    16'b11011010_11101011 : OUT <= 0;  //218 / 235 = 0
    16'b11011010_11101100 : OUT <= 0;  //218 / 236 = 0
    16'b11011010_11101101 : OUT <= 0;  //218 / 237 = 0
    16'b11011010_11101110 : OUT <= 0;  //218 / 238 = 0
    16'b11011010_11101111 : OUT <= 0;  //218 / 239 = 0
    16'b11011010_11110000 : OUT <= 0;  //218 / 240 = 0
    16'b11011010_11110001 : OUT <= 0;  //218 / 241 = 0
    16'b11011010_11110010 : OUT <= 0;  //218 / 242 = 0
    16'b11011010_11110011 : OUT <= 0;  //218 / 243 = 0
    16'b11011010_11110100 : OUT <= 0;  //218 / 244 = 0
    16'b11011010_11110101 : OUT <= 0;  //218 / 245 = 0
    16'b11011010_11110110 : OUT <= 0;  //218 / 246 = 0
    16'b11011010_11110111 : OUT <= 0;  //218 / 247 = 0
    16'b11011010_11111000 : OUT <= 0;  //218 / 248 = 0
    16'b11011010_11111001 : OUT <= 0;  //218 / 249 = 0
    16'b11011010_11111010 : OUT <= 0;  //218 / 250 = 0
    16'b11011010_11111011 : OUT <= 0;  //218 / 251 = 0
    16'b11011010_11111100 : OUT <= 0;  //218 / 252 = 0
    16'b11011010_11111101 : OUT <= 0;  //218 / 253 = 0
    16'b11011010_11111110 : OUT <= 0;  //218 / 254 = 0
    16'b11011010_11111111 : OUT <= 0;  //218 / 255 = 0
    16'b11011011_00000000 : OUT <= 0;  //219 / 0 = 0
    16'b11011011_00000001 : OUT <= 219;  //219 / 1 = 219
    16'b11011011_00000010 : OUT <= 109;  //219 / 2 = 109
    16'b11011011_00000011 : OUT <= 73;  //219 / 3 = 73
    16'b11011011_00000100 : OUT <= 54;  //219 / 4 = 54
    16'b11011011_00000101 : OUT <= 43;  //219 / 5 = 43
    16'b11011011_00000110 : OUT <= 36;  //219 / 6 = 36
    16'b11011011_00000111 : OUT <= 31;  //219 / 7 = 31
    16'b11011011_00001000 : OUT <= 27;  //219 / 8 = 27
    16'b11011011_00001001 : OUT <= 24;  //219 / 9 = 24
    16'b11011011_00001010 : OUT <= 21;  //219 / 10 = 21
    16'b11011011_00001011 : OUT <= 19;  //219 / 11 = 19
    16'b11011011_00001100 : OUT <= 18;  //219 / 12 = 18
    16'b11011011_00001101 : OUT <= 16;  //219 / 13 = 16
    16'b11011011_00001110 : OUT <= 15;  //219 / 14 = 15
    16'b11011011_00001111 : OUT <= 14;  //219 / 15 = 14
    16'b11011011_00010000 : OUT <= 13;  //219 / 16 = 13
    16'b11011011_00010001 : OUT <= 12;  //219 / 17 = 12
    16'b11011011_00010010 : OUT <= 12;  //219 / 18 = 12
    16'b11011011_00010011 : OUT <= 11;  //219 / 19 = 11
    16'b11011011_00010100 : OUT <= 10;  //219 / 20 = 10
    16'b11011011_00010101 : OUT <= 10;  //219 / 21 = 10
    16'b11011011_00010110 : OUT <= 9;  //219 / 22 = 9
    16'b11011011_00010111 : OUT <= 9;  //219 / 23 = 9
    16'b11011011_00011000 : OUT <= 9;  //219 / 24 = 9
    16'b11011011_00011001 : OUT <= 8;  //219 / 25 = 8
    16'b11011011_00011010 : OUT <= 8;  //219 / 26 = 8
    16'b11011011_00011011 : OUT <= 8;  //219 / 27 = 8
    16'b11011011_00011100 : OUT <= 7;  //219 / 28 = 7
    16'b11011011_00011101 : OUT <= 7;  //219 / 29 = 7
    16'b11011011_00011110 : OUT <= 7;  //219 / 30 = 7
    16'b11011011_00011111 : OUT <= 7;  //219 / 31 = 7
    16'b11011011_00100000 : OUT <= 6;  //219 / 32 = 6
    16'b11011011_00100001 : OUT <= 6;  //219 / 33 = 6
    16'b11011011_00100010 : OUT <= 6;  //219 / 34 = 6
    16'b11011011_00100011 : OUT <= 6;  //219 / 35 = 6
    16'b11011011_00100100 : OUT <= 6;  //219 / 36 = 6
    16'b11011011_00100101 : OUT <= 5;  //219 / 37 = 5
    16'b11011011_00100110 : OUT <= 5;  //219 / 38 = 5
    16'b11011011_00100111 : OUT <= 5;  //219 / 39 = 5
    16'b11011011_00101000 : OUT <= 5;  //219 / 40 = 5
    16'b11011011_00101001 : OUT <= 5;  //219 / 41 = 5
    16'b11011011_00101010 : OUT <= 5;  //219 / 42 = 5
    16'b11011011_00101011 : OUT <= 5;  //219 / 43 = 5
    16'b11011011_00101100 : OUT <= 4;  //219 / 44 = 4
    16'b11011011_00101101 : OUT <= 4;  //219 / 45 = 4
    16'b11011011_00101110 : OUT <= 4;  //219 / 46 = 4
    16'b11011011_00101111 : OUT <= 4;  //219 / 47 = 4
    16'b11011011_00110000 : OUT <= 4;  //219 / 48 = 4
    16'b11011011_00110001 : OUT <= 4;  //219 / 49 = 4
    16'b11011011_00110010 : OUT <= 4;  //219 / 50 = 4
    16'b11011011_00110011 : OUT <= 4;  //219 / 51 = 4
    16'b11011011_00110100 : OUT <= 4;  //219 / 52 = 4
    16'b11011011_00110101 : OUT <= 4;  //219 / 53 = 4
    16'b11011011_00110110 : OUT <= 4;  //219 / 54 = 4
    16'b11011011_00110111 : OUT <= 3;  //219 / 55 = 3
    16'b11011011_00111000 : OUT <= 3;  //219 / 56 = 3
    16'b11011011_00111001 : OUT <= 3;  //219 / 57 = 3
    16'b11011011_00111010 : OUT <= 3;  //219 / 58 = 3
    16'b11011011_00111011 : OUT <= 3;  //219 / 59 = 3
    16'b11011011_00111100 : OUT <= 3;  //219 / 60 = 3
    16'b11011011_00111101 : OUT <= 3;  //219 / 61 = 3
    16'b11011011_00111110 : OUT <= 3;  //219 / 62 = 3
    16'b11011011_00111111 : OUT <= 3;  //219 / 63 = 3
    16'b11011011_01000000 : OUT <= 3;  //219 / 64 = 3
    16'b11011011_01000001 : OUT <= 3;  //219 / 65 = 3
    16'b11011011_01000010 : OUT <= 3;  //219 / 66 = 3
    16'b11011011_01000011 : OUT <= 3;  //219 / 67 = 3
    16'b11011011_01000100 : OUT <= 3;  //219 / 68 = 3
    16'b11011011_01000101 : OUT <= 3;  //219 / 69 = 3
    16'b11011011_01000110 : OUT <= 3;  //219 / 70 = 3
    16'b11011011_01000111 : OUT <= 3;  //219 / 71 = 3
    16'b11011011_01001000 : OUT <= 3;  //219 / 72 = 3
    16'b11011011_01001001 : OUT <= 3;  //219 / 73 = 3
    16'b11011011_01001010 : OUT <= 2;  //219 / 74 = 2
    16'b11011011_01001011 : OUT <= 2;  //219 / 75 = 2
    16'b11011011_01001100 : OUT <= 2;  //219 / 76 = 2
    16'b11011011_01001101 : OUT <= 2;  //219 / 77 = 2
    16'b11011011_01001110 : OUT <= 2;  //219 / 78 = 2
    16'b11011011_01001111 : OUT <= 2;  //219 / 79 = 2
    16'b11011011_01010000 : OUT <= 2;  //219 / 80 = 2
    16'b11011011_01010001 : OUT <= 2;  //219 / 81 = 2
    16'b11011011_01010010 : OUT <= 2;  //219 / 82 = 2
    16'b11011011_01010011 : OUT <= 2;  //219 / 83 = 2
    16'b11011011_01010100 : OUT <= 2;  //219 / 84 = 2
    16'b11011011_01010101 : OUT <= 2;  //219 / 85 = 2
    16'b11011011_01010110 : OUT <= 2;  //219 / 86 = 2
    16'b11011011_01010111 : OUT <= 2;  //219 / 87 = 2
    16'b11011011_01011000 : OUT <= 2;  //219 / 88 = 2
    16'b11011011_01011001 : OUT <= 2;  //219 / 89 = 2
    16'b11011011_01011010 : OUT <= 2;  //219 / 90 = 2
    16'b11011011_01011011 : OUT <= 2;  //219 / 91 = 2
    16'b11011011_01011100 : OUT <= 2;  //219 / 92 = 2
    16'b11011011_01011101 : OUT <= 2;  //219 / 93 = 2
    16'b11011011_01011110 : OUT <= 2;  //219 / 94 = 2
    16'b11011011_01011111 : OUT <= 2;  //219 / 95 = 2
    16'b11011011_01100000 : OUT <= 2;  //219 / 96 = 2
    16'b11011011_01100001 : OUT <= 2;  //219 / 97 = 2
    16'b11011011_01100010 : OUT <= 2;  //219 / 98 = 2
    16'b11011011_01100011 : OUT <= 2;  //219 / 99 = 2
    16'b11011011_01100100 : OUT <= 2;  //219 / 100 = 2
    16'b11011011_01100101 : OUT <= 2;  //219 / 101 = 2
    16'b11011011_01100110 : OUT <= 2;  //219 / 102 = 2
    16'b11011011_01100111 : OUT <= 2;  //219 / 103 = 2
    16'b11011011_01101000 : OUT <= 2;  //219 / 104 = 2
    16'b11011011_01101001 : OUT <= 2;  //219 / 105 = 2
    16'b11011011_01101010 : OUT <= 2;  //219 / 106 = 2
    16'b11011011_01101011 : OUT <= 2;  //219 / 107 = 2
    16'b11011011_01101100 : OUT <= 2;  //219 / 108 = 2
    16'b11011011_01101101 : OUT <= 2;  //219 / 109 = 2
    16'b11011011_01101110 : OUT <= 1;  //219 / 110 = 1
    16'b11011011_01101111 : OUT <= 1;  //219 / 111 = 1
    16'b11011011_01110000 : OUT <= 1;  //219 / 112 = 1
    16'b11011011_01110001 : OUT <= 1;  //219 / 113 = 1
    16'b11011011_01110010 : OUT <= 1;  //219 / 114 = 1
    16'b11011011_01110011 : OUT <= 1;  //219 / 115 = 1
    16'b11011011_01110100 : OUT <= 1;  //219 / 116 = 1
    16'b11011011_01110101 : OUT <= 1;  //219 / 117 = 1
    16'b11011011_01110110 : OUT <= 1;  //219 / 118 = 1
    16'b11011011_01110111 : OUT <= 1;  //219 / 119 = 1
    16'b11011011_01111000 : OUT <= 1;  //219 / 120 = 1
    16'b11011011_01111001 : OUT <= 1;  //219 / 121 = 1
    16'b11011011_01111010 : OUT <= 1;  //219 / 122 = 1
    16'b11011011_01111011 : OUT <= 1;  //219 / 123 = 1
    16'b11011011_01111100 : OUT <= 1;  //219 / 124 = 1
    16'b11011011_01111101 : OUT <= 1;  //219 / 125 = 1
    16'b11011011_01111110 : OUT <= 1;  //219 / 126 = 1
    16'b11011011_01111111 : OUT <= 1;  //219 / 127 = 1
    16'b11011011_10000000 : OUT <= 1;  //219 / 128 = 1
    16'b11011011_10000001 : OUT <= 1;  //219 / 129 = 1
    16'b11011011_10000010 : OUT <= 1;  //219 / 130 = 1
    16'b11011011_10000011 : OUT <= 1;  //219 / 131 = 1
    16'b11011011_10000100 : OUT <= 1;  //219 / 132 = 1
    16'b11011011_10000101 : OUT <= 1;  //219 / 133 = 1
    16'b11011011_10000110 : OUT <= 1;  //219 / 134 = 1
    16'b11011011_10000111 : OUT <= 1;  //219 / 135 = 1
    16'b11011011_10001000 : OUT <= 1;  //219 / 136 = 1
    16'b11011011_10001001 : OUT <= 1;  //219 / 137 = 1
    16'b11011011_10001010 : OUT <= 1;  //219 / 138 = 1
    16'b11011011_10001011 : OUT <= 1;  //219 / 139 = 1
    16'b11011011_10001100 : OUT <= 1;  //219 / 140 = 1
    16'b11011011_10001101 : OUT <= 1;  //219 / 141 = 1
    16'b11011011_10001110 : OUT <= 1;  //219 / 142 = 1
    16'b11011011_10001111 : OUT <= 1;  //219 / 143 = 1
    16'b11011011_10010000 : OUT <= 1;  //219 / 144 = 1
    16'b11011011_10010001 : OUT <= 1;  //219 / 145 = 1
    16'b11011011_10010010 : OUT <= 1;  //219 / 146 = 1
    16'b11011011_10010011 : OUT <= 1;  //219 / 147 = 1
    16'b11011011_10010100 : OUT <= 1;  //219 / 148 = 1
    16'b11011011_10010101 : OUT <= 1;  //219 / 149 = 1
    16'b11011011_10010110 : OUT <= 1;  //219 / 150 = 1
    16'b11011011_10010111 : OUT <= 1;  //219 / 151 = 1
    16'b11011011_10011000 : OUT <= 1;  //219 / 152 = 1
    16'b11011011_10011001 : OUT <= 1;  //219 / 153 = 1
    16'b11011011_10011010 : OUT <= 1;  //219 / 154 = 1
    16'b11011011_10011011 : OUT <= 1;  //219 / 155 = 1
    16'b11011011_10011100 : OUT <= 1;  //219 / 156 = 1
    16'b11011011_10011101 : OUT <= 1;  //219 / 157 = 1
    16'b11011011_10011110 : OUT <= 1;  //219 / 158 = 1
    16'b11011011_10011111 : OUT <= 1;  //219 / 159 = 1
    16'b11011011_10100000 : OUT <= 1;  //219 / 160 = 1
    16'b11011011_10100001 : OUT <= 1;  //219 / 161 = 1
    16'b11011011_10100010 : OUT <= 1;  //219 / 162 = 1
    16'b11011011_10100011 : OUT <= 1;  //219 / 163 = 1
    16'b11011011_10100100 : OUT <= 1;  //219 / 164 = 1
    16'b11011011_10100101 : OUT <= 1;  //219 / 165 = 1
    16'b11011011_10100110 : OUT <= 1;  //219 / 166 = 1
    16'b11011011_10100111 : OUT <= 1;  //219 / 167 = 1
    16'b11011011_10101000 : OUT <= 1;  //219 / 168 = 1
    16'b11011011_10101001 : OUT <= 1;  //219 / 169 = 1
    16'b11011011_10101010 : OUT <= 1;  //219 / 170 = 1
    16'b11011011_10101011 : OUT <= 1;  //219 / 171 = 1
    16'b11011011_10101100 : OUT <= 1;  //219 / 172 = 1
    16'b11011011_10101101 : OUT <= 1;  //219 / 173 = 1
    16'b11011011_10101110 : OUT <= 1;  //219 / 174 = 1
    16'b11011011_10101111 : OUT <= 1;  //219 / 175 = 1
    16'b11011011_10110000 : OUT <= 1;  //219 / 176 = 1
    16'b11011011_10110001 : OUT <= 1;  //219 / 177 = 1
    16'b11011011_10110010 : OUT <= 1;  //219 / 178 = 1
    16'b11011011_10110011 : OUT <= 1;  //219 / 179 = 1
    16'b11011011_10110100 : OUT <= 1;  //219 / 180 = 1
    16'b11011011_10110101 : OUT <= 1;  //219 / 181 = 1
    16'b11011011_10110110 : OUT <= 1;  //219 / 182 = 1
    16'b11011011_10110111 : OUT <= 1;  //219 / 183 = 1
    16'b11011011_10111000 : OUT <= 1;  //219 / 184 = 1
    16'b11011011_10111001 : OUT <= 1;  //219 / 185 = 1
    16'b11011011_10111010 : OUT <= 1;  //219 / 186 = 1
    16'b11011011_10111011 : OUT <= 1;  //219 / 187 = 1
    16'b11011011_10111100 : OUT <= 1;  //219 / 188 = 1
    16'b11011011_10111101 : OUT <= 1;  //219 / 189 = 1
    16'b11011011_10111110 : OUT <= 1;  //219 / 190 = 1
    16'b11011011_10111111 : OUT <= 1;  //219 / 191 = 1
    16'b11011011_11000000 : OUT <= 1;  //219 / 192 = 1
    16'b11011011_11000001 : OUT <= 1;  //219 / 193 = 1
    16'b11011011_11000010 : OUT <= 1;  //219 / 194 = 1
    16'b11011011_11000011 : OUT <= 1;  //219 / 195 = 1
    16'b11011011_11000100 : OUT <= 1;  //219 / 196 = 1
    16'b11011011_11000101 : OUT <= 1;  //219 / 197 = 1
    16'b11011011_11000110 : OUT <= 1;  //219 / 198 = 1
    16'b11011011_11000111 : OUT <= 1;  //219 / 199 = 1
    16'b11011011_11001000 : OUT <= 1;  //219 / 200 = 1
    16'b11011011_11001001 : OUT <= 1;  //219 / 201 = 1
    16'b11011011_11001010 : OUT <= 1;  //219 / 202 = 1
    16'b11011011_11001011 : OUT <= 1;  //219 / 203 = 1
    16'b11011011_11001100 : OUT <= 1;  //219 / 204 = 1
    16'b11011011_11001101 : OUT <= 1;  //219 / 205 = 1
    16'b11011011_11001110 : OUT <= 1;  //219 / 206 = 1
    16'b11011011_11001111 : OUT <= 1;  //219 / 207 = 1
    16'b11011011_11010000 : OUT <= 1;  //219 / 208 = 1
    16'b11011011_11010001 : OUT <= 1;  //219 / 209 = 1
    16'b11011011_11010010 : OUT <= 1;  //219 / 210 = 1
    16'b11011011_11010011 : OUT <= 1;  //219 / 211 = 1
    16'b11011011_11010100 : OUT <= 1;  //219 / 212 = 1
    16'b11011011_11010101 : OUT <= 1;  //219 / 213 = 1
    16'b11011011_11010110 : OUT <= 1;  //219 / 214 = 1
    16'b11011011_11010111 : OUT <= 1;  //219 / 215 = 1
    16'b11011011_11011000 : OUT <= 1;  //219 / 216 = 1
    16'b11011011_11011001 : OUT <= 1;  //219 / 217 = 1
    16'b11011011_11011010 : OUT <= 1;  //219 / 218 = 1
    16'b11011011_11011011 : OUT <= 1;  //219 / 219 = 1
    16'b11011011_11011100 : OUT <= 0;  //219 / 220 = 0
    16'b11011011_11011101 : OUT <= 0;  //219 / 221 = 0
    16'b11011011_11011110 : OUT <= 0;  //219 / 222 = 0
    16'b11011011_11011111 : OUT <= 0;  //219 / 223 = 0
    16'b11011011_11100000 : OUT <= 0;  //219 / 224 = 0
    16'b11011011_11100001 : OUT <= 0;  //219 / 225 = 0
    16'b11011011_11100010 : OUT <= 0;  //219 / 226 = 0
    16'b11011011_11100011 : OUT <= 0;  //219 / 227 = 0
    16'b11011011_11100100 : OUT <= 0;  //219 / 228 = 0
    16'b11011011_11100101 : OUT <= 0;  //219 / 229 = 0
    16'b11011011_11100110 : OUT <= 0;  //219 / 230 = 0
    16'b11011011_11100111 : OUT <= 0;  //219 / 231 = 0
    16'b11011011_11101000 : OUT <= 0;  //219 / 232 = 0
    16'b11011011_11101001 : OUT <= 0;  //219 / 233 = 0
    16'b11011011_11101010 : OUT <= 0;  //219 / 234 = 0
    16'b11011011_11101011 : OUT <= 0;  //219 / 235 = 0
    16'b11011011_11101100 : OUT <= 0;  //219 / 236 = 0
    16'b11011011_11101101 : OUT <= 0;  //219 / 237 = 0
    16'b11011011_11101110 : OUT <= 0;  //219 / 238 = 0
    16'b11011011_11101111 : OUT <= 0;  //219 / 239 = 0
    16'b11011011_11110000 : OUT <= 0;  //219 / 240 = 0
    16'b11011011_11110001 : OUT <= 0;  //219 / 241 = 0
    16'b11011011_11110010 : OUT <= 0;  //219 / 242 = 0
    16'b11011011_11110011 : OUT <= 0;  //219 / 243 = 0
    16'b11011011_11110100 : OUT <= 0;  //219 / 244 = 0
    16'b11011011_11110101 : OUT <= 0;  //219 / 245 = 0
    16'b11011011_11110110 : OUT <= 0;  //219 / 246 = 0
    16'b11011011_11110111 : OUT <= 0;  //219 / 247 = 0
    16'b11011011_11111000 : OUT <= 0;  //219 / 248 = 0
    16'b11011011_11111001 : OUT <= 0;  //219 / 249 = 0
    16'b11011011_11111010 : OUT <= 0;  //219 / 250 = 0
    16'b11011011_11111011 : OUT <= 0;  //219 / 251 = 0
    16'b11011011_11111100 : OUT <= 0;  //219 / 252 = 0
    16'b11011011_11111101 : OUT <= 0;  //219 / 253 = 0
    16'b11011011_11111110 : OUT <= 0;  //219 / 254 = 0
    16'b11011011_11111111 : OUT <= 0;  //219 / 255 = 0
    16'b11011100_00000000 : OUT <= 0;  //220 / 0 = 0
    16'b11011100_00000001 : OUT <= 220;  //220 / 1 = 220
    16'b11011100_00000010 : OUT <= 110;  //220 / 2 = 110
    16'b11011100_00000011 : OUT <= 73;  //220 / 3 = 73
    16'b11011100_00000100 : OUT <= 55;  //220 / 4 = 55
    16'b11011100_00000101 : OUT <= 44;  //220 / 5 = 44
    16'b11011100_00000110 : OUT <= 36;  //220 / 6 = 36
    16'b11011100_00000111 : OUT <= 31;  //220 / 7 = 31
    16'b11011100_00001000 : OUT <= 27;  //220 / 8 = 27
    16'b11011100_00001001 : OUT <= 24;  //220 / 9 = 24
    16'b11011100_00001010 : OUT <= 22;  //220 / 10 = 22
    16'b11011100_00001011 : OUT <= 20;  //220 / 11 = 20
    16'b11011100_00001100 : OUT <= 18;  //220 / 12 = 18
    16'b11011100_00001101 : OUT <= 16;  //220 / 13 = 16
    16'b11011100_00001110 : OUT <= 15;  //220 / 14 = 15
    16'b11011100_00001111 : OUT <= 14;  //220 / 15 = 14
    16'b11011100_00010000 : OUT <= 13;  //220 / 16 = 13
    16'b11011100_00010001 : OUT <= 12;  //220 / 17 = 12
    16'b11011100_00010010 : OUT <= 12;  //220 / 18 = 12
    16'b11011100_00010011 : OUT <= 11;  //220 / 19 = 11
    16'b11011100_00010100 : OUT <= 11;  //220 / 20 = 11
    16'b11011100_00010101 : OUT <= 10;  //220 / 21 = 10
    16'b11011100_00010110 : OUT <= 10;  //220 / 22 = 10
    16'b11011100_00010111 : OUT <= 9;  //220 / 23 = 9
    16'b11011100_00011000 : OUT <= 9;  //220 / 24 = 9
    16'b11011100_00011001 : OUT <= 8;  //220 / 25 = 8
    16'b11011100_00011010 : OUT <= 8;  //220 / 26 = 8
    16'b11011100_00011011 : OUT <= 8;  //220 / 27 = 8
    16'b11011100_00011100 : OUT <= 7;  //220 / 28 = 7
    16'b11011100_00011101 : OUT <= 7;  //220 / 29 = 7
    16'b11011100_00011110 : OUT <= 7;  //220 / 30 = 7
    16'b11011100_00011111 : OUT <= 7;  //220 / 31 = 7
    16'b11011100_00100000 : OUT <= 6;  //220 / 32 = 6
    16'b11011100_00100001 : OUT <= 6;  //220 / 33 = 6
    16'b11011100_00100010 : OUT <= 6;  //220 / 34 = 6
    16'b11011100_00100011 : OUT <= 6;  //220 / 35 = 6
    16'b11011100_00100100 : OUT <= 6;  //220 / 36 = 6
    16'b11011100_00100101 : OUT <= 5;  //220 / 37 = 5
    16'b11011100_00100110 : OUT <= 5;  //220 / 38 = 5
    16'b11011100_00100111 : OUT <= 5;  //220 / 39 = 5
    16'b11011100_00101000 : OUT <= 5;  //220 / 40 = 5
    16'b11011100_00101001 : OUT <= 5;  //220 / 41 = 5
    16'b11011100_00101010 : OUT <= 5;  //220 / 42 = 5
    16'b11011100_00101011 : OUT <= 5;  //220 / 43 = 5
    16'b11011100_00101100 : OUT <= 5;  //220 / 44 = 5
    16'b11011100_00101101 : OUT <= 4;  //220 / 45 = 4
    16'b11011100_00101110 : OUT <= 4;  //220 / 46 = 4
    16'b11011100_00101111 : OUT <= 4;  //220 / 47 = 4
    16'b11011100_00110000 : OUT <= 4;  //220 / 48 = 4
    16'b11011100_00110001 : OUT <= 4;  //220 / 49 = 4
    16'b11011100_00110010 : OUT <= 4;  //220 / 50 = 4
    16'b11011100_00110011 : OUT <= 4;  //220 / 51 = 4
    16'b11011100_00110100 : OUT <= 4;  //220 / 52 = 4
    16'b11011100_00110101 : OUT <= 4;  //220 / 53 = 4
    16'b11011100_00110110 : OUT <= 4;  //220 / 54 = 4
    16'b11011100_00110111 : OUT <= 4;  //220 / 55 = 4
    16'b11011100_00111000 : OUT <= 3;  //220 / 56 = 3
    16'b11011100_00111001 : OUT <= 3;  //220 / 57 = 3
    16'b11011100_00111010 : OUT <= 3;  //220 / 58 = 3
    16'b11011100_00111011 : OUT <= 3;  //220 / 59 = 3
    16'b11011100_00111100 : OUT <= 3;  //220 / 60 = 3
    16'b11011100_00111101 : OUT <= 3;  //220 / 61 = 3
    16'b11011100_00111110 : OUT <= 3;  //220 / 62 = 3
    16'b11011100_00111111 : OUT <= 3;  //220 / 63 = 3
    16'b11011100_01000000 : OUT <= 3;  //220 / 64 = 3
    16'b11011100_01000001 : OUT <= 3;  //220 / 65 = 3
    16'b11011100_01000010 : OUT <= 3;  //220 / 66 = 3
    16'b11011100_01000011 : OUT <= 3;  //220 / 67 = 3
    16'b11011100_01000100 : OUT <= 3;  //220 / 68 = 3
    16'b11011100_01000101 : OUT <= 3;  //220 / 69 = 3
    16'b11011100_01000110 : OUT <= 3;  //220 / 70 = 3
    16'b11011100_01000111 : OUT <= 3;  //220 / 71 = 3
    16'b11011100_01001000 : OUT <= 3;  //220 / 72 = 3
    16'b11011100_01001001 : OUT <= 3;  //220 / 73 = 3
    16'b11011100_01001010 : OUT <= 2;  //220 / 74 = 2
    16'b11011100_01001011 : OUT <= 2;  //220 / 75 = 2
    16'b11011100_01001100 : OUT <= 2;  //220 / 76 = 2
    16'b11011100_01001101 : OUT <= 2;  //220 / 77 = 2
    16'b11011100_01001110 : OUT <= 2;  //220 / 78 = 2
    16'b11011100_01001111 : OUT <= 2;  //220 / 79 = 2
    16'b11011100_01010000 : OUT <= 2;  //220 / 80 = 2
    16'b11011100_01010001 : OUT <= 2;  //220 / 81 = 2
    16'b11011100_01010010 : OUT <= 2;  //220 / 82 = 2
    16'b11011100_01010011 : OUT <= 2;  //220 / 83 = 2
    16'b11011100_01010100 : OUT <= 2;  //220 / 84 = 2
    16'b11011100_01010101 : OUT <= 2;  //220 / 85 = 2
    16'b11011100_01010110 : OUT <= 2;  //220 / 86 = 2
    16'b11011100_01010111 : OUT <= 2;  //220 / 87 = 2
    16'b11011100_01011000 : OUT <= 2;  //220 / 88 = 2
    16'b11011100_01011001 : OUT <= 2;  //220 / 89 = 2
    16'b11011100_01011010 : OUT <= 2;  //220 / 90 = 2
    16'b11011100_01011011 : OUT <= 2;  //220 / 91 = 2
    16'b11011100_01011100 : OUT <= 2;  //220 / 92 = 2
    16'b11011100_01011101 : OUT <= 2;  //220 / 93 = 2
    16'b11011100_01011110 : OUT <= 2;  //220 / 94 = 2
    16'b11011100_01011111 : OUT <= 2;  //220 / 95 = 2
    16'b11011100_01100000 : OUT <= 2;  //220 / 96 = 2
    16'b11011100_01100001 : OUT <= 2;  //220 / 97 = 2
    16'b11011100_01100010 : OUT <= 2;  //220 / 98 = 2
    16'b11011100_01100011 : OUT <= 2;  //220 / 99 = 2
    16'b11011100_01100100 : OUT <= 2;  //220 / 100 = 2
    16'b11011100_01100101 : OUT <= 2;  //220 / 101 = 2
    16'b11011100_01100110 : OUT <= 2;  //220 / 102 = 2
    16'b11011100_01100111 : OUT <= 2;  //220 / 103 = 2
    16'b11011100_01101000 : OUT <= 2;  //220 / 104 = 2
    16'b11011100_01101001 : OUT <= 2;  //220 / 105 = 2
    16'b11011100_01101010 : OUT <= 2;  //220 / 106 = 2
    16'b11011100_01101011 : OUT <= 2;  //220 / 107 = 2
    16'b11011100_01101100 : OUT <= 2;  //220 / 108 = 2
    16'b11011100_01101101 : OUT <= 2;  //220 / 109 = 2
    16'b11011100_01101110 : OUT <= 2;  //220 / 110 = 2
    16'b11011100_01101111 : OUT <= 1;  //220 / 111 = 1
    16'b11011100_01110000 : OUT <= 1;  //220 / 112 = 1
    16'b11011100_01110001 : OUT <= 1;  //220 / 113 = 1
    16'b11011100_01110010 : OUT <= 1;  //220 / 114 = 1
    16'b11011100_01110011 : OUT <= 1;  //220 / 115 = 1
    16'b11011100_01110100 : OUT <= 1;  //220 / 116 = 1
    16'b11011100_01110101 : OUT <= 1;  //220 / 117 = 1
    16'b11011100_01110110 : OUT <= 1;  //220 / 118 = 1
    16'b11011100_01110111 : OUT <= 1;  //220 / 119 = 1
    16'b11011100_01111000 : OUT <= 1;  //220 / 120 = 1
    16'b11011100_01111001 : OUT <= 1;  //220 / 121 = 1
    16'b11011100_01111010 : OUT <= 1;  //220 / 122 = 1
    16'b11011100_01111011 : OUT <= 1;  //220 / 123 = 1
    16'b11011100_01111100 : OUT <= 1;  //220 / 124 = 1
    16'b11011100_01111101 : OUT <= 1;  //220 / 125 = 1
    16'b11011100_01111110 : OUT <= 1;  //220 / 126 = 1
    16'b11011100_01111111 : OUT <= 1;  //220 / 127 = 1
    16'b11011100_10000000 : OUT <= 1;  //220 / 128 = 1
    16'b11011100_10000001 : OUT <= 1;  //220 / 129 = 1
    16'b11011100_10000010 : OUT <= 1;  //220 / 130 = 1
    16'b11011100_10000011 : OUT <= 1;  //220 / 131 = 1
    16'b11011100_10000100 : OUT <= 1;  //220 / 132 = 1
    16'b11011100_10000101 : OUT <= 1;  //220 / 133 = 1
    16'b11011100_10000110 : OUT <= 1;  //220 / 134 = 1
    16'b11011100_10000111 : OUT <= 1;  //220 / 135 = 1
    16'b11011100_10001000 : OUT <= 1;  //220 / 136 = 1
    16'b11011100_10001001 : OUT <= 1;  //220 / 137 = 1
    16'b11011100_10001010 : OUT <= 1;  //220 / 138 = 1
    16'b11011100_10001011 : OUT <= 1;  //220 / 139 = 1
    16'b11011100_10001100 : OUT <= 1;  //220 / 140 = 1
    16'b11011100_10001101 : OUT <= 1;  //220 / 141 = 1
    16'b11011100_10001110 : OUT <= 1;  //220 / 142 = 1
    16'b11011100_10001111 : OUT <= 1;  //220 / 143 = 1
    16'b11011100_10010000 : OUT <= 1;  //220 / 144 = 1
    16'b11011100_10010001 : OUT <= 1;  //220 / 145 = 1
    16'b11011100_10010010 : OUT <= 1;  //220 / 146 = 1
    16'b11011100_10010011 : OUT <= 1;  //220 / 147 = 1
    16'b11011100_10010100 : OUT <= 1;  //220 / 148 = 1
    16'b11011100_10010101 : OUT <= 1;  //220 / 149 = 1
    16'b11011100_10010110 : OUT <= 1;  //220 / 150 = 1
    16'b11011100_10010111 : OUT <= 1;  //220 / 151 = 1
    16'b11011100_10011000 : OUT <= 1;  //220 / 152 = 1
    16'b11011100_10011001 : OUT <= 1;  //220 / 153 = 1
    16'b11011100_10011010 : OUT <= 1;  //220 / 154 = 1
    16'b11011100_10011011 : OUT <= 1;  //220 / 155 = 1
    16'b11011100_10011100 : OUT <= 1;  //220 / 156 = 1
    16'b11011100_10011101 : OUT <= 1;  //220 / 157 = 1
    16'b11011100_10011110 : OUT <= 1;  //220 / 158 = 1
    16'b11011100_10011111 : OUT <= 1;  //220 / 159 = 1
    16'b11011100_10100000 : OUT <= 1;  //220 / 160 = 1
    16'b11011100_10100001 : OUT <= 1;  //220 / 161 = 1
    16'b11011100_10100010 : OUT <= 1;  //220 / 162 = 1
    16'b11011100_10100011 : OUT <= 1;  //220 / 163 = 1
    16'b11011100_10100100 : OUT <= 1;  //220 / 164 = 1
    16'b11011100_10100101 : OUT <= 1;  //220 / 165 = 1
    16'b11011100_10100110 : OUT <= 1;  //220 / 166 = 1
    16'b11011100_10100111 : OUT <= 1;  //220 / 167 = 1
    16'b11011100_10101000 : OUT <= 1;  //220 / 168 = 1
    16'b11011100_10101001 : OUT <= 1;  //220 / 169 = 1
    16'b11011100_10101010 : OUT <= 1;  //220 / 170 = 1
    16'b11011100_10101011 : OUT <= 1;  //220 / 171 = 1
    16'b11011100_10101100 : OUT <= 1;  //220 / 172 = 1
    16'b11011100_10101101 : OUT <= 1;  //220 / 173 = 1
    16'b11011100_10101110 : OUT <= 1;  //220 / 174 = 1
    16'b11011100_10101111 : OUT <= 1;  //220 / 175 = 1
    16'b11011100_10110000 : OUT <= 1;  //220 / 176 = 1
    16'b11011100_10110001 : OUT <= 1;  //220 / 177 = 1
    16'b11011100_10110010 : OUT <= 1;  //220 / 178 = 1
    16'b11011100_10110011 : OUT <= 1;  //220 / 179 = 1
    16'b11011100_10110100 : OUT <= 1;  //220 / 180 = 1
    16'b11011100_10110101 : OUT <= 1;  //220 / 181 = 1
    16'b11011100_10110110 : OUT <= 1;  //220 / 182 = 1
    16'b11011100_10110111 : OUT <= 1;  //220 / 183 = 1
    16'b11011100_10111000 : OUT <= 1;  //220 / 184 = 1
    16'b11011100_10111001 : OUT <= 1;  //220 / 185 = 1
    16'b11011100_10111010 : OUT <= 1;  //220 / 186 = 1
    16'b11011100_10111011 : OUT <= 1;  //220 / 187 = 1
    16'b11011100_10111100 : OUT <= 1;  //220 / 188 = 1
    16'b11011100_10111101 : OUT <= 1;  //220 / 189 = 1
    16'b11011100_10111110 : OUT <= 1;  //220 / 190 = 1
    16'b11011100_10111111 : OUT <= 1;  //220 / 191 = 1
    16'b11011100_11000000 : OUT <= 1;  //220 / 192 = 1
    16'b11011100_11000001 : OUT <= 1;  //220 / 193 = 1
    16'b11011100_11000010 : OUT <= 1;  //220 / 194 = 1
    16'b11011100_11000011 : OUT <= 1;  //220 / 195 = 1
    16'b11011100_11000100 : OUT <= 1;  //220 / 196 = 1
    16'b11011100_11000101 : OUT <= 1;  //220 / 197 = 1
    16'b11011100_11000110 : OUT <= 1;  //220 / 198 = 1
    16'b11011100_11000111 : OUT <= 1;  //220 / 199 = 1
    16'b11011100_11001000 : OUT <= 1;  //220 / 200 = 1
    16'b11011100_11001001 : OUT <= 1;  //220 / 201 = 1
    16'b11011100_11001010 : OUT <= 1;  //220 / 202 = 1
    16'b11011100_11001011 : OUT <= 1;  //220 / 203 = 1
    16'b11011100_11001100 : OUT <= 1;  //220 / 204 = 1
    16'b11011100_11001101 : OUT <= 1;  //220 / 205 = 1
    16'b11011100_11001110 : OUT <= 1;  //220 / 206 = 1
    16'b11011100_11001111 : OUT <= 1;  //220 / 207 = 1
    16'b11011100_11010000 : OUT <= 1;  //220 / 208 = 1
    16'b11011100_11010001 : OUT <= 1;  //220 / 209 = 1
    16'b11011100_11010010 : OUT <= 1;  //220 / 210 = 1
    16'b11011100_11010011 : OUT <= 1;  //220 / 211 = 1
    16'b11011100_11010100 : OUT <= 1;  //220 / 212 = 1
    16'b11011100_11010101 : OUT <= 1;  //220 / 213 = 1
    16'b11011100_11010110 : OUT <= 1;  //220 / 214 = 1
    16'b11011100_11010111 : OUT <= 1;  //220 / 215 = 1
    16'b11011100_11011000 : OUT <= 1;  //220 / 216 = 1
    16'b11011100_11011001 : OUT <= 1;  //220 / 217 = 1
    16'b11011100_11011010 : OUT <= 1;  //220 / 218 = 1
    16'b11011100_11011011 : OUT <= 1;  //220 / 219 = 1
    16'b11011100_11011100 : OUT <= 1;  //220 / 220 = 1
    16'b11011100_11011101 : OUT <= 0;  //220 / 221 = 0
    16'b11011100_11011110 : OUT <= 0;  //220 / 222 = 0
    16'b11011100_11011111 : OUT <= 0;  //220 / 223 = 0
    16'b11011100_11100000 : OUT <= 0;  //220 / 224 = 0
    16'b11011100_11100001 : OUT <= 0;  //220 / 225 = 0
    16'b11011100_11100010 : OUT <= 0;  //220 / 226 = 0
    16'b11011100_11100011 : OUT <= 0;  //220 / 227 = 0
    16'b11011100_11100100 : OUT <= 0;  //220 / 228 = 0
    16'b11011100_11100101 : OUT <= 0;  //220 / 229 = 0
    16'b11011100_11100110 : OUT <= 0;  //220 / 230 = 0
    16'b11011100_11100111 : OUT <= 0;  //220 / 231 = 0
    16'b11011100_11101000 : OUT <= 0;  //220 / 232 = 0
    16'b11011100_11101001 : OUT <= 0;  //220 / 233 = 0
    16'b11011100_11101010 : OUT <= 0;  //220 / 234 = 0
    16'b11011100_11101011 : OUT <= 0;  //220 / 235 = 0
    16'b11011100_11101100 : OUT <= 0;  //220 / 236 = 0
    16'b11011100_11101101 : OUT <= 0;  //220 / 237 = 0
    16'b11011100_11101110 : OUT <= 0;  //220 / 238 = 0
    16'b11011100_11101111 : OUT <= 0;  //220 / 239 = 0
    16'b11011100_11110000 : OUT <= 0;  //220 / 240 = 0
    16'b11011100_11110001 : OUT <= 0;  //220 / 241 = 0
    16'b11011100_11110010 : OUT <= 0;  //220 / 242 = 0
    16'b11011100_11110011 : OUT <= 0;  //220 / 243 = 0
    16'b11011100_11110100 : OUT <= 0;  //220 / 244 = 0
    16'b11011100_11110101 : OUT <= 0;  //220 / 245 = 0
    16'b11011100_11110110 : OUT <= 0;  //220 / 246 = 0
    16'b11011100_11110111 : OUT <= 0;  //220 / 247 = 0
    16'b11011100_11111000 : OUT <= 0;  //220 / 248 = 0
    16'b11011100_11111001 : OUT <= 0;  //220 / 249 = 0
    16'b11011100_11111010 : OUT <= 0;  //220 / 250 = 0
    16'b11011100_11111011 : OUT <= 0;  //220 / 251 = 0
    16'b11011100_11111100 : OUT <= 0;  //220 / 252 = 0
    16'b11011100_11111101 : OUT <= 0;  //220 / 253 = 0
    16'b11011100_11111110 : OUT <= 0;  //220 / 254 = 0
    16'b11011100_11111111 : OUT <= 0;  //220 / 255 = 0
    16'b11011101_00000000 : OUT <= 0;  //221 / 0 = 0
    16'b11011101_00000001 : OUT <= 221;  //221 / 1 = 221
    16'b11011101_00000010 : OUT <= 110;  //221 / 2 = 110
    16'b11011101_00000011 : OUT <= 73;  //221 / 3 = 73
    16'b11011101_00000100 : OUT <= 55;  //221 / 4 = 55
    16'b11011101_00000101 : OUT <= 44;  //221 / 5 = 44
    16'b11011101_00000110 : OUT <= 36;  //221 / 6 = 36
    16'b11011101_00000111 : OUT <= 31;  //221 / 7 = 31
    16'b11011101_00001000 : OUT <= 27;  //221 / 8 = 27
    16'b11011101_00001001 : OUT <= 24;  //221 / 9 = 24
    16'b11011101_00001010 : OUT <= 22;  //221 / 10 = 22
    16'b11011101_00001011 : OUT <= 20;  //221 / 11 = 20
    16'b11011101_00001100 : OUT <= 18;  //221 / 12 = 18
    16'b11011101_00001101 : OUT <= 17;  //221 / 13 = 17
    16'b11011101_00001110 : OUT <= 15;  //221 / 14 = 15
    16'b11011101_00001111 : OUT <= 14;  //221 / 15 = 14
    16'b11011101_00010000 : OUT <= 13;  //221 / 16 = 13
    16'b11011101_00010001 : OUT <= 13;  //221 / 17 = 13
    16'b11011101_00010010 : OUT <= 12;  //221 / 18 = 12
    16'b11011101_00010011 : OUT <= 11;  //221 / 19 = 11
    16'b11011101_00010100 : OUT <= 11;  //221 / 20 = 11
    16'b11011101_00010101 : OUT <= 10;  //221 / 21 = 10
    16'b11011101_00010110 : OUT <= 10;  //221 / 22 = 10
    16'b11011101_00010111 : OUT <= 9;  //221 / 23 = 9
    16'b11011101_00011000 : OUT <= 9;  //221 / 24 = 9
    16'b11011101_00011001 : OUT <= 8;  //221 / 25 = 8
    16'b11011101_00011010 : OUT <= 8;  //221 / 26 = 8
    16'b11011101_00011011 : OUT <= 8;  //221 / 27 = 8
    16'b11011101_00011100 : OUT <= 7;  //221 / 28 = 7
    16'b11011101_00011101 : OUT <= 7;  //221 / 29 = 7
    16'b11011101_00011110 : OUT <= 7;  //221 / 30 = 7
    16'b11011101_00011111 : OUT <= 7;  //221 / 31 = 7
    16'b11011101_00100000 : OUT <= 6;  //221 / 32 = 6
    16'b11011101_00100001 : OUT <= 6;  //221 / 33 = 6
    16'b11011101_00100010 : OUT <= 6;  //221 / 34 = 6
    16'b11011101_00100011 : OUT <= 6;  //221 / 35 = 6
    16'b11011101_00100100 : OUT <= 6;  //221 / 36 = 6
    16'b11011101_00100101 : OUT <= 5;  //221 / 37 = 5
    16'b11011101_00100110 : OUT <= 5;  //221 / 38 = 5
    16'b11011101_00100111 : OUT <= 5;  //221 / 39 = 5
    16'b11011101_00101000 : OUT <= 5;  //221 / 40 = 5
    16'b11011101_00101001 : OUT <= 5;  //221 / 41 = 5
    16'b11011101_00101010 : OUT <= 5;  //221 / 42 = 5
    16'b11011101_00101011 : OUT <= 5;  //221 / 43 = 5
    16'b11011101_00101100 : OUT <= 5;  //221 / 44 = 5
    16'b11011101_00101101 : OUT <= 4;  //221 / 45 = 4
    16'b11011101_00101110 : OUT <= 4;  //221 / 46 = 4
    16'b11011101_00101111 : OUT <= 4;  //221 / 47 = 4
    16'b11011101_00110000 : OUT <= 4;  //221 / 48 = 4
    16'b11011101_00110001 : OUT <= 4;  //221 / 49 = 4
    16'b11011101_00110010 : OUT <= 4;  //221 / 50 = 4
    16'b11011101_00110011 : OUT <= 4;  //221 / 51 = 4
    16'b11011101_00110100 : OUT <= 4;  //221 / 52 = 4
    16'b11011101_00110101 : OUT <= 4;  //221 / 53 = 4
    16'b11011101_00110110 : OUT <= 4;  //221 / 54 = 4
    16'b11011101_00110111 : OUT <= 4;  //221 / 55 = 4
    16'b11011101_00111000 : OUT <= 3;  //221 / 56 = 3
    16'b11011101_00111001 : OUT <= 3;  //221 / 57 = 3
    16'b11011101_00111010 : OUT <= 3;  //221 / 58 = 3
    16'b11011101_00111011 : OUT <= 3;  //221 / 59 = 3
    16'b11011101_00111100 : OUT <= 3;  //221 / 60 = 3
    16'b11011101_00111101 : OUT <= 3;  //221 / 61 = 3
    16'b11011101_00111110 : OUT <= 3;  //221 / 62 = 3
    16'b11011101_00111111 : OUT <= 3;  //221 / 63 = 3
    16'b11011101_01000000 : OUT <= 3;  //221 / 64 = 3
    16'b11011101_01000001 : OUT <= 3;  //221 / 65 = 3
    16'b11011101_01000010 : OUT <= 3;  //221 / 66 = 3
    16'b11011101_01000011 : OUT <= 3;  //221 / 67 = 3
    16'b11011101_01000100 : OUT <= 3;  //221 / 68 = 3
    16'b11011101_01000101 : OUT <= 3;  //221 / 69 = 3
    16'b11011101_01000110 : OUT <= 3;  //221 / 70 = 3
    16'b11011101_01000111 : OUT <= 3;  //221 / 71 = 3
    16'b11011101_01001000 : OUT <= 3;  //221 / 72 = 3
    16'b11011101_01001001 : OUT <= 3;  //221 / 73 = 3
    16'b11011101_01001010 : OUT <= 2;  //221 / 74 = 2
    16'b11011101_01001011 : OUT <= 2;  //221 / 75 = 2
    16'b11011101_01001100 : OUT <= 2;  //221 / 76 = 2
    16'b11011101_01001101 : OUT <= 2;  //221 / 77 = 2
    16'b11011101_01001110 : OUT <= 2;  //221 / 78 = 2
    16'b11011101_01001111 : OUT <= 2;  //221 / 79 = 2
    16'b11011101_01010000 : OUT <= 2;  //221 / 80 = 2
    16'b11011101_01010001 : OUT <= 2;  //221 / 81 = 2
    16'b11011101_01010010 : OUT <= 2;  //221 / 82 = 2
    16'b11011101_01010011 : OUT <= 2;  //221 / 83 = 2
    16'b11011101_01010100 : OUT <= 2;  //221 / 84 = 2
    16'b11011101_01010101 : OUT <= 2;  //221 / 85 = 2
    16'b11011101_01010110 : OUT <= 2;  //221 / 86 = 2
    16'b11011101_01010111 : OUT <= 2;  //221 / 87 = 2
    16'b11011101_01011000 : OUT <= 2;  //221 / 88 = 2
    16'b11011101_01011001 : OUT <= 2;  //221 / 89 = 2
    16'b11011101_01011010 : OUT <= 2;  //221 / 90 = 2
    16'b11011101_01011011 : OUT <= 2;  //221 / 91 = 2
    16'b11011101_01011100 : OUT <= 2;  //221 / 92 = 2
    16'b11011101_01011101 : OUT <= 2;  //221 / 93 = 2
    16'b11011101_01011110 : OUT <= 2;  //221 / 94 = 2
    16'b11011101_01011111 : OUT <= 2;  //221 / 95 = 2
    16'b11011101_01100000 : OUT <= 2;  //221 / 96 = 2
    16'b11011101_01100001 : OUT <= 2;  //221 / 97 = 2
    16'b11011101_01100010 : OUT <= 2;  //221 / 98 = 2
    16'b11011101_01100011 : OUT <= 2;  //221 / 99 = 2
    16'b11011101_01100100 : OUT <= 2;  //221 / 100 = 2
    16'b11011101_01100101 : OUT <= 2;  //221 / 101 = 2
    16'b11011101_01100110 : OUT <= 2;  //221 / 102 = 2
    16'b11011101_01100111 : OUT <= 2;  //221 / 103 = 2
    16'b11011101_01101000 : OUT <= 2;  //221 / 104 = 2
    16'b11011101_01101001 : OUT <= 2;  //221 / 105 = 2
    16'b11011101_01101010 : OUT <= 2;  //221 / 106 = 2
    16'b11011101_01101011 : OUT <= 2;  //221 / 107 = 2
    16'b11011101_01101100 : OUT <= 2;  //221 / 108 = 2
    16'b11011101_01101101 : OUT <= 2;  //221 / 109 = 2
    16'b11011101_01101110 : OUT <= 2;  //221 / 110 = 2
    16'b11011101_01101111 : OUT <= 1;  //221 / 111 = 1
    16'b11011101_01110000 : OUT <= 1;  //221 / 112 = 1
    16'b11011101_01110001 : OUT <= 1;  //221 / 113 = 1
    16'b11011101_01110010 : OUT <= 1;  //221 / 114 = 1
    16'b11011101_01110011 : OUT <= 1;  //221 / 115 = 1
    16'b11011101_01110100 : OUT <= 1;  //221 / 116 = 1
    16'b11011101_01110101 : OUT <= 1;  //221 / 117 = 1
    16'b11011101_01110110 : OUT <= 1;  //221 / 118 = 1
    16'b11011101_01110111 : OUT <= 1;  //221 / 119 = 1
    16'b11011101_01111000 : OUT <= 1;  //221 / 120 = 1
    16'b11011101_01111001 : OUT <= 1;  //221 / 121 = 1
    16'b11011101_01111010 : OUT <= 1;  //221 / 122 = 1
    16'b11011101_01111011 : OUT <= 1;  //221 / 123 = 1
    16'b11011101_01111100 : OUT <= 1;  //221 / 124 = 1
    16'b11011101_01111101 : OUT <= 1;  //221 / 125 = 1
    16'b11011101_01111110 : OUT <= 1;  //221 / 126 = 1
    16'b11011101_01111111 : OUT <= 1;  //221 / 127 = 1
    16'b11011101_10000000 : OUT <= 1;  //221 / 128 = 1
    16'b11011101_10000001 : OUT <= 1;  //221 / 129 = 1
    16'b11011101_10000010 : OUT <= 1;  //221 / 130 = 1
    16'b11011101_10000011 : OUT <= 1;  //221 / 131 = 1
    16'b11011101_10000100 : OUT <= 1;  //221 / 132 = 1
    16'b11011101_10000101 : OUT <= 1;  //221 / 133 = 1
    16'b11011101_10000110 : OUT <= 1;  //221 / 134 = 1
    16'b11011101_10000111 : OUT <= 1;  //221 / 135 = 1
    16'b11011101_10001000 : OUT <= 1;  //221 / 136 = 1
    16'b11011101_10001001 : OUT <= 1;  //221 / 137 = 1
    16'b11011101_10001010 : OUT <= 1;  //221 / 138 = 1
    16'b11011101_10001011 : OUT <= 1;  //221 / 139 = 1
    16'b11011101_10001100 : OUT <= 1;  //221 / 140 = 1
    16'b11011101_10001101 : OUT <= 1;  //221 / 141 = 1
    16'b11011101_10001110 : OUT <= 1;  //221 / 142 = 1
    16'b11011101_10001111 : OUT <= 1;  //221 / 143 = 1
    16'b11011101_10010000 : OUT <= 1;  //221 / 144 = 1
    16'b11011101_10010001 : OUT <= 1;  //221 / 145 = 1
    16'b11011101_10010010 : OUT <= 1;  //221 / 146 = 1
    16'b11011101_10010011 : OUT <= 1;  //221 / 147 = 1
    16'b11011101_10010100 : OUT <= 1;  //221 / 148 = 1
    16'b11011101_10010101 : OUT <= 1;  //221 / 149 = 1
    16'b11011101_10010110 : OUT <= 1;  //221 / 150 = 1
    16'b11011101_10010111 : OUT <= 1;  //221 / 151 = 1
    16'b11011101_10011000 : OUT <= 1;  //221 / 152 = 1
    16'b11011101_10011001 : OUT <= 1;  //221 / 153 = 1
    16'b11011101_10011010 : OUT <= 1;  //221 / 154 = 1
    16'b11011101_10011011 : OUT <= 1;  //221 / 155 = 1
    16'b11011101_10011100 : OUT <= 1;  //221 / 156 = 1
    16'b11011101_10011101 : OUT <= 1;  //221 / 157 = 1
    16'b11011101_10011110 : OUT <= 1;  //221 / 158 = 1
    16'b11011101_10011111 : OUT <= 1;  //221 / 159 = 1
    16'b11011101_10100000 : OUT <= 1;  //221 / 160 = 1
    16'b11011101_10100001 : OUT <= 1;  //221 / 161 = 1
    16'b11011101_10100010 : OUT <= 1;  //221 / 162 = 1
    16'b11011101_10100011 : OUT <= 1;  //221 / 163 = 1
    16'b11011101_10100100 : OUT <= 1;  //221 / 164 = 1
    16'b11011101_10100101 : OUT <= 1;  //221 / 165 = 1
    16'b11011101_10100110 : OUT <= 1;  //221 / 166 = 1
    16'b11011101_10100111 : OUT <= 1;  //221 / 167 = 1
    16'b11011101_10101000 : OUT <= 1;  //221 / 168 = 1
    16'b11011101_10101001 : OUT <= 1;  //221 / 169 = 1
    16'b11011101_10101010 : OUT <= 1;  //221 / 170 = 1
    16'b11011101_10101011 : OUT <= 1;  //221 / 171 = 1
    16'b11011101_10101100 : OUT <= 1;  //221 / 172 = 1
    16'b11011101_10101101 : OUT <= 1;  //221 / 173 = 1
    16'b11011101_10101110 : OUT <= 1;  //221 / 174 = 1
    16'b11011101_10101111 : OUT <= 1;  //221 / 175 = 1
    16'b11011101_10110000 : OUT <= 1;  //221 / 176 = 1
    16'b11011101_10110001 : OUT <= 1;  //221 / 177 = 1
    16'b11011101_10110010 : OUT <= 1;  //221 / 178 = 1
    16'b11011101_10110011 : OUT <= 1;  //221 / 179 = 1
    16'b11011101_10110100 : OUT <= 1;  //221 / 180 = 1
    16'b11011101_10110101 : OUT <= 1;  //221 / 181 = 1
    16'b11011101_10110110 : OUT <= 1;  //221 / 182 = 1
    16'b11011101_10110111 : OUT <= 1;  //221 / 183 = 1
    16'b11011101_10111000 : OUT <= 1;  //221 / 184 = 1
    16'b11011101_10111001 : OUT <= 1;  //221 / 185 = 1
    16'b11011101_10111010 : OUT <= 1;  //221 / 186 = 1
    16'b11011101_10111011 : OUT <= 1;  //221 / 187 = 1
    16'b11011101_10111100 : OUT <= 1;  //221 / 188 = 1
    16'b11011101_10111101 : OUT <= 1;  //221 / 189 = 1
    16'b11011101_10111110 : OUT <= 1;  //221 / 190 = 1
    16'b11011101_10111111 : OUT <= 1;  //221 / 191 = 1
    16'b11011101_11000000 : OUT <= 1;  //221 / 192 = 1
    16'b11011101_11000001 : OUT <= 1;  //221 / 193 = 1
    16'b11011101_11000010 : OUT <= 1;  //221 / 194 = 1
    16'b11011101_11000011 : OUT <= 1;  //221 / 195 = 1
    16'b11011101_11000100 : OUT <= 1;  //221 / 196 = 1
    16'b11011101_11000101 : OUT <= 1;  //221 / 197 = 1
    16'b11011101_11000110 : OUT <= 1;  //221 / 198 = 1
    16'b11011101_11000111 : OUT <= 1;  //221 / 199 = 1
    16'b11011101_11001000 : OUT <= 1;  //221 / 200 = 1
    16'b11011101_11001001 : OUT <= 1;  //221 / 201 = 1
    16'b11011101_11001010 : OUT <= 1;  //221 / 202 = 1
    16'b11011101_11001011 : OUT <= 1;  //221 / 203 = 1
    16'b11011101_11001100 : OUT <= 1;  //221 / 204 = 1
    16'b11011101_11001101 : OUT <= 1;  //221 / 205 = 1
    16'b11011101_11001110 : OUT <= 1;  //221 / 206 = 1
    16'b11011101_11001111 : OUT <= 1;  //221 / 207 = 1
    16'b11011101_11010000 : OUT <= 1;  //221 / 208 = 1
    16'b11011101_11010001 : OUT <= 1;  //221 / 209 = 1
    16'b11011101_11010010 : OUT <= 1;  //221 / 210 = 1
    16'b11011101_11010011 : OUT <= 1;  //221 / 211 = 1
    16'b11011101_11010100 : OUT <= 1;  //221 / 212 = 1
    16'b11011101_11010101 : OUT <= 1;  //221 / 213 = 1
    16'b11011101_11010110 : OUT <= 1;  //221 / 214 = 1
    16'b11011101_11010111 : OUT <= 1;  //221 / 215 = 1
    16'b11011101_11011000 : OUT <= 1;  //221 / 216 = 1
    16'b11011101_11011001 : OUT <= 1;  //221 / 217 = 1
    16'b11011101_11011010 : OUT <= 1;  //221 / 218 = 1
    16'b11011101_11011011 : OUT <= 1;  //221 / 219 = 1
    16'b11011101_11011100 : OUT <= 1;  //221 / 220 = 1
    16'b11011101_11011101 : OUT <= 1;  //221 / 221 = 1
    16'b11011101_11011110 : OUT <= 0;  //221 / 222 = 0
    16'b11011101_11011111 : OUT <= 0;  //221 / 223 = 0
    16'b11011101_11100000 : OUT <= 0;  //221 / 224 = 0
    16'b11011101_11100001 : OUT <= 0;  //221 / 225 = 0
    16'b11011101_11100010 : OUT <= 0;  //221 / 226 = 0
    16'b11011101_11100011 : OUT <= 0;  //221 / 227 = 0
    16'b11011101_11100100 : OUT <= 0;  //221 / 228 = 0
    16'b11011101_11100101 : OUT <= 0;  //221 / 229 = 0
    16'b11011101_11100110 : OUT <= 0;  //221 / 230 = 0
    16'b11011101_11100111 : OUT <= 0;  //221 / 231 = 0
    16'b11011101_11101000 : OUT <= 0;  //221 / 232 = 0
    16'b11011101_11101001 : OUT <= 0;  //221 / 233 = 0
    16'b11011101_11101010 : OUT <= 0;  //221 / 234 = 0
    16'b11011101_11101011 : OUT <= 0;  //221 / 235 = 0
    16'b11011101_11101100 : OUT <= 0;  //221 / 236 = 0
    16'b11011101_11101101 : OUT <= 0;  //221 / 237 = 0
    16'b11011101_11101110 : OUT <= 0;  //221 / 238 = 0
    16'b11011101_11101111 : OUT <= 0;  //221 / 239 = 0
    16'b11011101_11110000 : OUT <= 0;  //221 / 240 = 0
    16'b11011101_11110001 : OUT <= 0;  //221 / 241 = 0
    16'b11011101_11110010 : OUT <= 0;  //221 / 242 = 0
    16'b11011101_11110011 : OUT <= 0;  //221 / 243 = 0
    16'b11011101_11110100 : OUT <= 0;  //221 / 244 = 0
    16'b11011101_11110101 : OUT <= 0;  //221 / 245 = 0
    16'b11011101_11110110 : OUT <= 0;  //221 / 246 = 0
    16'b11011101_11110111 : OUT <= 0;  //221 / 247 = 0
    16'b11011101_11111000 : OUT <= 0;  //221 / 248 = 0
    16'b11011101_11111001 : OUT <= 0;  //221 / 249 = 0
    16'b11011101_11111010 : OUT <= 0;  //221 / 250 = 0
    16'b11011101_11111011 : OUT <= 0;  //221 / 251 = 0
    16'b11011101_11111100 : OUT <= 0;  //221 / 252 = 0
    16'b11011101_11111101 : OUT <= 0;  //221 / 253 = 0
    16'b11011101_11111110 : OUT <= 0;  //221 / 254 = 0
    16'b11011101_11111111 : OUT <= 0;  //221 / 255 = 0
    16'b11011110_00000000 : OUT <= 0;  //222 / 0 = 0
    16'b11011110_00000001 : OUT <= 222;  //222 / 1 = 222
    16'b11011110_00000010 : OUT <= 111;  //222 / 2 = 111
    16'b11011110_00000011 : OUT <= 74;  //222 / 3 = 74
    16'b11011110_00000100 : OUT <= 55;  //222 / 4 = 55
    16'b11011110_00000101 : OUT <= 44;  //222 / 5 = 44
    16'b11011110_00000110 : OUT <= 37;  //222 / 6 = 37
    16'b11011110_00000111 : OUT <= 31;  //222 / 7 = 31
    16'b11011110_00001000 : OUT <= 27;  //222 / 8 = 27
    16'b11011110_00001001 : OUT <= 24;  //222 / 9 = 24
    16'b11011110_00001010 : OUT <= 22;  //222 / 10 = 22
    16'b11011110_00001011 : OUT <= 20;  //222 / 11 = 20
    16'b11011110_00001100 : OUT <= 18;  //222 / 12 = 18
    16'b11011110_00001101 : OUT <= 17;  //222 / 13 = 17
    16'b11011110_00001110 : OUT <= 15;  //222 / 14 = 15
    16'b11011110_00001111 : OUT <= 14;  //222 / 15 = 14
    16'b11011110_00010000 : OUT <= 13;  //222 / 16 = 13
    16'b11011110_00010001 : OUT <= 13;  //222 / 17 = 13
    16'b11011110_00010010 : OUT <= 12;  //222 / 18 = 12
    16'b11011110_00010011 : OUT <= 11;  //222 / 19 = 11
    16'b11011110_00010100 : OUT <= 11;  //222 / 20 = 11
    16'b11011110_00010101 : OUT <= 10;  //222 / 21 = 10
    16'b11011110_00010110 : OUT <= 10;  //222 / 22 = 10
    16'b11011110_00010111 : OUT <= 9;  //222 / 23 = 9
    16'b11011110_00011000 : OUT <= 9;  //222 / 24 = 9
    16'b11011110_00011001 : OUT <= 8;  //222 / 25 = 8
    16'b11011110_00011010 : OUT <= 8;  //222 / 26 = 8
    16'b11011110_00011011 : OUT <= 8;  //222 / 27 = 8
    16'b11011110_00011100 : OUT <= 7;  //222 / 28 = 7
    16'b11011110_00011101 : OUT <= 7;  //222 / 29 = 7
    16'b11011110_00011110 : OUT <= 7;  //222 / 30 = 7
    16'b11011110_00011111 : OUT <= 7;  //222 / 31 = 7
    16'b11011110_00100000 : OUT <= 6;  //222 / 32 = 6
    16'b11011110_00100001 : OUT <= 6;  //222 / 33 = 6
    16'b11011110_00100010 : OUT <= 6;  //222 / 34 = 6
    16'b11011110_00100011 : OUT <= 6;  //222 / 35 = 6
    16'b11011110_00100100 : OUT <= 6;  //222 / 36 = 6
    16'b11011110_00100101 : OUT <= 6;  //222 / 37 = 6
    16'b11011110_00100110 : OUT <= 5;  //222 / 38 = 5
    16'b11011110_00100111 : OUT <= 5;  //222 / 39 = 5
    16'b11011110_00101000 : OUT <= 5;  //222 / 40 = 5
    16'b11011110_00101001 : OUT <= 5;  //222 / 41 = 5
    16'b11011110_00101010 : OUT <= 5;  //222 / 42 = 5
    16'b11011110_00101011 : OUT <= 5;  //222 / 43 = 5
    16'b11011110_00101100 : OUT <= 5;  //222 / 44 = 5
    16'b11011110_00101101 : OUT <= 4;  //222 / 45 = 4
    16'b11011110_00101110 : OUT <= 4;  //222 / 46 = 4
    16'b11011110_00101111 : OUT <= 4;  //222 / 47 = 4
    16'b11011110_00110000 : OUT <= 4;  //222 / 48 = 4
    16'b11011110_00110001 : OUT <= 4;  //222 / 49 = 4
    16'b11011110_00110010 : OUT <= 4;  //222 / 50 = 4
    16'b11011110_00110011 : OUT <= 4;  //222 / 51 = 4
    16'b11011110_00110100 : OUT <= 4;  //222 / 52 = 4
    16'b11011110_00110101 : OUT <= 4;  //222 / 53 = 4
    16'b11011110_00110110 : OUT <= 4;  //222 / 54 = 4
    16'b11011110_00110111 : OUT <= 4;  //222 / 55 = 4
    16'b11011110_00111000 : OUT <= 3;  //222 / 56 = 3
    16'b11011110_00111001 : OUT <= 3;  //222 / 57 = 3
    16'b11011110_00111010 : OUT <= 3;  //222 / 58 = 3
    16'b11011110_00111011 : OUT <= 3;  //222 / 59 = 3
    16'b11011110_00111100 : OUT <= 3;  //222 / 60 = 3
    16'b11011110_00111101 : OUT <= 3;  //222 / 61 = 3
    16'b11011110_00111110 : OUT <= 3;  //222 / 62 = 3
    16'b11011110_00111111 : OUT <= 3;  //222 / 63 = 3
    16'b11011110_01000000 : OUT <= 3;  //222 / 64 = 3
    16'b11011110_01000001 : OUT <= 3;  //222 / 65 = 3
    16'b11011110_01000010 : OUT <= 3;  //222 / 66 = 3
    16'b11011110_01000011 : OUT <= 3;  //222 / 67 = 3
    16'b11011110_01000100 : OUT <= 3;  //222 / 68 = 3
    16'b11011110_01000101 : OUT <= 3;  //222 / 69 = 3
    16'b11011110_01000110 : OUT <= 3;  //222 / 70 = 3
    16'b11011110_01000111 : OUT <= 3;  //222 / 71 = 3
    16'b11011110_01001000 : OUT <= 3;  //222 / 72 = 3
    16'b11011110_01001001 : OUT <= 3;  //222 / 73 = 3
    16'b11011110_01001010 : OUT <= 3;  //222 / 74 = 3
    16'b11011110_01001011 : OUT <= 2;  //222 / 75 = 2
    16'b11011110_01001100 : OUT <= 2;  //222 / 76 = 2
    16'b11011110_01001101 : OUT <= 2;  //222 / 77 = 2
    16'b11011110_01001110 : OUT <= 2;  //222 / 78 = 2
    16'b11011110_01001111 : OUT <= 2;  //222 / 79 = 2
    16'b11011110_01010000 : OUT <= 2;  //222 / 80 = 2
    16'b11011110_01010001 : OUT <= 2;  //222 / 81 = 2
    16'b11011110_01010010 : OUT <= 2;  //222 / 82 = 2
    16'b11011110_01010011 : OUT <= 2;  //222 / 83 = 2
    16'b11011110_01010100 : OUT <= 2;  //222 / 84 = 2
    16'b11011110_01010101 : OUT <= 2;  //222 / 85 = 2
    16'b11011110_01010110 : OUT <= 2;  //222 / 86 = 2
    16'b11011110_01010111 : OUT <= 2;  //222 / 87 = 2
    16'b11011110_01011000 : OUT <= 2;  //222 / 88 = 2
    16'b11011110_01011001 : OUT <= 2;  //222 / 89 = 2
    16'b11011110_01011010 : OUT <= 2;  //222 / 90 = 2
    16'b11011110_01011011 : OUT <= 2;  //222 / 91 = 2
    16'b11011110_01011100 : OUT <= 2;  //222 / 92 = 2
    16'b11011110_01011101 : OUT <= 2;  //222 / 93 = 2
    16'b11011110_01011110 : OUT <= 2;  //222 / 94 = 2
    16'b11011110_01011111 : OUT <= 2;  //222 / 95 = 2
    16'b11011110_01100000 : OUT <= 2;  //222 / 96 = 2
    16'b11011110_01100001 : OUT <= 2;  //222 / 97 = 2
    16'b11011110_01100010 : OUT <= 2;  //222 / 98 = 2
    16'b11011110_01100011 : OUT <= 2;  //222 / 99 = 2
    16'b11011110_01100100 : OUT <= 2;  //222 / 100 = 2
    16'b11011110_01100101 : OUT <= 2;  //222 / 101 = 2
    16'b11011110_01100110 : OUT <= 2;  //222 / 102 = 2
    16'b11011110_01100111 : OUT <= 2;  //222 / 103 = 2
    16'b11011110_01101000 : OUT <= 2;  //222 / 104 = 2
    16'b11011110_01101001 : OUT <= 2;  //222 / 105 = 2
    16'b11011110_01101010 : OUT <= 2;  //222 / 106 = 2
    16'b11011110_01101011 : OUT <= 2;  //222 / 107 = 2
    16'b11011110_01101100 : OUT <= 2;  //222 / 108 = 2
    16'b11011110_01101101 : OUT <= 2;  //222 / 109 = 2
    16'b11011110_01101110 : OUT <= 2;  //222 / 110 = 2
    16'b11011110_01101111 : OUT <= 2;  //222 / 111 = 2
    16'b11011110_01110000 : OUT <= 1;  //222 / 112 = 1
    16'b11011110_01110001 : OUT <= 1;  //222 / 113 = 1
    16'b11011110_01110010 : OUT <= 1;  //222 / 114 = 1
    16'b11011110_01110011 : OUT <= 1;  //222 / 115 = 1
    16'b11011110_01110100 : OUT <= 1;  //222 / 116 = 1
    16'b11011110_01110101 : OUT <= 1;  //222 / 117 = 1
    16'b11011110_01110110 : OUT <= 1;  //222 / 118 = 1
    16'b11011110_01110111 : OUT <= 1;  //222 / 119 = 1
    16'b11011110_01111000 : OUT <= 1;  //222 / 120 = 1
    16'b11011110_01111001 : OUT <= 1;  //222 / 121 = 1
    16'b11011110_01111010 : OUT <= 1;  //222 / 122 = 1
    16'b11011110_01111011 : OUT <= 1;  //222 / 123 = 1
    16'b11011110_01111100 : OUT <= 1;  //222 / 124 = 1
    16'b11011110_01111101 : OUT <= 1;  //222 / 125 = 1
    16'b11011110_01111110 : OUT <= 1;  //222 / 126 = 1
    16'b11011110_01111111 : OUT <= 1;  //222 / 127 = 1
    16'b11011110_10000000 : OUT <= 1;  //222 / 128 = 1
    16'b11011110_10000001 : OUT <= 1;  //222 / 129 = 1
    16'b11011110_10000010 : OUT <= 1;  //222 / 130 = 1
    16'b11011110_10000011 : OUT <= 1;  //222 / 131 = 1
    16'b11011110_10000100 : OUT <= 1;  //222 / 132 = 1
    16'b11011110_10000101 : OUT <= 1;  //222 / 133 = 1
    16'b11011110_10000110 : OUT <= 1;  //222 / 134 = 1
    16'b11011110_10000111 : OUT <= 1;  //222 / 135 = 1
    16'b11011110_10001000 : OUT <= 1;  //222 / 136 = 1
    16'b11011110_10001001 : OUT <= 1;  //222 / 137 = 1
    16'b11011110_10001010 : OUT <= 1;  //222 / 138 = 1
    16'b11011110_10001011 : OUT <= 1;  //222 / 139 = 1
    16'b11011110_10001100 : OUT <= 1;  //222 / 140 = 1
    16'b11011110_10001101 : OUT <= 1;  //222 / 141 = 1
    16'b11011110_10001110 : OUT <= 1;  //222 / 142 = 1
    16'b11011110_10001111 : OUT <= 1;  //222 / 143 = 1
    16'b11011110_10010000 : OUT <= 1;  //222 / 144 = 1
    16'b11011110_10010001 : OUT <= 1;  //222 / 145 = 1
    16'b11011110_10010010 : OUT <= 1;  //222 / 146 = 1
    16'b11011110_10010011 : OUT <= 1;  //222 / 147 = 1
    16'b11011110_10010100 : OUT <= 1;  //222 / 148 = 1
    16'b11011110_10010101 : OUT <= 1;  //222 / 149 = 1
    16'b11011110_10010110 : OUT <= 1;  //222 / 150 = 1
    16'b11011110_10010111 : OUT <= 1;  //222 / 151 = 1
    16'b11011110_10011000 : OUT <= 1;  //222 / 152 = 1
    16'b11011110_10011001 : OUT <= 1;  //222 / 153 = 1
    16'b11011110_10011010 : OUT <= 1;  //222 / 154 = 1
    16'b11011110_10011011 : OUT <= 1;  //222 / 155 = 1
    16'b11011110_10011100 : OUT <= 1;  //222 / 156 = 1
    16'b11011110_10011101 : OUT <= 1;  //222 / 157 = 1
    16'b11011110_10011110 : OUT <= 1;  //222 / 158 = 1
    16'b11011110_10011111 : OUT <= 1;  //222 / 159 = 1
    16'b11011110_10100000 : OUT <= 1;  //222 / 160 = 1
    16'b11011110_10100001 : OUT <= 1;  //222 / 161 = 1
    16'b11011110_10100010 : OUT <= 1;  //222 / 162 = 1
    16'b11011110_10100011 : OUT <= 1;  //222 / 163 = 1
    16'b11011110_10100100 : OUT <= 1;  //222 / 164 = 1
    16'b11011110_10100101 : OUT <= 1;  //222 / 165 = 1
    16'b11011110_10100110 : OUT <= 1;  //222 / 166 = 1
    16'b11011110_10100111 : OUT <= 1;  //222 / 167 = 1
    16'b11011110_10101000 : OUT <= 1;  //222 / 168 = 1
    16'b11011110_10101001 : OUT <= 1;  //222 / 169 = 1
    16'b11011110_10101010 : OUT <= 1;  //222 / 170 = 1
    16'b11011110_10101011 : OUT <= 1;  //222 / 171 = 1
    16'b11011110_10101100 : OUT <= 1;  //222 / 172 = 1
    16'b11011110_10101101 : OUT <= 1;  //222 / 173 = 1
    16'b11011110_10101110 : OUT <= 1;  //222 / 174 = 1
    16'b11011110_10101111 : OUT <= 1;  //222 / 175 = 1
    16'b11011110_10110000 : OUT <= 1;  //222 / 176 = 1
    16'b11011110_10110001 : OUT <= 1;  //222 / 177 = 1
    16'b11011110_10110010 : OUT <= 1;  //222 / 178 = 1
    16'b11011110_10110011 : OUT <= 1;  //222 / 179 = 1
    16'b11011110_10110100 : OUT <= 1;  //222 / 180 = 1
    16'b11011110_10110101 : OUT <= 1;  //222 / 181 = 1
    16'b11011110_10110110 : OUT <= 1;  //222 / 182 = 1
    16'b11011110_10110111 : OUT <= 1;  //222 / 183 = 1
    16'b11011110_10111000 : OUT <= 1;  //222 / 184 = 1
    16'b11011110_10111001 : OUT <= 1;  //222 / 185 = 1
    16'b11011110_10111010 : OUT <= 1;  //222 / 186 = 1
    16'b11011110_10111011 : OUT <= 1;  //222 / 187 = 1
    16'b11011110_10111100 : OUT <= 1;  //222 / 188 = 1
    16'b11011110_10111101 : OUT <= 1;  //222 / 189 = 1
    16'b11011110_10111110 : OUT <= 1;  //222 / 190 = 1
    16'b11011110_10111111 : OUT <= 1;  //222 / 191 = 1
    16'b11011110_11000000 : OUT <= 1;  //222 / 192 = 1
    16'b11011110_11000001 : OUT <= 1;  //222 / 193 = 1
    16'b11011110_11000010 : OUT <= 1;  //222 / 194 = 1
    16'b11011110_11000011 : OUT <= 1;  //222 / 195 = 1
    16'b11011110_11000100 : OUT <= 1;  //222 / 196 = 1
    16'b11011110_11000101 : OUT <= 1;  //222 / 197 = 1
    16'b11011110_11000110 : OUT <= 1;  //222 / 198 = 1
    16'b11011110_11000111 : OUT <= 1;  //222 / 199 = 1
    16'b11011110_11001000 : OUT <= 1;  //222 / 200 = 1
    16'b11011110_11001001 : OUT <= 1;  //222 / 201 = 1
    16'b11011110_11001010 : OUT <= 1;  //222 / 202 = 1
    16'b11011110_11001011 : OUT <= 1;  //222 / 203 = 1
    16'b11011110_11001100 : OUT <= 1;  //222 / 204 = 1
    16'b11011110_11001101 : OUT <= 1;  //222 / 205 = 1
    16'b11011110_11001110 : OUT <= 1;  //222 / 206 = 1
    16'b11011110_11001111 : OUT <= 1;  //222 / 207 = 1
    16'b11011110_11010000 : OUT <= 1;  //222 / 208 = 1
    16'b11011110_11010001 : OUT <= 1;  //222 / 209 = 1
    16'b11011110_11010010 : OUT <= 1;  //222 / 210 = 1
    16'b11011110_11010011 : OUT <= 1;  //222 / 211 = 1
    16'b11011110_11010100 : OUT <= 1;  //222 / 212 = 1
    16'b11011110_11010101 : OUT <= 1;  //222 / 213 = 1
    16'b11011110_11010110 : OUT <= 1;  //222 / 214 = 1
    16'b11011110_11010111 : OUT <= 1;  //222 / 215 = 1
    16'b11011110_11011000 : OUT <= 1;  //222 / 216 = 1
    16'b11011110_11011001 : OUT <= 1;  //222 / 217 = 1
    16'b11011110_11011010 : OUT <= 1;  //222 / 218 = 1
    16'b11011110_11011011 : OUT <= 1;  //222 / 219 = 1
    16'b11011110_11011100 : OUT <= 1;  //222 / 220 = 1
    16'b11011110_11011101 : OUT <= 1;  //222 / 221 = 1
    16'b11011110_11011110 : OUT <= 1;  //222 / 222 = 1
    16'b11011110_11011111 : OUT <= 0;  //222 / 223 = 0
    16'b11011110_11100000 : OUT <= 0;  //222 / 224 = 0
    16'b11011110_11100001 : OUT <= 0;  //222 / 225 = 0
    16'b11011110_11100010 : OUT <= 0;  //222 / 226 = 0
    16'b11011110_11100011 : OUT <= 0;  //222 / 227 = 0
    16'b11011110_11100100 : OUT <= 0;  //222 / 228 = 0
    16'b11011110_11100101 : OUT <= 0;  //222 / 229 = 0
    16'b11011110_11100110 : OUT <= 0;  //222 / 230 = 0
    16'b11011110_11100111 : OUT <= 0;  //222 / 231 = 0
    16'b11011110_11101000 : OUT <= 0;  //222 / 232 = 0
    16'b11011110_11101001 : OUT <= 0;  //222 / 233 = 0
    16'b11011110_11101010 : OUT <= 0;  //222 / 234 = 0
    16'b11011110_11101011 : OUT <= 0;  //222 / 235 = 0
    16'b11011110_11101100 : OUT <= 0;  //222 / 236 = 0
    16'b11011110_11101101 : OUT <= 0;  //222 / 237 = 0
    16'b11011110_11101110 : OUT <= 0;  //222 / 238 = 0
    16'b11011110_11101111 : OUT <= 0;  //222 / 239 = 0
    16'b11011110_11110000 : OUT <= 0;  //222 / 240 = 0
    16'b11011110_11110001 : OUT <= 0;  //222 / 241 = 0
    16'b11011110_11110010 : OUT <= 0;  //222 / 242 = 0
    16'b11011110_11110011 : OUT <= 0;  //222 / 243 = 0
    16'b11011110_11110100 : OUT <= 0;  //222 / 244 = 0
    16'b11011110_11110101 : OUT <= 0;  //222 / 245 = 0
    16'b11011110_11110110 : OUT <= 0;  //222 / 246 = 0
    16'b11011110_11110111 : OUT <= 0;  //222 / 247 = 0
    16'b11011110_11111000 : OUT <= 0;  //222 / 248 = 0
    16'b11011110_11111001 : OUT <= 0;  //222 / 249 = 0
    16'b11011110_11111010 : OUT <= 0;  //222 / 250 = 0
    16'b11011110_11111011 : OUT <= 0;  //222 / 251 = 0
    16'b11011110_11111100 : OUT <= 0;  //222 / 252 = 0
    16'b11011110_11111101 : OUT <= 0;  //222 / 253 = 0
    16'b11011110_11111110 : OUT <= 0;  //222 / 254 = 0
    16'b11011110_11111111 : OUT <= 0;  //222 / 255 = 0
    16'b11011111_00000000 : OUT <= 0;  //223 / 0 = 0
    16'b11011111_00000001 : OUT <= 223;  //223 / 1 = 223
    16'b11011111_00000010 : OUT <= 111;  //223 / 2 = 111
    16'b11011111_00000011 : OUT <= 74;  //223 / 3 = 74
    16'b11011111_00000100 : OUT <= 55;  //223 / 4 = 55
    16'b11011111_00000101 : OUT <= 44;  //223 / 5 = 44
    16'b11011111_00000110 : OUT <= 37;  //223 / 6 = 37
    16'b11011111_00000111 : OUT <= 31;  //223 / 7 = 31
    16'b11011111_00001000 : OUT <= 27;  //223 / 8 = 27
    16'b11011111_00001001 : OUT <= 24;  //223 / 9 = 24
    16'b11011111_00001010 : OUT <= 22;  //223 / 10 = 22
    16'b11011111_00001011 : OUT <= 20;  //223 / 11 = 20
    16'b11011111_00001100 : OUT <= 18;  //223 / 12 = 18
    16'b11011111_00001101 : OUT <= 17;  //223 / 13 = 17
    16'b11011111_00001110 : OUT <= 15;  //223 / 14 = 15
    16'b11011111_00001111 : OUT <= 14;  //223 / 15 = 14
    16'b11011111_00010000 : OUT <= 13;  //223 / 16 = 13
    16'b11011111_00010001 : OUT <= 13;  //223 / 17 = 13
    16'b11011111_00010010 : OUT <= 12;  //223 / 18 = 12
    16'b11011111_00010011 : OUT <= 11;  //223 / 19 = 11
    16'b11011111_00010100 : OUT <= 11;  //223 / 20 = 11
    16'b11011111_00010101 : OUT <= 10;  //223 / 21 = 10
    16'b11011111_00010110 : OUT <= 10;  //223 / 22 = 10
    16'b11011111_00010111 : OUT <= 9;  //223 / 23 = 9
    16'b11011111_00011000 : OUT <= 9;  //223 / 24 = 9
    16'b11011111_00011001 : OUT <= 8;  //223 / 25 = 8
    16'b11011111_00011010 : OUT <= 8;  //223 / 26 = 8
    16'b11011111_00011011 : OUT <= 8;  //223 / 27 = 8
    16'b11011111_00011100 : OUT <= 7;  //223 / 28 = 7
    16'b11011111_00011101 : OUT <= 7;  //223 / 29 = 7
    16'b11011111_00011110 : OUT <= 7;  //223 / 30 = 7
    16'b11011111_00011111 : OUT <= 7;  //223 / 31 = 7
    16'b11011111_00100000 : OUT <= 6;  //223 / 32 = 6
    16'b11011111_00100001 : OUT <= 6;  //223 / 33 = 6
    16'b11011111_00100010 : OUT <= 6;  //223 / 34 = 6
    16'b11011111_00100011 : OUT <= 6;  //223 / 35 = 6
    16'b11011111_00100100 : OUT <= 6;  //223 / 36 = 6
    16'b11011111_00100101 : OUT <= 6;  //223 / 37 = 6
    16'b11011111_00100110 : OUT <= 5;  //223 / 38 = 5
    16'b11011111_00100111 : OUT <= 5;  //223 / 39 = 5
    16'b11011111_00101000 : OUT <= 5;  //223 / 40 = 5
    16'b11011111_00101001 : OUT <= 5;  //223 / 41 = 5
    16'b11011111_00101010 : OUT <= 5;  //223 / 42 = 5
    16'b11011111_00101011 : OUT <= 5;  //223 / 43 = 5
    16'b11011111_00101100 : OUT <= 5;  //223 / 44 = 5
    16'b11011111_00101101 : OUT <= 4;  //223 / 45 = 4
    16'b11011111_00101110 : OUT <= 4;  //223 / 46 = 4
    16'b11011111_00101111 : OUT <= 4;  //223 / 47 = 4
    16'b11011111_00110000 : OUT <= 4;  //223 / 48 = 4
    16'b11011111_00110001 : OUT <= 4;  //223 / 49 = 4
    16'b11011111_00110010 : OUT <= 4;  //223 / 50 = 4
    16'b11011111_00110011 : OUT <= 4;  //223 / 51 = 4
    16'b11011111_00110100 : OUT <= 4;  //223 / 52 = 4
    16'b11011111_00110101 : OUT <= 4;  //223 / 53 = 4
    16'b11011111_00110110 : OUT <= 4;  //223 / 54 = 4
    16'b11011111_00110111 : OUT <= 4;  //223 / 55 = 4
    16'b11011111_00111000 : OUT <= 3;  //223 / 56 = 3
    16'b11011111_00111001 : OUT <= 3;  //223 / 57 = 3
    16'b11011111_00111010 : OUT <= 3;  //223 / 58 = 3
    16'b11011111_00111011 : OUT <= 3;  //223 / 59 = 3
    16'b11011111_00111100 : OUT <= 3;  //223 / 60 = 3
    16'b11011111_00111101 : OUT <= 3;  //223 / 61 = 3
    16'b11011111_00111110 : OUT <= 3;  //223 / 62 = 3
    16'b11011111_00111111 : OUT <= 3;  //223 / 63 = 3
    16'b11011111_01000000 : OUT <= 3;  //223 / 64 = 3
    16'b11011111_01000001 : OUT <= 3;  //223 / 65 = 3
    16'b11011111_01000010 : OUT <= 3;  //223 / 66 = 3
    16'b11011111_01000011 : OUT <= 3;  //223 / 67 = 3
    16'b11011111_01000100 : OUT <= 3;  //223 / 68 = 3
    16'b11011111_01000101 : OUT <= 3;  //223 / 69 = 3
    16'b11011111_01000110 : OUT <= 3;  //223 / 70 = 3
    16'b11011111_01000111 : OUT <= 3;  //223 / 71 = 3
    16'b11011111_01001000 : OUT <= 3;  //223 / 72 = 3
    16'b11011111_01001001 : OUT <= 3;  //223 / 73 = 3
    16'b11011111_01001010 : OUT <= 3;  //223 / 74 = 3
    16'b11011111_01001011 : OUT <= 2;  //223 / 75 = 2
    16'b11011111_01001100 : OUT <= 2;  //223 / 76 = 2
    16'b11011111_01001101 : OUT <= 2;  //223 / 77 = 2
    16'b11011111_01001110 : OUT <= 2;  //223 / 78 = 2
    16'b11011111_01001111 : OUT <= 2;  //223 / 79 = 2
    16'b11011111_01010000 : OUT <= 2;  //223 / 80 = 2
    16'b11011111_01010001 : OUT <= 2;  //223 / 81 = 2
    16'b11011111_01010010 : OUT <= 2;  //223 / 82 = 2
    16'b11011111_01010011 : OUT <= 2;  //223 / 83 = 2
    16'b11011111_01010100 : OUT <= 2;  //223 / 84 = 2
    16'b11011111_01010101 : OUT <= 2;  //223 / 85 = 2
    16'b11011111_01010110 : OUT <= 2;  //223 / 86 = 2
    16'b11011111_01010111 : OUT <= 2;  //223 / 87 = 2
    16'b11011111_01011000 : OUT <= 2;  //223 / 88 = 2
    16'b11011111_01011001 : OUT <= 2;  //223 / 89 = 2
    16'b11011111_01011010 : OUT <= 2;  //223 / 90 = 2
    16'b11011111_01011011 : OUT <= 2;  //223 / 91 = 2
    16'b11011111_01011100 : OUT <= 2;  //223 / 92 = 2
    16'b11011111_01011101 : OUT <= 2;  //223 / 93 = 2
    16'b11011111_01011110 : OUT <= 2;  //223 / 94 = 2
    16'b11011111_01011111 : OUT <= 2;  //223 / 95 = 2
    16'b11011111_01100000 : OUT <= 2;  //223 / 96 = 2
    16'b11011111_01100001 : OUT <= 2;  //223 / 97 = 2
    16'b11011111_01100010 : OUT <= 2;  //223 / 98 = 2
    16'b11011111_01100011 : OUT <= 2;  //223 / 99 = 2
    16'b11011111_01100100 : OUT <= 2;  //223 / 100 = 2
    16'b11011111_01100101 : OUT <= 2;  //223 / 101 = 2
    16'b11011111_01100110 : OUT <= 2;  //223 / 102 = 2
    16'b11011111_01100111 : OUT <= 2;  //223 / 103 = 2
    16'b11011111_01101000 : OUT <= 2;  //223 / 104 = 2
    16'b11011111_01101001 : OUT <= 2;  //223 / 105 = 2
    16'b11011111_01101010 : OUT <= 2;  //223 / 106 = 2
    16'b11011111_01101011 : OUT <= 2;  //223 / 107 = 2
    16'b11011111_01101100 : OUT <= 2;  //223 / 108 = 2
    16'b11011111_01101101 : OUT <= 2;  //223 / 109 = 2
    16'b11011111_01101110 : OUT <= 2;  //223 / 110 = 2
    16'b11011111_01101111 : OUT <= 2;  //223 / 111 = 2
    16'b11011111_01110000 : OUT <= 1;  //223 / 112 = 1
    16'b11011111_01110001 : OUT <= 1;  //223 / 113 = 1
    16'b11011111_01110010 : OUT <= 1;  //223 / 114 = 1
    16'b11011111_01110011 : OUT <= 1;  //223 / 115 = 1
    16'b11011111_01110100 : OUT <= 1;  //223 / 116 = 1
    16'b11011111_01110101 : OUT <= 1;  //223 / 117 = 1
    16'b11011111_01110110 : OUT <= 1;  //223 / 118 = 1
    16'b11011111_01110111 : OUT <= 1;  //223 / 119 = 1
    16'b11011111_01111000 : OUT <= 1;  //223 / 120 = 1
    16'b11011111_01111001 : OUT <= 1;  //223 / 121 = 1
    16'b11011111_01111010 : OUT <= 1;  //223 / 122 = 1
    16'b11011111_01111011 : OUT <= 1;  //223 / 123 = 1
    16'b11011111_01111100 : OUT <= 1;  //223 / 124 = 1
    16'b11011111_01111101 : OUT <= 1;  //223 / 125 = 1
    16'b11011111_01111110 : OUT <= 1;  //223 / 126 = 1
    16'b11011111_01111111 : OUT <= 1;  //223 / 127 = 1
    16'b11011111_10000000 : OUT <= 1;  //223 / 128 = 1
    16'b11011111_10000001 : OUT <= 1;  //223 / 129 = 1
    16'b11011111_10000010 : OUT <= 1;  //223 / 130 = 1
    16'b11011111_10000011 : OUT <= 1;  //223 / 131 = 1
    16'b11011111_10000100 : OUT <= 1;  //223 / 132 = 1
    16'b11011111_10000101 : OUT <= 1;  //223 / 133 = 1
    16'b11011111_10000110 : OUT <= 1;  //223 / 134 = 1
    16'b11011111_10000111 : OUT <= 1;  //223 / 135 = 1
    16'b11011111_10001000 : OUT <= 1;  //223 / 136 = 1
    16'b11011111_10001001 : OUT <= 1;  //223 / 137 = 1
    16'b11011111_10001010 : OUT <= 1;  //223 / 138 = 1
    16'b11011111_10001011 : OUT <= 1;  //223 / 139 = 1
    16'b11011111_10001100 : OUT <= 1;  //223 / 140 = 1
    16'b11011111_10001101 : OUT <= 1;  //223 / 141 = 1
    16'b11011111_10001110 : OUT <= 1;  //223 / 142 = 1
    16'b11011111_10001111 : OUT <= 1;  //223 / 143 = 1
    16'b11011111_10010000 : OUT <= 1;  //223 / 144 = 1
    16'b11011111_10010001 : OUT <= 1;  //223 / 145 = 1
    16'b11011111_10010010 : OUT <= 1;  //223 / 146 = 1
    16'b11011111_10010011 : OUT <= 1;  //223 / 147 = 1
    16'b11011111_10010100 : OUT <= 1;  //223 / 148 = 1
    16'b11011111_10010101 : OUT <= 1;  //223 / 149 = 1
    16'b11011111_10010110 : OUT <= 1;  //223 / 150 = 1
    16'b11011111_10010111 : OUT <= 1;  //223 / 151 = 1
    16'b11011111_10011000 : OUT <= 1;  //223 / 152 = 1
    16'b11011111_10011001 : OUT <= 1;  //223 / 153 = 1
    16'b11011111_10011010 : OUT <= 1;  //223 / 154 = 1
    16'b11011111_10011011 : OUT <= 1;  //223 / 155 = 1
    16'b11011111_10011100 : OUT <= 1;  //223 / 156 = 1
    16'b11011111_10011101 : OUT <= 1;  //223 / 157 = 1
    16'b11011111_10011110 : OUT <= 1;  //223 / 158 = 1
    16'b11011111_10011111 : OUT <= 1;  //223 / 159 = 1
    16'b11011111_10100000 : OUT <= 1;  //223 / 160 = 1
    16'b11011111_10100001 : OUT <= 1;  //223 / 161 = 1
    16'b11011111_10100010 : OUT <= 1;  //223 / 162 = 1
    16'b11011111_10100011 : OUT <= 1;  //223 / 163 = 1
    16'b11011111_10100100 : OUT <= 1;  //223 / 164 = 1
    16'b11011111_10100101 : OUT <= 1;  //223 / 165 = 1
    16'b11011111_10100110 : OUT <= 1;  //223 / 166 = 1
    16'b11011111_10100111 : OUT <= 1;  //223 / 167 = 1
    16'b11011111_10101000 : OUT <= 1;  //223 / 168 = 1
    16'b11011111_10101001 : OUT <= 1;  //223 / 169 = 1
    16'b11011111_10101010 : OUT <= 1;  //223 / 170 = 1
    16'b11011111_10101011 : OUT <= 1;  //223 / 171 = 1
    16'b11011111_10101100 : OUT <= 1;  //223 / 172 = 1
    16'b11011111_10101101 : OUT <= 1;  //223 / 173 = 1
    16'b11011111_10101110 : OUT <= 1;  //223 / 174 = 1
    16'b11011111_10101111 : OUT <= 1;  //223 / 175 = 1
    16'b11011111_10110000 : OUT <= 1;  //223 / 176 = 1
    16'b11011111_10110001 : OUT <= 1;  //223 / 177 = 1
    16'b11011111_10110010 : OUT <= 1;  //223 / 178 = 1
    16'b11011111_10110011 : OUT <= 1;  //223 / 179 = 1
    16'b11011111_10110100 : OUT <= 1;  //223 / 180 = 1
    16'b11011111_10110101 : OUT <= 1;  //223 / 181 = 1
    16'b11011111_10110110 : OUT <= 1;  //223 / 182 = 1
    16'b11011111_10110111 : OUT <= 1;  //223 / 183 = 1
    16'b11011111_10111000 : OUT <= 1;  //223 / 184 = 1
    16'b11011111_10111001 : OUT <= 1;  //223 / 185 = 1
    16'b11011111_10111010 : OUT <= 1;  //223 / 186 = 1
    16'b11011111_10111011 : OUT <= 1;  //223 / 187 = 1
    16'b11011111_10111100 : OUT <= 1;  //223 / 188 = 1
    16'b11011111_10111101 : OUT <= 1;  //223 / 189 = 1
    16'b11011111_10111110 : OUT <= 1;  //223 / 190 = 1
    16'b11011111_10111111 : OUT <= 1;  //223 / 191 = 1
    16'b11011111_11000000 : OUT <= 1;  //223 / 192 = 1
    16'b11011111_11000001 : OUT <= 1;  //223 / 193 = 1
    16'b11011111_11000010 : OUT <= 1;  //223 / 194 = 1
    16'b11011111_11000011 : OUT <= 1;  //223 / 195 = 1
    16'b11011111_11000100 : OUT <= 1;  //223 / 196 = 1
    16'b11011111_11000101 : OUT <= 1;  //223 / 197 = 1
    16'b11011111_11000110 : OUT <= 1;  //223 / 198 = 1
    16'b11011111_11000111 : OUT <= 1;  //223 / 199 = 1
    16'b11011111_11001000 : OUT <= 1;  //223 / 200 = 1
    16'b11011111_11001001 : OUT <= 1;  //223 / 201 = 1
    16'b11011111_11001010 : OUT <= 1;  //223 / 202 = 1
    16'b11011111_11001011 : OUT <= 1;  //223 / 203 = 1
    16'b11011111_11001100 : OUT <= 1;  //223 / 204 = 1
    16'b11011111_11001101 : OUT <= 1;  //223 / 205 = 1
    16'b11011111_11001110 : OUT <= 1;  //223 / 206 = 1
    16'b11011111_11001111 : OUT <= 1;  //223 / 207 = 1
    16'b11011111_11010000 : OUT <= 1;  //223 / 208 = 1
    16'b11011111_11010001 : OUT <= 1;  //223 / 209 = 1
    16'b11011111_11010010 : OUT <= 1;  //223 / 210 = 1
    16'b11011111_11010011 : OUT <= 1;  //223 / 211 = 1
    16'b11011111_11010100 : OUT <= 1;  //223 / 212 = 1
    16'b11011111_11010101 : OUT <= 1;  //223 / 213 = 1
    16'b11011111_11010110 : OUT <= 1;  //223 / 214 = 1
    16'b11011111_11010111 : OUT <= 1;  //223 / 215 = 1
    16'b11011111_11011000 : OUT <= 1;  //223 / 216 = 1
    16'b11011111_11011001 : OUT <= 1;  //223 / 217 = 1
    16'b11011111_11011010 : OUT <= 1;  //223 / 218 = 1
    16'b11011111_11011011 : OUT <= 1;  //223 / 219 = 1
    16'b11011111_11011100 : OUT <= 1;  //223 / 220 = 1
    16'b11011111_11011101 : OUT <= 1;  //223 / 221 = 1
    16'b11011111_11011110 : OUT <= 1;  //223 / 222 = 1
    16'b11011111_11011111 : OUT <= 1;  //223 / 223 = 1
    16'b11011111_11100000 : OUT <= 0;  //223 / 224 = 0
    16'b11011111_11100001 : OUT <= 0;  //223 / 225 = 0
    16'b11011111_11100010 : OUT <= 0;  //223 / 226 = 0
    16'b11011111_11100011 : OUT <= 0;  //223 / 227 = 0
    16'b11011111_11100100 : OUT <= 0;  //223 / 228 = 0
    16'b11011111_11100101 : OUT <= 0;  //223 / 229 = 0
    16'b11011111_11100110 : OUT <= 0;  //223 / 230 = 0
    16'b11011111_11100111 : OUT <= 0;  //223 / 231 = 0
    16'b11011111_11101000 : OUT <= 0;  //223 / 232 = 0
    16'b11011111_11101001 : OUT <= 0;  //223 / 233 = 0
    16'b11011111_11101010 : OUT <= 0;  //223 / 234 = 0
    16'b11011111_11101011 : OUT <= 0;  //223 / 235 = 0
    16'b11011111_11101100 : OUT <= 0;  //223 / 236 = 0
    16'b11011111_11101101 : OUT <= 0;  //223 / 237 = 0
    16'b11011111_11101110 : OUT <= 0;  //223 / 238 = 0
    16'b11011111_11101111 : OUT <= 0;  //223 / 239 = 0
    16'b11011111_11110000 : OUT <= 0;  //223 / 240 = 0
    16'b11011111_11110001 : OUT <= 0;  //223 / 241 = 0
    16'b11011111_11110010 : OUT <= 0;  //223 / 242 = 0
    16'b11011111_11110011 : OUT <= 0;  //223 / 243 = 0
    16'b11011111_11110100 : OUT <= 0;  //223 / 244 = 0
    16'b11011111_11110101 : OUT <= 0;  //223 / 245 = 0
    16'b11011111_11110110 : OUT <= 0;  //223 / 246 = 0
    16'b11011111_11110111 : OUT <= 0;  //223 / 247 = 0
    16'b11011111_11111000 : OUT <= 0;  //223 / 248 = 0
    16'b11011111_11111001 : OUT <= 0;  //223 / 249 = 0
    16'b11011111_11111010 : OUT <= 0;  //223 / 250 = 0
    16'b11011111_11111011 : OUT <= 0;  //223 / 251 = 0
    16'b11011111_11111100 : OUT <= 0;  //223 / 252 = 0
    16'b11011111_11111101 : OUT <= 0;  //223 / 253 = 0
    16'b11011111_11111110 : OUT <= 0;  //223 / 254 = 0
    16'b11011111_11111111 : OUT <= 0;  //223 / 255 = 0
    16'b11100000_00000000 : OUT <= 0;  //224 / 0 = 0
    16'b11100000_00000001 : OUT <= 224;  //224 / 1 = 224
    16'b11100000_00000010 : OUT <= 112;  //224 / 2 = 112
    16'b11100000_00000011 : OUT <= 74;  //224 / 3 = 74
    16'b11100000_00000100 : OUT <= 56;  //224 / 4 = 56
    16'b11100000_00000101 : OUT <= 44;  //224 / 5 = 44
    16'b11100000_00000110 : OUT <= 37;  //224 / 6 = 37
    16'b11100000_00000111 : OUT <= 32;  //224 / 7 = 32
    16'b11100000_00001000 : OUT <= 28;  //224 / 8 = 28
    16'b11100000_00001001 : OUT <= 24;  //224 / 9 = 24
    16'b11100000_00001010 : OUT <= 22;  //224 / 10 = 22
    16'b11100000_00001011 : OUT <= 20;  //224 / 11 = 20
    16'b11100000_00001100 : OUT <= 18;  //224 / 12 = 18
    16'b11100000_00001101 : OUT <= 17;  //224 / 13 = 17
    16'b11100000_00001110 : OUT <= 16;  //224 / 14 = 16
    16'b11100000_00001111 : OUT <= 14;  //224 / 15 = 14
    16'b11100000_00010000 : OUT <= 14;  //224 / 16 = 14
    16'b11100000_00010001 : OUT <= 13;  //224 / 17 = 13
    16'b11100000_00010010 : OUT <= 12;  //224 / 18 = 12
    16'b11100000_00010011 : OUT <= 11;  //224 / 19 = 11
    16'b11100000_00010100 : OUT <= 11;  //224 / 20 = 11
    16'b11100000_00010101 : OUT <= 10;  //224 / 21 = 10
    16'b11100000_00010110 : OUT <= 10;  //224 / 22 = 10
    16'b11100000_00010111 : OUT <= 9;  //224 / 23 = 9
    16'b11100000_00011000 : OUT <= 9;  //224 / 24 = 9
    16'b11100000_00011001 : OUT <= 8;  //224 / 25 = 8
    16'b11100000_00011010 : OUT <= 8;  //224 / 26 = 8
    16'b11100000_00011011 : OUT <= 8;  //224 / 27 = 8
    16'b11100000_00011100 : OUT <= 8;  //224 / 28 = 8
    16'b11100000_00011101 : OUT <= 7;  //224 / 29 = 7
    16'b11100000_00011110 : OUT <= 7;  //224 / 30 = 7
    16'b11100000_00011111 : OUT <= 7;  //224 / 31 = 7
    16'b11100000_00100000 : OUT <= 7;  //224 / 32 = 7
    16'b11100000_00100001 : OUT <= 6;  //224 / 33 = 6
    16'b11100000_00100010 : OUT <= 6;  //224 / 34 = 6
    16'b11100000_00100011 : OUT <= 6;  //224 / 35 = 6
    16'b11100000_00100100 : OUT <= 6;  //224 / 36 = 6
    16'b11100000_00100101 : OUT <= 6;  //224 / 37 = 6
    16'b11100000_00100110 : OUT <= 5;  //224 / 38 = 5
    16'b11100000_00100111 : OUT <= 5;  //224 / 39 = 5
    16'b11100000_00101000 : OUT <= 5;  //224 / 40 = 5
    16'b11100000_00101001 : OUT <= 5;  //224 / 41 = 5
    16'b11100000_00101010 : OUT <= 5;  //224 / 42 = 5
    16'b11100000_00101011 : OUT <= 5;  //224 / 43 = 5
    16'b11100000_00101100 : OUT <= 5;  //224 / 44 = 5
    16'b11100000_00101101 : OUT <= 4;  //224 / 45 = 4
    16'b11100000_00101110 : OUT <= 4;  //224 / 46 = 4
    16'b11100000_00101111 : OUT <= 4;  //224 / 47 = 4
    16'b11100000_00110000 : OUT <= 4;  //224 / 48 = 4
    16'b11100000_00110001 : OUT <= 4;  //224 / 49 = 4
    16'b11100000_00110010 : OUT <= 4;  //224 / 50 = 4
    16'b11100000_00110011 : OUT <= 4;  //224 / 51 = 4
    16'b11100000_00110100 : OUT <= 4;  //224 / 52 = 4
    16'b11100000_00110101 : OUT <= 4;  //224 / 53 = 4
    16'b11100000_00110110 : OUT <= 4;  //224 / 54 = 4
    16'b11100000_00110111 : OUT <= 4;  //224 / 55 = 4
    16'b11100000_00111000 : OUT <= 4;  //224 / 56 = 4
    16'b11100000_00111001 : OUT <= 3;  //224 / 57 = 3
    16'b11100000_00111010 : OUT <= 3;  //224 / 58 = 3
    16'b11100000_00111011 : OUT <= 3;  //224 / 59 = 3
    16'b11100000_00111100 : OUT <= 3;  //224 / 60 = 3
    16'b11100000_00111101 : OUT <= 3;  //224 / 61 = 3
    16'b11100000_00111110 : OUT <= 3;  //224 / 62 = 3
    16'b11100000_00111111 : OUT <= 3;  //224 / 63 = 3
    16'b11100000_01000000 : OUT <= 3;  //224 / 64 = 3
    16'b11100000_01000001 : OUT <= 3;  //224 / 65 = 3
    16'b11100000_01000010 : OUT <= 3;  //224 / 66 = 3
    16'b11100000_01000011 : OUT <= 3;  //224 / 67 = 3
    16'b11100000_01000100 : OUT <= 3;  //224 / 68 = 3
    16'b11100000_01000101 : OUT <= 3;  //224 / 69 = 3
    16'b11100000_01000110 : OUT <= 3;  //224 / 70 = 3
    16'b11100000_01000111 : OUT <= 3;  //224 / 71 = 3
    16'b11100000_01001000 : OUT <= 3;  //224 / 72 = 3
    16'b11100000_01001001 : OUT <= 3;  //224 / 73 = 3
    16'b11100000_01001010 : OUT <= 3;  //224 / 74 = 3
    16'b11100000_01001011 : OUT <= 2;  //224 / 75 = 2
    16'b11100000_01001100 : OUT <= 2;  //224 / 76 = 2
    16'b11100000_01001101 : OUT <= 2;  //224 / 77 = 2
    16'b11100000_01001110 : OUT <= 2;  //224 / 78 = 2
    16'b11100000_01001111 : OUT <= 2;  //224 / 79 = 2
    16'b11100000_01010000 : OUT <= 2;  //224 / 80 = 2
    16'b11100000_01010001 : OUT <= 2;  //224 / 81 = 2
    16'b11100000_01010010 : OUT <= 2;  //224 / 82 = 2
    16'b11100000_01010011 : OUT <= 2;  //224 / 83 = 2
    16'b11100000_01010100 : OUT <= 2;  //224 / 84 = 2
    16'b11100000_01010101 : OUT <= 2;  //224 / 85 = 2
    16'b11100000_01010110 : OUT <= 2;  //224 / 86 = 2
    16'b11100000_01010111 : OUT <= 2;  //224 / 87 = 2
    16'b11100000_01011000 : OUT <= 2;  //224 / 88 = 2
    16'b11100000_01011001 : OUT <= 2;  //224 / 89 = 2
    16'b11100000_01011010 : OUT <= 2;  //224 / 90 = 2
    16'b11100000_01011011 : OUT <= 2;  //224 / 91 = 2
    16'b11100000_01011100 : OUT <= 2;  //224 / 92 = 2
    16'b11100000_01011101 : OUT <= 2;  //224 / 93 = 2
    16'b11100000_01011110 : OUT <= 2;  //224 / 94 = 2
    16'b11100000_01011111 : OUT <= 2;  //224 / 95 = 2
    16'b11100000_01100000 : OUT <= 2;  //224 / 96 = 2
    16'b11100000_01100001 : OUT <= 2;  //224 / 97 = 2
    16'b11100000_01100010 : OUT <= 2;  //224 / 98 = 2
    16'b11100000_01100011 : OUT <= 2;  //224 / 99 = 2
    16'b11100000_01100100 : OUT <= 2;  //224 / 100 = 2
    16'b11100000_01100101 : OUT <= 2;  //224 / 101 = 2
    16'b11100000_01100110 : OUT <= 2;  //224 / 102 = 2
    16'b11100000_01100111 : OUT <= 2;  //224 / 103 = 2
    16'b11100000_01101000 : OUT <= 2;  //224 / 104 = 2
    16'b11100000_01101001 : OUT <= 2;  //224 / 105 = 2
    16'b11100000_01101010 : OUT <= 2;  //224 / 106 = 2
    16'b11100000_01101011 : OUT <= 2;  //224 / 107 = 2
    16'b11100000_01101100 : OUT <= 2;  //224 / 108 = 2
    16'b11100000_01101101 : OUT <= 2;  //224 / 109 = 2
    16'b11100000_01101110 : OUT <= 2;  //224 / 110 = 2
    16'b11100000_01101111 : OUT <= 2;  //224 / 111 = 2
    16'b11100000_01110000 : OUT <= 2;  //224 / 112 = 2
    16'b11100000_01110001 : OUT <= 1;  //224 / 113 = 1
    16'b11100000_01110010 : OUT <= 1;  //224 / 114 = 1
    16'b11100000_01110011 : OUT <= 1;  //224 / 115 = 1
    16'b11100000_01110100 : OUT <= 1;  //224 / 116 = 1
    16'b11100000_01110101 : OUT <= 1;  //224 / 117 = 1
    16'b11100000_01110110 : OUT <= 1;  //224 / 118 = 1
    16'b11100000_01110111 : OUT <= 1;  //224 / 119 = 1
    16'b11100000_01111000 : OUT <= 1;  //224 / 120 = 1
    16'b11100000_01111001 : OUT <= 1;  //224 / 121 = 1
    16'b11100000_01111010 : OUT <= 1;  //224 / 122 = 1
    16'b11100000_01111011 : OUT <= 1;  //224 / 123 = 1
    16'b11100000_01111100 : OUT <= 1;  //224 / 124 = 1
    16'b11100000_01111101 : OUT <= 1;  //224 / 125 = 1
    16'b11100000_01111110 : OUT <= 1;  //224 / 126 = 1
    16'b11100000_01111111 : OUT <= 1;  //224 / 127 = 1
    16'b11100000_10000000 : OUT <= 1;  //224 / 128 = 1
    16'b11100000_10000001 : OUT <= 1;  //224 / 129 = 1
    16'b11100000_10000010 : OUT <= 1;  //224 / 130 = 1
    16'b11100000_10000011 : OUT <= 1;  //224 / 131 = 1
    16'b11100000_10000100 : OUT <= 1;  //224 / 132 = 1
    16'b11100000_10000101 : OUT <= 1;  //224 / 133 = 1
    16'b11100000_10000110 : OUT <= 1;  //224 / 134 = 1
    16'b11100000_10000111 : OUT <= 1;  //224 / 135 = 1
    16'b11100000_10001000 : OUT <= 1;  //224 / 136 = 1
    16'b11100000_10001001 : OUT <= 1;  //224 / 137 = 1
    16'b11100000_10001010 : OUT <= 1;  //224 / 138 = 1
    16'b11100000_10001011 : OUT <= 1;  //224 / 139 = 1
    16'b11100000_10001100 : OUT <= 1;  //224 / 140 = 1
    16'b11100000_10001101 : OUT <= 1;  //224 / 141 = 1
    16'b11100000_10001110 : OUT <= 1;  //224 / 142 = 1
    16'b11100000_10001111 : OUT <= 1;  //224 / 143 = 1
    16'b11100000_10010000 : OUT <= 1;  //224 / 144 = 1
    16'b11100000_10010001 : OUT <= 1;  //224 / 145 = 1
    16'b11100000_10010010 : OUT <= 1;  //224 / 146 = 1
    16'b11100000_10010011 : OUT <= 1;  //224 / 147 = 1
    16'b11100000_10010100 : OUT <= 1;  //224 / 148 = 1
    16'b11100000_10010101 : OUT <= 1;  //224 / 149 = 1
    16'b11100000_10010110 : OUT <= 1;  //224 / 150 = 1
    16'b11100000_10010111 : OUT <= 1;  //224 / 151 = 1
    16'b11100000_10011000 : OUT <= 1;  //224 / 152 = 1
    16'b11100000_10011001 : OUT <= 1;  //224 / 153 = 1
    16'b11100000_10011010 : OUT <= 1;  //224 / 154 = 1
    16'b11100000_10011011 : OUT <= 1;  //224 / 155 = 1
    16'b11100000_10011100 : OUT <= 1;  //224 / 156 = 1
    16'b11100000_10011101 : OUT <= 1;  //224 / 157 = 1
    16'b11100000_10011110 : OUT <= 1;  //224 / 158 = 1
    16'b11100000_10011111 : OUT <= 1;  //224 / 159 = 1
    16'b11100000_10100000 : OUT <= 1;  //224 / 160 = 1
    16'b11100000_10100001 : OUT <= 1;  //224 / 161 = 1
    16'b11100000_10100010 : OUT <= 1;  //224 / 162 = 1
    16'b11100000_10100011 : OUT <= 1;  //224 / 163 = 1
    16'b11100000_10100100 : OUT <= 1;  //224 / 164 = 1
    16'b11100000_10100101 : OUT <= 1;  //224 / 165 = 1
    16'b11100000_10100110 : OUT <= 1;  //224 / 166 = 1
    16'b11100000_10100111 : OUT <= 1;  //224 / 167 = 1
    16'b11100000_10101000 : OUT <= 1;  //224 / 168 = 1
    16'b11100000_10101001 : OUT <= 1;  //224 / 169 = 1
    16'b11100000_10101010 : OUT <= 1;  //224 / 170 = 1
    16'b11100000_10101011 : OUT <= 1;  //224 / 171 = 1
    16'b11100000_10101100 : OUT <= 1;  //224 / 172 = 1
    16'b11100000_10101101 : OUT <= 1;  //224 / 173 = 1
    16'b11100000_10101110 : OUT <= 1;  //224 / 174 = 1
    16'b11100000_10101111 : OUT <= 1;  //224 / 175 = 1
    16'b11100000_10110000 : OUT <= 1;  //224 / 176 = 1
    16'b11100000_10110001 : OUT <= 1;  //224 / 177 = 1
    16'b11100000_10110010 : OUT <= 1;  //224 / 178 = 1
    16'b11100000_10110011 : OUT <= 1;  //224 / 179 = 1
    16'b11100000_10110100 : OUT <= 1;  //224 / 180 = 1
    16'b11100000_10110101 : OUT <= 1;  //224 / 181 = 1
    16'b11100000_10110110 : OUT <= 1;  //224 / 182 = 1
    16'b11100000_10110111 : OUT <= 1;  //224 / 183 = 1
    16'b11100000_10111000 : OUT <= 1;  //224 / 184 = 1
    16'b11100000_10111001 : OUT <= 1;  //224 / 185 = 1
    16'b11100000_10111010 : OUT <= 1;  //224 / 186 = 1
    16'b11100000_10111011 : OUT <= 1;  //224 / 187 = 1
    16'b11100000_10111100 : OUT <= 1;  //224 / 188 = 1
    16'b11100000_10111101 : OUT <= 1;  //224 / 189 = 1
    16'b11100000_10111110 : OUT <= 1;  //224 / 190 = 1
    16'b11100000_10111111 : OUT <= 1;  //224 / 191 = 1
    16'b11100000_11000000 : OUT <= 1;  //224 / 192 = 1
    16'b11100000_11000001 : OUT <= 1;  //224 / 193 = 1
    16'b11100000_11000010 : OUT <= 1;  //224 / 194 = 1
    16'b11100000_11000011 : OUT <= 1;  //224 / 195 = 1
    16'b11100000_11000100 : OUT <= 1;  //224 / 196 = 1
    16'b11100000_11000101 : OUT <= 1;  //224 / 197 = 1
    16'b11100000_11000110 : OUT <= 1;  //224 / 198 = 1
    16'b11100000_11000111 : OUT <= 1;  //224 / 199 = 1
    16'b11100000_11001000 : OUT <= 1;  //224 / 200 = 1
    16'b11100000_11001001 : OUT <= 1;  //224 / 201 = 1
    16'b11100000_11001010 : OUT <= 1;  //224 / 202 = 1
    16'b11100000_11001011 : OUT <= 1;  //224 / 203 = 1
    16'b11100000_11001100 : OUT <= 1;  //224 / 204 = 1
    16'b11100000_11001101 : OUT <= 1;  //224 / 205 = 1
    16'b11100000_11001110 : OUT <= 1;  //224 / 206 = 1
    16'b11100000_11001111 : OUT <= 1;  //224 / 207 = 1
    16'b11100000_11010000 : OUT <= 1;  //224 / 208 = 1
    16'b11100000_11010001 : OUT <= 1;  //224 / 209 = 1
    16'b11100000_11010010 : OUT <= 1;  //224 / 210 = 1
    16'b11100000_11010011 : OUT <= 1;  //224 / 211 = 1
    16'b11100000_11010100 : OUT <= 1;  //224 / 212 = 1
    16'b11100000_11010101 : OUT <= 1;  //224 / 213 = 1
    16'b11100000_11010110 : OUT <= 1;  //224 / 214 = 1
    16'b11100000_11010111 : OUT <= 1;  //224 / 215 = 1
    16'b11100000_11011000 : OUT <= 1;  //224 / 216 = 1
    16'b11100000_11011001 : OUT <= 1;  //224 / 217 = 1
    16'b11100000_11011010 : OUT <= 1;  //224 / 218 = 1
    16'b11100000_11011011 : OUT <= 1;  //224 / 219 = 1
    16'b11100000_11011100 : OUT <= 1;  //224 / 220 = 1
    16'b11100000_11011101 : OUT <= 1;  //224 / 221 = 1
    16'b11100000_11011110 : OUT <= 1;  //224 / 222 = 1
    16'b11100000_11011111 : OUT <= 1;  //224 / 223 = 1
    16'b11100000_11100000 : OUT <= 1;  //224 / 224 = 1
    16'b11100000_11100001 : OUT <= 0;  //224 / 225 = 0
    16'b11100000_11100010 : OUT <= 0;  //224 / 226 = 0
    16'b11100000_11100011 : OUT <= 0;  //224 / 227 = 0
    16'b11100000_11100100 : OUT <= 0;  //224 / 228 = 0
    16'b11100000_11100101 : OUT <= 0;  //224 / 229 = 0
    16'b11100000_11100110 : OUT <= 0;  //224 / 230 = 0
    16'b11100000_11100111 : OUT <= 0;  //224 / 231 = 0
    16'b11100000_11101000 : OUT <= 0;  //224 / 232 = 0
    16'b11100000_11101001 : OUT <= 0;  //224 / 233 = 0
    16'b11100000_11101010 : OUT <= 0;  //224 / 234 = 0
    16'b11100000_11101011 : OUT <= 0;  //224 / 235 = 0
    16'b11100000_11101100 : OUT <= 0;  //224 / 236 = 0
    16'b11100000_11101101 : OUT <= 0;  //224 / 237 = 0
    16'b11100000_11101110 : OUT <= 0;  //224 / 238 = 0
    16'b11100000_11101111 : OUT <= 0;  //224 / 239 = 0
    16'b11100000_11110000 : OUT <= 0;  //224 / 240 = 0
    16'b11100000_11110001 : OUT <= 0;  //224 / 241 = 0
    16'b11100000_11110010 : OUT <= 0;  //224 / 242 = 0
    16'b11100000_11110011 : OUT <= 0;  //224 / 243 = 0
    16'b11100000_11110100 : OUT <= 0;  //224 / 244 = 0
    16'b11100000_11110101 : OUT <= 0;  //224 / 245 = 0
    16'b11100000_11110110 : OUT <= 0;  //224 / 246 = 0
    16'b11100000_11110111 : OUT <= 0;  //224 / 247 = 0
    16'b11100000_11111000 : OUT <= 0;  //224 / 248 = 0
    16'b11100000_11111001 : OUT <= 0;  //224 / 249 = 0
    16'b11100000_11111010 : OUT <= 0;  //224 / 250 = 0
    16'b11100000_11111011 : OUT <= 0;  //224 / 251 = 0
    16'b11100000_11111100 : OUT <= 0;  //224 / 252 = 0
    16'b11100000_11111101 : OUT <= 0;  //224 / 253 = 0
    16'b11100000_11111110 : OUT <= 0;  //224 / 254 = 0
    16'b11100000_11111111 : OUT <= 0;  //224 / 255 = 0
    16'b11100001_00000000 : OUT <= 0;  //225 / 0 = 0
    16'b11100001_00000001 : OUT <= 225;  //225 / 1 = 225
    16'b11100001_00000010 : OUT <= 112;  //225 / 2 = 112
    16'b11100001_00000011 : OUT <= 75;  //225 / 3 = 75
    16'b11100001_00000100 : OUT <= 56;  //225 / 4 = 56
    16'b11100001_00000101 : OUT <= 45;  //225 / 5 = 45
    16'b11100001_00000110 : OUT <= 37;  //225 / 6 = 37
    16'b11100001_00000111 : OUT <= 32;  //225 / 7 = 32
    16'b11100001_00001000 : OUT <= 28;  //225 / 8 = 28
    16'b11100001_00001001 : OUT <= 25;  //225 / 9 = 25
    16'b11100001_00001010 : OUT <= 22;  //225 / 10 = 22
    16'b11100001_00001011 : OUT <= 20;  //225 / 11 = 20
    16'b11100001_00001100 : OUT <= 18;  //225 / 12 = 18
    16'b11100001_00001101 : OUT <= 17;  //225 / 13 = 17
    16'b11100001_00001110 : OUT <= 16;  //225 / 14 = 16
    16'b11100001_00001111 : OUT <= 15;  //225 / 15 = 15
    16'b11100001_00010000 : OUT <= 14;  //225 / 16 = 14
    16'b11100001_00010001 : OUT <= 13;  //225 / 17 = 13
    16'b11100001_00010010 : OUT <= 12;  //225 / 18 = 12
    16'b11100001_00010011 : OUT <= 11;  //225 / 19 = 11
    16'b11100001_00010100 : OUT <= 11;  //225 / 20 = 11
    16'b11100001_00010101 : OUT <= 10;  //225 / 21 = 10
    16'b11100001_00010110 : OUT <= 10;  //225 / 22 = 10
    16'b11100001_00010111 : OUT <= 9;  //225 / 23 = 9
    16'b11100001_00011000 : OUT <= 9;  //225 / 24 = 9
    16'b11100001_00011001 : OUT <= 9;  //225 / 25 = 9
    16'b11100001_00011010 : OUT <= 8;  //225 / 26 = 8
    16'b11100001_00011011 : OUT <= 8;  //225 / 27 = 8
    16'b11100001_00011100 : OUT <= 8;  //225 / 28 = 8
    16'b11100001_00011101 : OUT <= 7;  //225 / 29 = 7
    16'b11100001_00011110 : OUT <= 7;  //225 / 30 = 7
    16'b11100001_00011111 : OUT <= 7;  //225 / 31 = 7
    16'b11100001_00100000 : OUT <= 7;  //225 / 32 = 7
    16'b11100001_00100001 : OUT <= 6;  //225 / 33 = 6
    16'b11100001_00100010 : OUT <= 6;  //225 / 34 = 6
    16'b11100001_00100011 : OUT <= 6;  //225 / 35 = 6
    16'b11100001_00100100 : OUT <= 6;  //225 / 36 = 6
    16'b11100001_00100101 : OUT <= 6;  //225 / 37 = 6
    16'b11100001_00100110 : OUT <= 5;  //225 / 38 = 5
    16'b11100001_00100111 : OUT <= 5;  //225 / 39 = 5
    16'b11100001_00101000 : OUT <= 5;  //225 / 40 = 5
    16'b11100001_00101001 : OUT <= 5;  //225 / 41 = 5
    16'b11100001_00101010 : OUT <= 5;  //225 / 42 = 5
    16'b11100001_00101011 : OUT <= 5;  //225 / 43 = 5
    16'b11100001_00101100 : OUT <= 5;  //225 / 44 = 5
    16'b11100001_00101101 : OUT <= 5;  //225 / 45 = 5
    16'b11100001_00101110 : OUT <= 4;  //225 / 46 = 4
    16'b11100001_00101111 : OUT <= 4;  //225 / 47 = 4
    16'b11100001_00110000 : OUT <= 4;  //225 / 48 = 4
    16'b11100001_00110001 : OUT <= 4;  //225 / 49 = 4
    16'b11100001_00110010 : OUT <= 4;  //225 / 50 = 4
    16'b11100001_00110011 : OUT <= 4;  //225 / 51 = 4
    16'b11100001_00110100 : OUT <= 4;  //225 / 52 = 4
    16'b11100001_00110101 : OUT <= 4;  //225 / 53 = 4
    16'b11100001_00110110 : OUT <= 4;  //225 / 54 = 4
    16'b11100001_00110111 : OUT <= 4;  //225 / 55 = 4
    16'b11100001_00111000 : OUT <= 4;  //225 / 56 = 4
    16'b11100001_00111001 : OUT <= 3;  //225 / 57 = 3
    16'b11100001_00111010 : OUT <= 3;  //225 / 58 = 3
    16'b11100001_00111011 : OUT <= 3;  //225 / 59 = 3
    16'b11100001_00111100 : OUT <= 3;  //225 / 60 = 3
    16'b11100001_00111101 : OUT <= 3;  //225 / 61 = 3
    16'b11100001_00111110 : OUT <= 3;  //225 / 62 = 3
    16'b11100001_00111111 : OUT <= 3;  //225 / 63 = 3
    16'b11100001_01000000 : OUT <= 3;  //225 / 64 = 3
    16'b11100001_01000001 : OUT <= 3;  //225 / 65 = 3
    16'b11100001_01000010 : OUT <= 3;  //225 / 66 = 3
    16'b11100001_01000011 : OUT <= 3;  //225 / 67 = 3
    16'b11100001_01000100 : OUT <= 3;  //225 / 68 = 3
    16'b11100001_01000101 : OUT <= 3;  //225 / 69 = 3
    16'b11100001_01000110 : OUT <= 3;  //225 / 70 = 3
    16'b11100001_01000111 : OUT <= 3;  //225 / 71 = 3
    16'b11100001_01001000 : OUT <= 3;  //225 / 72 = 3
    16'b11100001_01001001 : OUT <= 3;  //225 / 73 = 3
    16'b11100001_01001010 : OUT <= 3;  //225 / 74 = 3
    16'b11100001_01001011 : OUT <= 3;  //225 / 75 = 3
    16'b11100001_01001100 : OUT <= 2;  //225 / 76 = 2
    16'b11100001_01001101 : OUT <= 2;  //225 / 77 = 2
    16'b11100001_01001110 : OUT <= 2;  //225 / 78 = 2
    16'b11100001_01001111 : OUT <= 2;  //225 / 79 = 2
    16'b11100001_01010000 : OUT <= 2;  //225 / 80 = 2
    16'b11100001_01010001 : OUT <= 2;  //225 / 81 = 2
    16'b11100001_01010010 : OUT <= 2;  //225 / 82 = 2
    16'b11100001_01010011 : OUT <= 2;  //225 / 83 = 2
    16'b11100001_01010100 : OUT <= 2;  //225 / 84 = 2
    16'b11100001_01010101 : OUT <= 2;  //225 / 85 = 2
    16'b11100001_01010110 : OUT <= 2;  //225 / 86 = 2
    16'b11100001_01010111 : OUT <= 2;  //225 / 87 = 2
    16'b11100001_01011000 : OUT <= 2;  //225 / 88 = 2
    16'b11100001_01011001 : OUT <= 2;  //225 / 89 = 2
    16'b11100001_01011010 : OUT <= 2;  //225 / 90 = 2
    16'b11100001_01011011 : OUT <= 2;  //225 / 91 = 2
    16'b11100001_01011100 : OUT <= 2;  //225 / 92 = 2
    16'b11100001_01011101 : OUT <= 2;  //225 / 93 = 2
    16'b11100001_01011110 : OUT <= 2;  //225 / 94 = 2
    16'b11100001_01011111 : OUT <= 2;  //225 / 95 = 2
    16'b11100001_01100000 : OUT <= 2;  //225 / 96 = 2
    16'b11100001_01100001 : OUT <= 2;  //225 / 97 = 2
    16'b11100001_01100010 : OUT <= 2;  //225 / 98 = 2
    16'b11100001_01100011 : OUT <= 2;  //225 / 99 = 2
    16'b11100001_01100100 : OUT <= 2;  //225 / 100 = 2
    16'b11100001_01100101 : OUT <= 2;  //225 / 101 = 2
    16'b11100001_01100110 : OUT <= 2;  //225 / 102 = 2
    16'b11100001_01100111 : OUT <= 2;  //225 / 103 = 2
    16'b11100001_01101000 : OUT <= 2;  //225 / 104 = 2
    16'b11100001_01101001 : OUT <= 2;  //225 / 105 = 2
    16'b11100001_01101010 : OUT <= 2;  //225 / 106 = 2
    16'b11100001_01101011 : OUT <= 2;  //225 / 107 = 2
    16'b11100001_01101100 : OUT <= 2;  //225 / 108 = 2
    16'b11100001_01101101 : OUT <= 2;  //225 / 109 = 2
    16'b11100001_01101110 : OUT <= 2;  //225 / 110 = 2
    16'b11100001_01101111 : OUT <= 2;  //225 / 111 = 2
    16'b11100001_01110000 : OUT <= 2;  //225 / 112 = 2
    16'b11100001_01110001 : OUT <= 1;  //225 / 113 = 1
    16'b11100001_01110010 : OUT <= 1;  //225 / 114 = 1
    16'b11100001_01110011 : OUT <= 1;  //225 / 115 = 1
    16'b11100001_01110100 : OUT <= 1;  //225 / 116 = 1
    16'b11100001_01110101 : OUT <= 1;  //225 / 117 = 1
    16'b11100001_01110110 : OUT <= 1;  //225 / 118 = 1
    16'b11100001_01110111 : OUT <= 1;  //225 / 119 = 1
    16'b11100001_01111000 : OUT <= 1;  //225 / 120 = 1
    16'b11100001_01111001 : OUT <= 1;  //225 / 121 = 1
    16'b11100001_01111010 : OUT <= 1;  //225 / 122 = 1
    16'b11100001_01111011 : OUT <= 1;  //225 / 123 = 1
    16'b11100001_01111100 : OUT <= 1;  //225 / 124 = 1
    16'b11100001_01111101 : OUT <= 1;  //225 / 125 = 1
    16'b11100001_01111110 : OUT <= 1;  //225 / 126 = 1
    16'b11100001_01111111 : OUT <= 1;  //225 / 127 = 1
    16'b11100001_10000000 : OUT <= 1;  //225 / 128 = 1
    16'b11100001_10000001 : OUT <= 1;  //225 / 129 = 1
    16'b11100001_10000010 : OUT <= 1;  //225 / 130 = 1
    16'b11100001_10000011 : OUT <= 1;  //225 / 131 = 1
    16'b11100001_10000100 : OUT <= 1;  //225 / 132 = 1
    16'b11100001_10000101 : OUT <= 1;  //225 / 133 = 1
    16'b11100001_10000110 : OUT <= 1;  //225 / 134 = 1
    16'b11100001_10000111 : OUT <= 1;  //225 / 135 = 1
    16'b11100001_10001000 : OUT <= 1;  //225 / 136 = 1
    16'b11100001_10001001 : OUT <= 1;  //225 / 137 = 1
    16'b11100001_10001010 : OUT <= 1;  //225 / 138 = 1
    16'b11100001_10001011 : OUT <= 1;  //225 / 139 = 1
    16'b11100001_10001100 : OUT <= 1;  //225 / 140 = 1
    16'b11100001_10001101 : OUT <= 1;  //225 / 141 = 1
    16'b11100001_10001110 : OUT <= 1;  //225 / 142 = 1
    16'b11100001_10001111 : OUT <= 1;  //225 / 143 = 1
    16'b11100001_10010000 : OUT <= 1;  //225 / 144 = 1
    16'b11100001_10010001 : OUT <= 1;  //225 / 145 = 1
    16'b11100001_10010010 : OUT <= 1;  //225 / 146 = 1
    16'b11100001_10010011 : OUT <= 1;  //225 / 147 = 1
    16'b11100001_10010100 : OUT <= 1;  //225 / 148 = 1
    16'b11100001_10010101 : OUT <= 1;  //225 / 149 = 1
    16'b11100001_10010110 : OUT <= 1;  //225 / 150 = 1
    16'b11100001_10010111 : OUT <= 1;  //225 / 151 = 1
    16'b11100001_10011000 : OUT <= 1;  //225 / 152 = 1
    16'b11100001_10011001 : OUT <= 1;  //225 / 153 = 1
    16'b11100001_10011010 : OUT <= 1;  //225 / 154 = 1
    16'b11100001_10011011 : OUT <= 1;  //225 / 155 = 1
    16'b11100001_10011100 : OUT <= 1;  //225 / 156 = 1
    16'b11100001_10011101 : OUT <= 1;  //225 / 157 = 1
    16'b11100001_10011110 : OUT <= 1;  //225 / 158 = 1
    16'b11100001_10011111 : OUT <= 1;  //225 / 159 = 1
    16'b11100001_10100000 : OUT <= 1;  //225 / 160 = 1
    16'b11100001_10100001 : OUT <= 1;  //225 / 161 = 1
    16'b11100001_10100010 : OUT <= 1;  //225 / 162 = 1
    16'b11100001_10100011 : OUT <= 1;  //225 / 163 = 1
    16'b11100001_10100100 : OUT <= 1;  //225 / 164 = 1
    16'b11100001_10100101 : OUT <= 1;  //225 / 165 = 1
    16'b11100001_10100110 : OUT <= 1;  //225 / 166 = 1
    16'b11100001_10100111 : OUT <= 1;  //225 / 167 = 1
    16'b11100001_10101000 : OUT <= 1;  //225 / 168 = 1
    16'b11100001_10101001 : OUT <= 1;  //225 / 169 = 1
    16'b11100001_10101010 : OUT <= 1;  //225 / 170 = 1
    16'b11100001_10101011 : OUT <= 1;  //225 / 171 = 1
    16'b11100001_10101100 : OUT <= 1;  //225 / 172 = 1
    16'b11100001_10101101 : OUT <= 1;  //225 / 173 = 1
    16'b11100001_10101110 : OUT <= 1;  //225 / 174 = 1
    16'b11100001_10101111 : OUT <= 1;  //225 / 175 = 1
    16'b11100001_10110000 : OUT <= 1;  //225 / 176 = 1
    16'b11100001_10110001 : OUT <= 1;  //225 / 177 = 1
    16'b11100001_10110010 : OUT <= 1;  //225 / 178 = 1
    16'b11100001_10110011 : OUT <= 1;  //225 / 179 = 1
    16'b11100001_10110100 : OUT <= 1;  //225 / 180 = 1
    16'b11100001_10110101 : OUT <= 1;  //225 / 181 = 1
    16'b11100001_10110110 : OUT <= 1;  //225 / 182 = 1
    16'b11100001_10110111 : OUT <= 1;  //225 / 183 = 1
    16'b11100001_10111000 : OUT <= 1;  //225 / 184 = 1
    16'b11100001_10111001 : OUT <= 1;  //225 / 185 = 1
    16'b11100001_10111010 : OUT <= 1;  //225 / 186 = 1
    16'b11100001_10111011 : OUT <= 1;  //225 / 187 = 1
    16'b11100001_10111100 : OUT <= 1;  //225 / 188 = 1
    16'b11100001_10111101 : OUT <= 1;  //225 / 189 = 1
    16'b11100001_10111110 : OUT <= 1;  //225 / 190 = 1
    16'b11100001_10111111 : OUT <= 1;  //225 / 191 = 1
    16'b11100001_11000000 : OUT <= 1;  //225 / 192 = 1
    16'b11100001_11000001 : OUT <= 1;  //225 / 193 = 1
    16'b11100001_11000010 : OUT <= 1;  //225 / 194 = 1
    16'b11100001_11000011 : OUT <= 1;  //225 / 195 = 1
    16'b11100001_11000100 : OUT <= 1;  //225 / 196 = 1
    16'b11100001_11000101 : OUT <= 1;  //225 / 197 = 1
    16'b11100001_11000110 : OUT <= 1;  //225 / 198 = 1
    16'b11100001_11000111 : OUT <= 1;  //225 / 199 = 1
    16'b11100001_11001000 : OUT <= 1;  //225 / 200 = 1
    16'b11100001_11001001 : OUT <= 1;  //225 / 201 = 1
    16'b11100001_11001010 : OUT <= 1;  //225 / 202 = 1
    16'b11100001_11001011 : OUT <= 1;  //225 / 203 = 1
    16'b11100001_11001100 : OUT <= 1;  //225 / 204 = 1
    16'b11100001_11001101 : OUT <= 1;  //225 / 205 = 1
    16'b11100001_11001110 : OUT <= 1;  //225 / 206 = 1
    16'b11100001_11001111 : OUT <= 1;  //225 / 207 = 1
    16'b11100001_11010000 : OUT <= 1;  //225 / 208 = 1
    16'b11100001_11010001 : OUT <= 1;  //225 / 209 = 1
    16'b11100001_11010010 : OUT <= 1;  //225 / 210 = 1
    16'b11100001_11010011 : OUT <= 1;  //225 / 211 = 1
    16'b11100001_11010100 : OUT <= 1;  //225 / 212 = 1
    16'b11100001_11010101 : OUT <= 1;  //225 / 213 = 1
    16'b11100001_11010110 : OUT <= 1;  //225 / 214 = 1
    16'b11100001_11010111 : OUT <= 1;  //225 / 215 = 1
    16'b11100001_11011000 : OUT <= 1;  //225 / 216 = 1
    16'b11100001_11011001 : OUT <= 1;  //225 / 217 = 1
    16'b11100001_11011010 : OUT <= 1;  //225 / 218 = 1
    16'b11100001_11011011 : OUT <= 1;  //225 / 219 = 1
    16'b11100001_11011100 : OUT <= 1;  //225 / 220 = 1
    16'b11100001_11011101 : OUT <= 1;  //225 / 221 = 1
    16'b11100001_11011110 : OUT <= 1;  //225 / 222 = 1
    16'b11100001_11011111 : OUT <= 1;  //225 / 223 = 1
    16'b11100001_11100000 : OUT <= 1;  //225 / 224 = 1
    16'b11100001_11100001 : OUT <= 1;  //225 / 225 = 1
    16'b11100001_11100010 : OUT <= 0;  //225 / 226 = 0
    16'b11100001_11100011 : OUT <= 0;  //225 / 227 = 0
    16'b11100001_11100100 : OUT <= 0;  //225 / 228 = 0
    16'b11100001_11100101 : OUT <= 0;  //225 / 229 = 0
    16'b11100001_11100110 : OUT <= 0;  //225 / 230 = 0
    16'b11100001_11100111 : OUT <= 0;  //225 / 231 = 0
    16'b11100001_11101000 : OUT <= 0;  //225 / 232 = 0
    16'b11100001_11101001 : OUT <= 0;  //225 / 233 = 0
    16'b11100001_11101010 : OUT <= 0;  //225 / 234 = 0
    16'b11100001_11101011 : OUT <= 0;  //225 / 235 = 0
    16'b11100001_11101100 : OUT <= 0;  //225 / 236 = 0
    16'b11100001_11101101 : OUT <= 0;  //225 / 237 = 0
    16'b11100001_11101110 : OUT <= 0;  //225 / 238 = 0
    16'b11100001_11101111 : OUT <= 0;  //225 / 239 = 0
    16'b11100001_11110000 : OUT <= 0;  //225 / 240 = 0
    16'b11100001_11110001 : OUT <= 0;  //225 / 241 = 0
    16'b11100001_11110010 : OUT <= 0;  //225 / 242 = 0
    16'b11100001_11110011 : OUT <= 0;  //225 / 243 = 0
    16'b11100001_11110100 : OUT <= 0;  //225 / 244 = 0
    16'b11100001_11110101 : OUT <= 0;  //225 / 245 = 0
    16'b11100001_11110110 : OUT <= 0;  //225 / 246 = 0
    16'b11100001_11110111 : OUT <= 0;  //225 / 247 = 0
    16'b11100001_11111000 : OUT <= 0;  //225 / 248 = 0
    16'b11100001_11111001 : OUT <= 0;  //225 / 249 = 0
    16'b11100001_11111010 : OUT <= 0;  //225 / 250 = 0
    16'b11100001_11111011 : OUT <= 0;  //225 / 251 = 0
    16'b11100001_11111100 : OUT <= 0;  //225 / 252 = 0
    16'b11100001_11111101 : OUT <= 0;  //225 / 253 = 0
    16'b11100001_11111110 : OUT <= 0;  //225 / 254 = 0
    16'b11100001_11111111 : OUT <= 0;  //225 / 255 = 0
    16'b11100010_00000000 : OUT <= 0;  //226 / 0 = 0
    16'b11100010_00000001 : OUT <= 226;  //226 / 1 = 226
    16'b11100010_00000010 : OUT <= 113;  //226 / 2 = 113
    16'b11100010_00000011 : OUT <= 75;  //226 / 3 = 75
    16'b11100010_00000100 : OUT <= 56;  //226 / 4 = 56
    16'b11100010_00000101 : OUT <= 45;  //226 / 5 = 45
    16'b11100010_00000110 : OUT <= 37;  //226 / 6 = 37
    16'b11100010_00000111 : OUT <= 32;  //226 / 7 = 32
    16'b11100010_00001000 : OUT <= 28;  //226 / 8 = 28
    16'b11100010_00001001 : OUT <= 25;  //226 / 9 = 25
    16'b11100010_00001010 : OUT <= 22;  //226 / 10 = 22
    16'b11100010_00001011 : OUT <= 20;  //226 / 11 = 20
    16'b11100010_00001100 : OUT <= 18;  //226 / 12 = 18
    16'b11100010_00001101 : OUT <= 17;  //226 / 13 = 17
    16'b11100010_00001110 : OUT <= 16;  //226 / 14 = 16
    16'b11100010_00001111 : OUT <= 15;  //226 / 15 = 15
    16'b11100010_00010000 : OUT <= 14;  //226 / 16 = 14
    16'b11100010_00010001 : OUT <= 13;  //226 / 17 = 13
    16'b11100010_00010010 : OUT <= 12;  //226 / 18 = 12
    16'b11100010_00010011 : OUT <= 11;  //226 / 19 = 11
    16'b11100010_00010100 : OUT <= 11;  //226 / 20 = 11
    16'b11100010_00010101 : OUT <= 10;  //226 / 21 = 10
    16'b11100010_00010110 : OUT <= 10;  //226 / 22 = 10
    16'b11100010_00010111 : OUT <= 9;  //226 / 23 = 9
    16'b11100010_00011000 : OUT <= 9;  //226 / 24 = 9
    16'b11100010_00011001 : OUT <= 9;  //226 / 25 = 9
    16'b11100010_00011010 : OUT <= 8;  //226 / 26 = 8
    16'b11100010_00011011 : OUT <= 8;  //226 / 27 = 8
    16'b11100010_00011100 : OUT <= 8;  //226 / 28 = 8
    16'b11100010_00011101 : OUT <= 7;  //226 / 29 = 7
    16'b11100010_00011110 : OUT <= 7;  //226 / 30 = 7
    16'b11100010_00011111 : OUT <= 7;  //226 / 31 = 7
    16'b11100010_00100000 : OUT <= 7;  //226 / 32 = 7
    16'b11100010_00100001 : OUT <= 6;  //226 / 33 = 6
    16'b11100010_00100010 : OUT <= 6;  //226 / 34 = 6
    16'b11100010_00100011 : OUT <= 6;  //226 / 35 = 6
    16'b11100010_00100100 : OUT <= 6;  //226 / 36 = 6
    16'b11100010_00100101 : OUT <= 6;  //226 / 37 = 6
    16'b11100010_00100110 : OUT <= 5;  //226 / 38 = 5
    16'b11100010_00100111 : OUT <= 5;  //226 / 39 = 5
    16'b11100010_00101000 : OUT <= 5;  //226 / 40 = 5
    16'b11100010_00101001 : OUT <= 5;  //226 / 41 = 5
    16'b11100010_00101010 : OUT <= 5;  //226 / 42 = 5
    16'b11100010_00101011 : OUT <= 5;  //226 / 43 = 5
    16'b11100010_00101100 : OUT <= 5;  //226 / 44 = 5
    16'b11100010_00101101 : OUT <= 5;  //226 / 45 = 5
    16'b11100010_00101110 : OUT <= 4;  //226 / 46 = 4
    16'b11100010_00101111 : OUT <= 4;  //226 / 47 = 4
    16'b11100010_00110000 : OUT <= 4;  //226 / 48 = 4
    16'b11100010_00110001 : OUT <= 4;  //226 / 49 = 4
    16'b11100010_00110010 : OUT <= 4;  //226 / 50 = 4
    16'b11100010_00110011 : OUT <= 4;  //226 / 51 = 4
    16'b11100010_00110100 : OUT <= 4;  //226 / 52 = 4
    16'b11100010_00110101 : OUT <= 4;  //226 / 53 = 4
    16'b11100010_00110110 : OUT <= 4;  //226 / 54 = 4
    16'b11100010_00110111 : OUT <= 4;  //226 / 55 = 4
    16'b11100010_00111000 : OUT <= 4;  //226 / 56 = 4
    16'b11100010_00111001 : OUT <= 3;  //226 / 57 = 3
    16'b11100010_00111010 : OUT <= 3;  //226 / 58 = 3
    16'b11100010_00111011 : OUT <= 3;  //226 / 59 = 3
    16'b11100010_00111100 : OUT <= 3;  //226 / 60 = 3
    16'b11100010_00111101 : OUT <= 3;  //226 / 61 = 3
    16'b11100010_00111110 : OUT <= 3;  //226 / 62 = 3
    16'b11100010_00111111 : OUT <= 3;  //226 / 63 = 3
    16'b11100010_01000000 : OUT <= 3;  //226 / 64 = 3
    16'b11100010_01000001 : OUT <= 3;  //226 / 65 = 3
    16'b11100010_01000010 : OUT <= 3;  //226 / 66 = 3
    16'b11100010_01000011 : OUT <= 3;  //226 / 67 = 3
    16'b11100010_01000100 : OUT <= 3;  //226 / 68 = 3
    16'b11100010_01000101 : OUT <= 3;  //226 / 69 = 3
    16'b11100010_01000110 : OUT <= 3;  //226 / 70 = 3
    16'b11100010_01000111 : OUT <= 3;  //226 / 71 = 3
    16'b11100010_01001000 : OUT <= 3;  //226 / 72 = 3
    16'b11100010_01001001 : OUT <= 3;  //226 / 73 = 3
    16'b11100010_01001010 : OUT <= 3;  //226 / 74 = 3
    16'b11100010_01001011 : OUT <= 3;  //226 / 75 = 3
    16'b11100010_01001100 : OUT <= 2;  //226 / 76 = 2
    16'b11100010_01001101 : OUT <= 2;  //226 / 77 = 2
    16'b11100010_01001110 : OUT <= 2;  //226 / 78 = 2
    16'b11100010_01001111 : OUT <= 2;  //226 / 79 = 2
    16'b11100010_01010000 : OUT <= 2;  //226 / 80 = 2
    16'b11100010_01010001 : OUT <= 2;  //226 / 81 = 2
    16'b11100010_01010010 : OUT <= 2;  //226 / 82 = 2
    16'b11100010_01010011 : OUT <= 2;  //226 / 83 = 2
    16'b11100010_01010100 : OUT <= 2;  //226 / 84 = 2
    16'b11100010_01010101 : OUT <= 2;  //226 / 85 = 2
    16'b11100010_01010110 : OUT <= 2;  //226 / 86 = 2
    16'b11100010_01010111 : OUT <= 2;  //226 / 87 = 2
    16'b11100010_01011000 : OUT <= 2;  //226 / 88 = 2
    16'b11100010_01011001 : OUT <= 2;  //226 / 89 = 2
    16'b11100010_01011010 : OUT <= 2;  //226 / 90 = 2
    16'b11100010_01011011 : OUT <= 2;  //226 / 91 = 2
    16'b11100010_01011100 : OUT <= 2;  //226 / 92 = 2
    16'b11100010_01011101 : OUT <= 2;  //226 / 93 = 2
    16'b11100010_01011110 : OUT <= 2;  //226 / 94 = 2
    16'b11100010_01011111 : OUT <= 2;  //226 / 95 = 2
    16'b11100010_01100000 : OUT <= 2;  //226 / 96 = 2
    16'b11100010_01100001 : OUT <= 2;  //226 / 97 = 2
    16'b11100010_01100010 : OUT <= 2;  //226 / 98 = 2
    16'b11100010_01100011 : OUT <= 2;  //226 / 99 = 2
    16'b11100010_01100100 : OUT <= 2;  //226 / 100 = 2
    16'b11100010_01100101 : OUT <= 2;  //226 / 101 = 2
    16'b11100010_01100110 : OUT <= 2;  //226 / 102 = 2
    16'b11100010_01100111 : OUT <= 2;  //226 / 103 = 2
    16'b11100010_01101000 : OUT <= 2;  //226 / 104 = 2
    16'b11100010_01101001 : OUT <= 2;  //226 / 105 = 2
    16'b11100010_01101010 : OUT <= 2;  //226 / 106 = 2
    16'b11100010_01101011 : OUT <= 2;  //226 / 107 = 2
    16'b11100010_01101100 : OUT <= 2;  //226 / 108 = 2
    16'b11100010_01101101 : OUT <= 2;  //226 / 109 = 2
    16'b11100010_01101110 : OUT <= 2;  //226 / 110 = 2
    16'b11100010_01101111 : OUT <= 2;  //226 / 111 = 2
    16'b11100010_01110000 : OUT <= 2;  //226 / 112 = 2
    16'b11100010_01110001 : OUT <= 2;  //226 / 113 = 2
    16'b11100010_01110010 : OUT <= 1;  //226 / 114 = 1
    16'b11100010_01110011 : OUT <= 1;  //226 / 115 = 1
    16'b11100010_01110100 : OUT <= 1;  //226 / 116 = 1
    16'b11100010_01110101 : OUT <= 1;  //226 / 117 = 1
    16'b11100010_01110110 : OUT <= 1;  //226 / 118 = 1
    16'b11100010_01110111 : OUT <= 1;  //226 / 119 = 1
    16'b11100010_01111000 : OUT <= 1;  //226 / 120 = 1
    16'b11100010_01111001 : OUT <= 1;  //226 / 121 = 1
    16'b11100010_01111010 : OUT <= 1;  //226 / 122 = 1
    16'b11100010_01111011 : OUT <= 1;  //226 / 123 = 1
    16'b11100010_01111100 : OUT <= 1;  //226 / 124 = 1
    16'b11100010_01111101 : OUT <= 1;  //226 / 125 = 1
    16'b11100010_01111110 : OUT <= 1;  //226 / 126 = 1
    16'b11100010_01111111 : OUT <= 1;  //226 / 127 = 1
    16'b11100010_10000000 : OUT <= 1;  //226 / 128 = 1
    16'b11100010_10000001 : OUT <= 1;  //226 / 129 = 1
    16'b11100010_10000010 : OUT <= 1;  //226 / 130 = 1
    16'b11100010_10000011 : OUT <= 1;  //226 / 131 = 1
    16'b11100010_10000100 : OUT <= 1;  //226 / 132 = 1
    16'b11100010_10000101 : OUT <= 1;  //226 / 133 = 1
    16'b11100010_10000110 : OUT <= 1;  //226 / 134 = 1
    16'b11100010_10000111 : OUT <= 1;  //226 / 135 = 1
    16'b11100010_10001000 : OUT <= 1;  //226 / 136 = 1
    16'b11100010_10001001 : OUT <= 1;  //226 / 137 = 1
    16'b11100010_10001010 : OUT <= 1;  //226 / 138 = 1
    16'b11100010_10001011 : OUT <= 1;  //226 / 139 = 1
    16'b11100010_10001100 : OUT <= 1;  //226 / 140 = 1
    16'b11100010_10001101 : OUT <= 1;  //226 / 141 = 1
    16'b11100010_10001110 : OUT <= 1;  //226 / 142 = 1
    16'b11100010_10001111 : OUT <= 1;  //226 / 143 = 1
    16'b11100010_10010000 : OUT <= 1;  //226 / 144 = 1
    16'b11100010_10010001 : OUT <= 1;  //226 / 145 = 1
    16'b11100010_10010010 : OUT <= 1;  //226 / 146 = 1
    16'b11100010_10010011 : OUT <= 1;  //226 / 147 = 1
    16'b11100010_10010100 : OUT <= 1;  //226 / 148 = 1
    16'b11100010_10010101 : OUT <= 1;  //226 / 149 = 1
    16'b11100010_10010110 : OUT <= 1;  //226 / 150 = 1
    16'b11100010_10010111 : OUT <= 1;  //226 / 151 = 1
    16'b11100010_10011000 : OUT <= 1;  //226 / 152 = 1
    16'b11100010_10011001 : OUT <= 1;  //226 / 153 = 1
    16'b11100010_10011010 : OUT <= 1;  //226 / 154 = 1
    16'b11100010_10011011 : OUT <= 1;  //226 / 155 = 1
    16'b11100010_10011100 : OUT <= 1;  //226 / 156 = 1
    16'b11100010_10011101 : OUT <= 1;  //226 / 157 = 1
    16'b11100010_10011110 : OUT <= 1;  //226 / 158 = 1
    16'b11100010_10011111 : OUT <= 1;  //226 / 159 = 1
    16'b11100010_10100000 : OUT <= 1;  //226 / 160 = 1
    16'b11100010_10100001 : OUT <= 1;  //226 / 161 = 1
    16'b11100010_10100010 : OUT <= 1;  //226 / 162 = 1
    16'b11100010_10100011 : OUT <= 1;  //226 / 163 = 1
    16'b11100010_10100100 : OUT <= 1;  //226 / 164 = 1
    16'b11100010_10100101 : OUT <= 1;  //226 / 165 = 1
    16'b11100010_10100110 : OUT <= 1;  //226 / 166 = 1
    16'b11100010_10100111 : OUT <= 1;  //226 / 167 = 1
    16'b11100010_10101000 : OUT <= 1;  //226 / 168 = 1
    16'b11100010_10101001 : OUT <= 1;  //226 / 169 = 1
    16'b11100010_10101010 : OUT <= 1;  //226 / 170 = 1
    16'b11100010_10101011 : OUT <= 1;  //226 / 171 = 1
    16'b11100010_10101100 : OUT <= 1;  //226 / 172 = 1
    16'b11100010_10101101 : OUT <= 1;  //226 / 173 = 1
    16'b11100010_10101110 : OUT <= 1;  //226 / 174 = 1
    16'b11100010_10101111 : OUT <= 1;  //226 / 175 = 1
    16'b11100010_10110000 : OUT <= 1;  //226 / 176 = 1
    16'b11100010_10110001 : OUT <= 1;  //226 / 177 = 1
    16'b11100010_10110010 : OUT <= 1;  //226 / 178 = 1
    16'b11100010_10110011 : OUT <= 1;  //226 / 179 = 1
    16'b11100010_10110100 : OUT <= 1;  //226 / 180 = 1
    16'b11100010_10110101 : OUT <= 1;  //226 / 181 = 1
    16'b11100010_10110110 : OUT <= 1;  //226 / 182 = 1
    16'b11100010_10110111 : OUT <= 1;  //226 / 183 = 1
    16'b11100010_10111000 : OUT <= 1;  //226 / 184 = 1
    16'b11100010_10111001 : OUT <= 1;  //226 / 185 = 1
    16'b11100010_10111010 : OUT <= 1;  //226 / 186 = 1
    16'b11100010_10111011 : OUT <= 1;  //226 / 187 = 1
    16'b11100010_10111100 : OUT <= 1;  //226 / 188 = 1
    16'b11100010_10111101 : OUT <= 1;  //226 / 189 = 1
    16'b11100010_10111110 : OUT <= 1;  //226 / 190 = 1
    16'b11100010_10111111 : OUT <= 1;  //226 / 191 = 1
    16'b11100010_11000000 : OUT <= 1;  //226 / 192 = 1
    16'b11100010_11000001 : OUT <= 1;  //226 / 193 = 1
    16'b11100010_11000010 : OUT <= 1;  //226 / 194 = 1
    16'b11100010_11000011 : OUT <= 1;  //226 / 195 = 1
    16'b11100010_11000100 : OUT <= 1;  //226 / 196 = 1
    16'b11100010_11000101 : OUT <= 1;  //226 / 197 = 1
    16'b11100010_11000110 : OUT <= 1;  //226 / 198 = 1
    16'b11100010_11000111 : OUT <= 1;  //226 / 199 = 1
    16'b11100010_11001000 : OUT <= 1;  //226 / 200 = 1
    16'b11100010_11001001 : OUT <= 1;  //226 / 201 = 1
    16'b11100010_11001010 : OUT <= 1;  //226 / 202 = 1
    16'b11100010_11001011 : OUT <= 1;  //226 / 203 = 1
    16'b11100010_11001100 : OUT <= 1;  //226 / 204 = 1
    16'b11100010_11001101 : OUT <= 1;  //226 / 205 = 1
    16'b11100010_11001110 : OUT <= 1;  //226 / 206 = 1
    16'b11100010_11001111 : OUT <= 1;  //226 / 207 = 1
    16'b11100010_11010000 : OUT <= 1;  //226 / 208 = 1
    16'b11100010_11010001 : OUT <= 1;  //226 / 209 = 1
    16'b11100010_11010010 : OUT <= 1;  //226 / 210 = 1
    16'b11100010_11010011 : OUT <= 1;  //226 / 211 = 1
    16'b11100010_11010100 : OUT <= 1;  //226 / 212 = 1
    16'b11100010_11010101 : OUT <= 1;  //226 / 213 = 1
    16'b11100010_11010110 : OUT <= 1;  //226 / 214 = 1
    16'b11100010_11010111 : OUT <= 1;  //226 / 215 = 1
    16'b11100010_11011000 : OUT <= 1;  //226 / 216 = 1
    16'b11100010_11011001 : OUT <= 1;  //226 / 217 = 1
    16'b11100010_11011010 : OUT <= 1;  //226 / 218 = 1
    16'b11100010_11011011 : OUT <= 1;  //226 / 219 = 1
    16'b11100010_11011100 : OUT <= 1;  //226 / 220 = 1
    16'b11100010_11011101 : OUT <= 1;  //226 / 221 = 1
    16'b11100010_11011110 : OUT <= 1;  //226 / 222 = 1
    16'b11100010_11011111 : OUT <= 1;  //226 / 223 = 1
    16'b11100010_11100000 : OUT <= 1;  //226 / 224 = 1
    16'b11100010_11100001 : OUT <= 1;  //226 / 225 = 1
    16'b11100010_11100010 : OUT <= 1;  //226 / 226 = 1
    16'b11100010_11100011 : OUT <= 0;  //226 / 227 = 0
    16'b11100010_11100100 : OUT <= 0;  //226 / 228 = 0
    16'b11100010_11100101 : OUT <= 0;  //226 / 229 = 0
    16'b11100010_11100110 : OUT <= 0;  //226 / 230 = 0
    16'b11100010_11100111 : OUT <= 0;  //226 / 231 = 0
    16'b11100010_11101000 : OUT <= 0;  //226 / 232 = 0
    16'b11100010_11101001 : OUT <= 0;  //226 / 233 = 0
    16'b11100010_11101010 : OUT <= 0;  //226 / 234 = 0
    16'b11100010_11101011 : OUT <= 0;  //226 / 235 = 0
    16'b11100010_11101100 : OUT <= 0;  //226 / 236 = 0
    16'b11100010_11101101 : OUT <= 0;  //226 / 237 = 0
    16'b11100010_11101110 : OUT <= 0;  //226 / 238 = 0
    16'b11100010_11101111 : OUT <= 0;  //226 / 239 = 0
    16'b11100010_11110000 : OUT <= 0;  //226 / 240 = 0
    16'b11100010_11110001 : OUT <= 0;  //226 / 241 = 0
    16'b11100010_11110010 : OUT <= 0;  //226 / 242 = 0
    16'b11100010_11110011 : OUT <= 0;  //226 / 243 = 0
    16'b11100010_11110100 : OUT <= 0;  //226 / 244 = 0
    16'b11100010_11110101 : OUT <= 0;  //226 / 245 = 0
    16'b11100010_11110110 : OUT <= 0;  //226 / 246 = 0
    16'b11100010_11110111 : OUT <= 0;  //226 / 247 = 0
    16'b11100010_11111000 : OUT <= 0;  //226 / 248 = 0
    16'b11100010_11111001 : OUT <= 0;  //226 / 249 = 0
    16'b11100010_11111010 : OUT <= 0;  //226 / 250 = 0
    16'b11100010_11111011 : OUT <= 0;  //226 / 251 = 0
    16'b11100010_11111100 : OUT <= 0;  //226 / 252 = 0
    16'b11100010_11111101 : OUT <= 0;  //226 / 253 = 0
    16'b11100010_11111110 : OUT <= 0;  //226 / 254 = 0
    16'b11100010_11111111 : OUT <= 0;  //226 / 255 = 0
    16'b11100011_00000000 : OUT <= 0;  //227 / 0 = 0
    16'b11100011_00000001 : OUT <= 227;  //227 / 1 = 227
    16'b11100011_00000010 : OUT <= 113;  //227 / 2 = 113
    16'b11100011_00000011 : OUT <= 75;  //227 / 3 = 75
    16'b11100011_00000100 : OUT <= 56;  //227 / 4 = 56
    16'b11100011_00000101 : OUT <= 45;  //227 / 5 = 45
    16'b11100011_00000110 : OUT <= 37;  //227 / 6 = 37
    16'b11100011_00000111 : OUT <= 32;  //227 / 7 = 32
    16'b11100011_00001000 : OUT <= 28;  //227 / 8 = 28
    16'b11100011_00001001 : OUT <= 25;  //227 / 9 = 25
    16'b11100011_00001010 : OUT <= 22;  //227 / 10 = 22
    16'b11100011_00001011 : OUT <= 20;  //227 / 11 = 20
    16'b11100011_00001100 : OUT <= 18;  //227 / 12 = 18
    16'b11100011_00001101 : OUT <= 17;  //227 / 13 = 17
    16'b11100011_00001110 : OUT <= 16;  //227 / 14 = 16
    16'b11100011_00001111 : OUT <= 15;  //227 / 15 = 15
    16'b11100011_00010000 : OUT <= 14;  //227 / 16 = 14
    16'b11100011_00010001 : OUT <= 13;  //227 / 17 = 13
    16'b11100011_00010010 : OUT <= 12;  //227 / 18 = 12
    16'b11100011_00010011 : OUT <= 11;  //227 / 19 = 11
    16'b11100011_00010100 : OUT <= 11;  //227 / 20 = 11
    16'b11100011_00010101 : OUT <= 10;  //227 / 21 = 10
    16'b11100011_00010110 : OUT <= 10;  //227 / 22 = 10
    16'b11100011_00010111 : OUT <= 9;  //227 / 23 = 9
    16'b11100011_00011000 : OUT <= 9;  //227 / 24 = 9
    16'b11100011_00011001 : OUT <= 9;  //227 / 25 = 9
    16'b11100011_00011010 : OUT <= 8;  //227 / 26 = 8
    16'b11100011_00011011 : OUT <= 8;  //227 / 27 = 8
    16'b11100011_00011100 : OUT <= 8;  //227 / 28 = 8
    16'b11100011_00011101 : OUT <= 7;  //227 / 29 = 7
    16'b11100011_00011110 : OUT <= 7;  //227 / 30 = 7
    16'b11100011_00011111 : OUT <= 7;  //227 / 31 = 7
    16'b11100011_00100000 : OUT <= 7;  //227 / 32 = 7
    16'b11100011_00100001 : OUT <= 6;  //227 / 33 = 6
    16'b11100011_00100010 : OUT <= 6;  //227 / 34 = 6
    16'b11100011_00100011 : OUT <= 6;  //227 / 35 = 6
    16'b11100011_00100100 : OUT <= 6;  //227 / 36 = 6
    16'b11100011_00100101 : OUT <= 6;  //227 / 37 = 6
    16'b11100011_00100110 : OUT <= 5;  //227 / 38 = 5
    16'b11100011_00100111 : OUT <= 5;  //227 / 39 = 5
    16'b11100011_00101000 : OUT <= 5;  //227 / 40 = 5
    16'b11100011_00101001 : OUT <= 5;  //227 / 41 = 5
    16'b11100011_00101010 : OUT <= 5;  //227 / 42 = 5
    16'b11100011_00101011 : OUT <= 5;  //227 / 43 = 5
    16'b11100011_00101100 : OUT <= 5;  //227 / 44 = 5
    16'b11100011_00101101 : OUT <= 5;  //227 / 45 = 5
    16'b11100011_00101110 : OUT <= 4;  //227 / 46 = 4
    16'b11100011_00101111 : OUT <= 4;  //227 / 47 = 4
    16'b11100011_00110000 : OUT <= 4;  //227 / 48 = 4
    16'b11100011_00110001 : OUT <= 4;  //227 / 49 = 4
    16'b11100011_00110010 : OUT <= 4;  //227 / 50 = 4
    16'b11100011_00110011 : OUT <= 4;  //227 / 51 = 4
    16'b11100011_00110100 : OUT <= 4;  //227 / 52 = 4
    16'b11100011_00110101 : OUT <= 4;  //227 / 53 = 4
    16'b11100011_00110110 : OUT <= 4;  //227 / 54 = 4
    16'b11100011_00110111 : OUT <= 4;  //227 / 55 = 4
    16'b11100011_00111000 : OUT <= 4;  //227 / 56 = 4
    16'b11100011_00111001 : OUT <= 3;  //227 / 57 = 3
    16'b11100011_00111010 : OUT <= 3;  //227 / 58 = 3
    16'b11100011_00111011 : OUT <= 3;  //227 / 59 = 3
    16'b11100011_00111100 : OUT <= 3;  //227 / 60 = 3
    16'b11100011_00111101 : OUT <= 3;  //227 / 61 = 3
    16'b11100011_00111110 : OUT <= 3;  //227 / 62 = 3
    16'b11100011_00111111 : OUT <= 3;  //227 / 63 = 3
    16'b11100011_01000000 : OUT <= 3;  //227 / 64 = 3
    16'b11100011_01000001 : OUT <= 3;  //227 / 65 = 3
    16'b11100011_01000010 : OUT <= 3;  //227 / 66 = 3
    16'b11100011_01000011 : OUT <= 3;  //227 / 67 = 3
    16'b11100011_01000100 : OUT <= 3;  //227 / 68 = 3
    16'b11100011_01000101 : OUT <= 3;  //227 / 69 = 3
    16'b11100011_01000110 : OUT <= 3;  //227 / 70 = 3
    16'b11100011_01000111 : OUT <= 3;  //227 / 71 = 3
    16'b11100011_01001000 : OUT <= 3;  //227 / 72 = 3
    16'b11100011_01001001 : OUT <= 3;  //227 / 73 = 3
    16'b11100011_01001010 : OUT <= 3;  //227 / 74 = 3
    16'b11100011_01001011 : OUT <= 3;  //227 / 75 = 3
    16'b11100011_01001100 : OUT <= 2;  //227 / 76 = 2
    16'b11100011_01001101 : OUT <= 2;  //227 / 77 = 2
    16'b11100011_01001110 : OUT <= 2;  //227 / 78 = 2
    16'b11100011_01001111 : OUT <= 2;  //227 / 79 = 2
    16'b11100011_01010000 : OUT <= 2;  //227 / 80 = 2
    16'b11100011_01010001 : OUT <= 2;  //227 / 81 = 2
    16'b11100011_01010010 : OUT <= 2;  //227 / 82 = 2
    16'b11100011_01010011 : OUT <= 2;  //227 / 83 = 2
    16'b11100011_01010100 : OUT <= 2;  //227 / 84 = 2
    16'b11100011_01010101 : OUT <= 2;  //227 / 85 = 2
    16'b11100011_01010110 : OUT <= 2;  //227 / 86 = 2
    16'b11100011_01010111 : OUT <= 2;  //227 / 87 = 2
    16'b11100011_01011000 : OUT <= 2;  //227 / 88 = 2
    16'b11100011_01011001 : OUT <= 2;  //227 / 89 = 2
    16'b11100011_01011010 : OUT <= 2;  //227 / 90 = 2
    16'b11100011_01011011 : OUT <= 2;  //227 / 91 = 2
    16'b11100011_01011100 : OUT <= 2;  //227 / 92 = 2
    16'b11100011_01011101 : OUT <= 2;  //227 / 93 = 2
    16'b11100011_01011110 : OUT <= 2;  //227 / 94 = 2
    16'b11100011_01011111 : OUT <= 2;  //227 / 95 = 2
    16'b11100011_01100000 : OUT <= 2;  //227 / 96 = 2
    16'b11100011_01100001 : OUT <= 2;  //227 / 97 = 2
    16'b11100011_01100010 : OUT <= 2;  //227 / 98 = 2
    16'b11100011_01100011 : OUT <= 2;  //227 / 99 = 2
    16'b11100011_01100100 : OUT <= 2;  //227 / 100 = 2
    16'b11100011_01100101 : OUT <= 2;  //227 / 101 = 2
    16'b11100011_01100110 : OUT <= 2;  //227 / 102 = 2
    16'b11100011_01100111 : OUT <= 2;  //227 / 103 = 2
    16'b11100011_01101000 : OUT <= 2;  //227 / 104 = 2
    16'b11100011_01101001 : OUT <= 2;  //227 / 105 = 2
    16'b11100011_01101010 : OUT <= 2;  //227 / 106 = 2
    16'b11100011_01101011 : OUT <= 2;  //227 / 107 = 2
    16'b11100011_01101100 : OUT <= 2;  //227 / 108 = 2
    16'b11100011_01101101 : OUT <= 2;  //227 / 109 = 2
    16'b11100011_01101110 : OUT <= 2;  //227 / 110 = 2
    16'b11100011_01101111 : OUT <= 2;  //227 / 111 = 2
    16'b11100011_01110000 : OUT <= 2;  //227 / 112 = 2
    16'b11100011_01110001 : OUT <= 2;  //227 / 113 = 2
    16'b11100011_01110010 : OUT <= 1;  //227 / 114 = 1
    16'b11100011_01110011 : OUT <= 1;  //227 / 115 = 1
    16'b11100011_01110100 : OUT <= 1;  //227 / 116 = 1
    16'b11100011_01110101 : OUT <= 1;  //227 / 117 = 1
    16'b11100011_01110110 : OUT <= 1;  //227 / 118 = 1
    16'b11100011_01110111 : OUT <= 1;  //227 / 119 = 1
    16'b11100011_01111000 : OUT <= 1;  //227 / 120 = 1
    16'b11100011_01111001 : OUT <= 1;  //227 / 121 = 1
    16'b11100011_01111010 : OUT <= 1;  //227 / 122 = 1
    16'b11100011_01111011 : OUT <= 1;  //227 / 123 = 1
    16'b11100011_01111100 : OUT <= 1;  //227 / 124 = 1
    16'b11100011_01111101 : OUT <= 1;  //227 / 125 = 1
    16'b11100011_01111110 : OUT <= 1;  //227 / 126 = 1
    16'b11100011_01111111 : OUT <= 1;  //227 / 127 = 1
    16'b11100011_10000000 : OUT <= 1;  //227 / 128 = 1
    16'b11100011_10000001 : OUT <= 1;  //227 / 129 = 1
    16'b11100011_10000010 : OUT <= 1;  //227 / 130 = 1
    16'b11100011_10000011 : OUT <= 1;  //227 / 131 = 1
    16'b11100011_10000100 : OUT <= 1;  //227 / 132 = 1
    16'b11100011_10000101 : OUT <= 1;  //227 / 133 = 1
    16'b11100011_10000110 : OUT <= 1;  //227 / 134 = 1
    16'b11100011_10000111 : OUT <= 1;  //227 / 135 = 1
    16'b11100011_10001000 : OUT <= 1;  //227 / 136 = 1
    16'b11100011_10001001 : OUT <= 1;  //227 / 137 = 1
    16'b11100011_10001010 : OUT <= 1;  //227 / 138 = 1
    16'b11100011_10001011 : OUT <= 1;  //227 / 139 = 1
    16'b11100011_10001100 : OUT <= 1;  //227 / 140 = 1
    16'b11100011_10001101 : OUT <= 1;  //227 / 141 = 1
    16'b11100011_10001110 : OUT <= 1;  //227 / 142 = 1
    16'b11100011_10001111 : OUT <= 1;  //227 / 143 = 1
    16'b11100011_10010000 : OUT <= 1;  //227 / 144 = 1
    16'b11100011_10010001 : OUT <= 1;  //227 / 145 = 1
    16'b11100011_10010010 : OUT <= 1;  //227 / 146 = 1
    16'b11100011_10010011 : OUT <= 1;  //227 / 147 = 1
    16'b11100011_10010100 : OUT <= 1;  //227 / 148 = 1
    16'b11100011_10010101 : OUT <= 1;  //227 / 149 = 1
    16'b11100011_10010110 : OUT <= 1;  //227 / 150 = 1
    16'b11100011_10010111 : OUT <= 1;  //227 / 151 = 1
    16'b11100011_10011000 : OUT <= 1;  //227 / 152 = 1
    16'b11100011_10011001 : OUT <= 1;  //227 / 153 = 1
    16'b11100011_10011010 : OUT <= 1;  //227 / 154 = 1
    16'b11100011_10011011 : OUT <= 1;  //227 / 155 = 1
    16'b11100011_10011100 : OUT <= 1;  //227 / 156 = 1
    16'b11100011_10011101 : OUT <= 1;  //227 / 157 = 1
    16'b11100011_10011110 : OUT <= 1;  //227 / 158 = 1
    16'b11100011_10011111 : OUT <= 1;  //227 / 159 = 1
    16'b11100011_10100000 : OUT <= 1;  //227 / 160 = 1
    16'b11100011_10100001 : OUT <= 1;  //227 / 161 = 1
    16'b11100011_10100010 : OUT <= 1;  //227 / 162 = 1
    16'b11100011_10100011 : OUT <= 1;  //227 / 163 = 1
    16'b11100011_10100100 : OUT <= 1;  //227 / 164 = 1
    16'b11100011_10100101 : OUT <= 1;  //227 / 165 = 1
    16'b11100011_10100110 : OUT <= 1;  //227 / 166 = 1
    16'b11100011_10100111 : OUT <= 1;  //227 / 167 = 1
    16'b11100011_10101000 : OUT <= 1;  //227 / 168 = 1
    16'b11100011_10101001 : OUT <= 1;  //227 / 169 = 1
    16'b11100011_10101010 : OUT <= 1;  //227 / 170 = 1
    16'b11100011_10101011 : OUT <= 1;  //227 / 171 = 1
    16'b11100011_10101100 : OUT <= 1;  //227 / 172 = 1
    16'b11100011_10101101 : OUT <= 1;  //227 / 173 = 1
    16'b11100011_10101110 : OUT <= 1;  //227 / 174 = 1
    16'b11100011_10101111 : OUT <= 1;  //227 / 175 = 1
    16'b11100011_10110000 : OUT <= 1;  //227 / 176 = 1
    16'b11100011_10110001 : OUT <= 1;  //227 / 177 = 1
    16'b11100011_10110010 : OUT <= 1;  //227 / 178 = 1
    16'b11100011_10110011 : OUT <= 1;  //227 / 179 = 1
    16'b11100011_10110100 : OUT <= 1;  //227 / 180 = 1
    16'b11100011_10110101 : OUT <= 1;  //227 / 181 = 1
    16'b11100011_10110110 : OUT <= 1;  //227 / 182 = 1
    16'b11100011_10110111 : OUT <= 1;  //227 / 183 = 1
    16'b11100011_10111000 : OUT <= 1;  //227 / 184 = 1
    16'b11100011_10111001 : OUT <= 1;  //227 / 185 = 1
    16'b11100011_10111010 : OUT <= 1;  //227 / 186 = 1
    16'b11100011_10111011 : OUT <= 1;  //227 / 187 = 1
    16'b11100011_10111100 : OUT <= 1;  //227 / 188 = 1
    16'b11100011_10111101 : OUT <= 1;  //227 / 189 = 1
    16'b11100011_10111110 : OUT <= 1;  //227 / 190 = 1
    16'b11100011_10111111 : OUT <= 1;  //227 / 191 = 1
    16'b11100011_11000000 : OUT <= 1;  //227 / 192 = 1
    16'b11100011_11000001 : OUT <= 1;  //227 / 193 = 1
    16'b11100011_11000010 : OUT <= 1;  //227 / 194 = 1
    16'b11100011_11000011 : OUT <= 1;  //227 / 195 = 1
    16'b11100011_11000100 : OUT <= 1;  //227 / 196 = 1
    16'b11100011_11000101 : OUT <= 1;  //227 / 197 = 1
    16'b11100011_11000110 : OUT <= 1;  //227 / 198 = 1
    16'b11100011_11000111 : OUT <= 1;  //227 / 199 = 1
    16'b11100011_11001000 : OUT <= 1;  //227 / 200 = 1
    16'b11100011_11001001 : OUT <= 1;  //227 / 201 = 1
    16'b11100011_11001010 : OUT <= 1;  //227 / 202 = 1
    16'b11100011_11001011 : OUT <= 1;  //227 / 203 = 1
    16'b11100011_11001100 : OUT <= 1;  //227 / 204 = 1
    16'b11100011_11001101 : OUT <= 1;  //227 / 205 = 1
    16'b11100011_11001110 : OUT <= 1;  //227 / 206 = 1
    16'b11100011_11001111 : OUT <= 1;  //227 / 207 = 1
    16'b11100011_11010000 : OUT <= 1;  //227 / 208 = 1
    16'b11100011_11010001 : OUT <= 1;  //227 / 209 = 1
    16'b11100011_11010010 : OUT <= 1;  //227 / 210 = 1
    16'b11100011_11010011 : OUT <= 1;  //227 / 211 = 1
    16'b11100011_11010100 : OUT <= 1;  //227 / 212 = 1
    16'b11100011_11010101 : OUT <= 1;  //227 / 213 = 1
    16'b11100011_11010110 : OUT <= 1;  //227 / 214 = 1
    16'b11100011_11010111 : OUT <= 1;  //227 / 215 = 1
    16'b11100011_11011000 : OUT <= 1;  //227 / 216 = 1
    16'b11100011_11011001 : OUT <= 1;  //227 / 217 = 1
    16'b11100011_11011010 : OUT <= 1;  //227 / 218 = 1
    16'b11100011_11011011 : OUT <= 1;  //227 / 219 = 1
    16'b11100011_11011100 : OUT <= 1;  //227 / 220 = 1
    16'b11100011_11011101 : OUT <= 1;  //227 / 221 = 1
    16'b11100011_11011110 : OUT <= 1;  //227 / 222 = 1
    16'b11100011_11011111 : OUT <= 1;  //227 / 223 = 1
    16'b11100011_11100000 : OUT <= 1;  //227 / 224 = 1
    16'b11100011_11100001 : OUT <= 1;  //227 / 225 = 1
    16'b11100011_11100010 : OUT <= 1;  //227 / 226 = 1
    16'b11100011_11100011 : OUT <= 1;  //227 / 227 = 1
    16'b11100011_11100100 : OUT <= 0;  //227 / 228 = 0
    16'b11100011_11100101 : OUT <= 0;  //227 / 229 = 0
    16'b11100011_11100110 : OUT <= 0;  //227 / 230 = 0
    16'b11100011_11100111 : OUT <= 0;  //227 / 231 = 0
    16'b11100011_11101000 : OUT <= 0;  //227 / 232 = 0
    16'b11100011_11101001 : OUT <= 0;  //227 / 233 = 0
    16'b11100011_11101010 : OUT <= 0;  //227 / 234 = 0
    16'b11100011_11101011 : OUT <= 0;  //227 / 235 = 0
    16'b11100011_11101100 : OUT <= 0;  //227 / 236 = 0
    16'b11100011_11101101 : OUT <= 0;  //227 / 237 = 0
    16'b11100011_11101110 : OUT <= 0;  //227 / 238 = 0
    16'b11100011_11101111 : OUT <= 0;  //227 / 239 = 0
    16'b11100011_11110000 : OUT <= 0;  //227 / 240 = 0
    16'b11100011_11110001 : OUT <= 0;  //227 / 241 = 0
    16'b11100011_11110010 : OUT <= 0;  //227 / 242 = 0
    16'b11100011_11110011 : OUT <= 0;  //227 / 243 = 0
    16'b11100011_11110100 : OUT <= 0;  //227 / 244 = 0
    16'b11100011_11110101 : OUT <= 0;  //227 / 245 = 0
    16'b11100011_11110110 : OUT <= 0;  //227 / 246 = 0
    16'b11100011_11110111 : OUT <= 0;  //227 / 247 = 0
    16'b11100011_11111000 : OUT <= 0;  //227 / 248 = 0
    16'b11100011_11111001 : OUT <= 0;  //227 / 249 = 0
    16'b11100011_11111010 : OUT <= 0;  //227 / 250 = 0
    16'b11100011_11111011 : OUT <= 0;  //227 / 251 = 0
    16'b11100011_11111100 : OUT <= 0;  //227 / 252 = 0
    16'b11100011_11111101 : OUT <= 0;  //227 / 253 = 0
    16'b11100011_11111110 : OUT <= 0;  //227 / 254 = 0
    16'b11100011_11111111 : OUT <= 0;  //227 / 255 = 0
    16'b11100100_00000000 : OUT <= 0;  //228 / 0 = 0
    16'b11100100_00000001 : OUT <= 228;  //228 / 1 = 228
    16'b11100100_00000010 : OUT <= 114;  //228 / 2 = 114
    16'b11100100_00000011 : OUT <= 76;  //228 / 3 = 76
    16'b11100100_00000100 : OUT <= 57;  //228 / 4 = 57
    16'b11100100_00000101 : OUT <= 45;  //228 / 5 = 45
    16'b11100100_00000110 : OUT <= 38;  //228 / 6 = 38
    16'b11100100_00000111 : OUT <= 32;  //228 / 7 = 32
    16'b11100100_00001000 : OUT <= 28;  //228 / 8 = 28
    16'b11100100_00001001 : OUT <= 25;  //228 / 9 = 25
    16'b11100100_00001010 : OUT <= 22;  //228 / 10 = 22
    16'b11100100_00001011 : OUT <= 20;  //228 / 11 = 20
    16'b11100100_00001100 : OUT <= 19;  //228 / 12 = 19
    16'b11100100_00001101 : OUT <= 17;  //228 / 13 = 17
    16'b11100100_00001110 : OUT <= 16;  //228 / 14 = 16
    16'b11100100_00001111 : OUT <= 15;  //228 / 15 = 15
    16'b11100100_00010000 : OUT <= 14;  //228 / 16 = 14
    16'b11100100_00010001 : OUT <= 13;  //228 / 17 = 13
    16'b11100100_00010010 : OUT <= 12;  //228 / 18 = 12
    16'b11100100_00010011 : OUT <= 12;  //228 / 19 = 12
    16'b11100100_00010100 : OUT <= 11;  //228 / 20 = 11
    16'b11100100_00010101 : OUT <= 10;  //228 / 21 = 10
    16'b11100100_00010110 : OUT <= 10;  //228 / 22 = 10
    16'b11100100_00010111 : OUT <= 9;  //228 / 23 = 9
    16'b11100100_00011000 : OUT <= 9;  //228 / 24 = 9
    16'b11100100_00011001 : OUT <= 9;  //228 / 25 = 9
    16'b11100100_00011010 : OUT <= 8;  //228 / 26 = 8
    16'b11100100_00011011 : OUT <= 8;  //228 / 27 = 8
    16'b11100100_00011100 : OUT <= 8;  //228 / 28 = 8
    16'b11100100_00011101 : OUT <= 7;  //228 / 29 = 7
    16'b11100100_00011110 : OUT <= 7;  //228 / 30 = 7
    16'b11100100_00011111 : OUT <= 7;  //228 / 31 = 7
    16'b11100100_00100000 : OUT <= 7;  //228 / 32 = 7
    16'b11100100_00100001 : OUT <= 6;  //228 / 33 = 6
    16'b11100100_00100010 : OUT <= 6;  //228 / 34 = 6
    16'b11100100_00100011 : OUT <= 6;  //228 / 35 = 6
    16'b11100100_00100100 : OUT <= 6;  //228 / 36 = 6
    16'b11100100_00100101 : OUT <= 6;  //228 / 37 = 6
    16'b11100100_00100110 : OUT <= 6;  //228 / 38 = 6
    16'b11100100_00100111 : OUT <= 5;  //228 / 39 = 5
    16'b11100100_00101000 : OUT <= 5;  //228 / 40 = 5
    16'b11100100_00101001 : OUT <= 5;  //228 / 41 = 5
    16'b11100100_00101010 : OUT <= 5;  //228 / 42 = 5
    16'b11100100_00101011 : OUT <= 5;  //228 / 43 = 5
    16'b11100100_00101100 : OUT <= 5;  //228 / 44 = 5
    16'b11100100_00101101 : OUT <= 5;  //228 / 45 = 5
    16'b11100100_00101110 : OUT <= 4;  //228 / 46 = 4
    16'b11100100_00101111 : OUT <= 4;  //228 / 47 = 4
    16'b11100100_00110000 : OUT <= 4;  //228 / 48 = 4
    16'b11100100_00110001 : OUT <= 4;  //228 / 49 = 4
    16'b11100100_00110010 : OUT <= 4;  //228 / 50 = 4
    16'b11100100_00110011 : OUT <= 4;  //228 / 51 = 4
    16'b11100100_00110100 : OUT <= 4;  //228 / 52 = 4
    16'b11100100_00110101 : OUT <= 4;  //228 / 53 = 4
    16'b11100100_00110110 : OUT <= 4;  //228 / 54 = 4
    16'b11100100_00110111 : OUT <= 4;  //228 / 55 = 4
    16'b11100100_00111000 : OUT <= 4;  //228 / 56 = 4
    16'b11100100_00111001 : OUT <= 4;  //228 / 57 = 4
    16'b11100100_00111010 : OUT <= 3;  //228 / 58 = 3
    16'b11100100_00111011 : OUT <= 3;  //228 / 59 = 3
    16'b11100100_00111100 : OUT <= 3;  //228 / 60 = 3
    16'b11100100_00111101 : OUT <= 3;  //228 / 61 = 3
    16'b11100100_00111110 : OUT <= 3;  //228 / 62 = 3
    16'b11100100_00111111 : OUT <= 3;  //228 / 63 = 3
    16'b11100100_01000000 : OUT <= 3;  //228 / 64 = 3
    16'b11100100_01000001 : OUT <= 3;  //228 / 65 = 3
    16'b11100100_01000010 : OUT <= 3;  //228 / 66 = 3
    16'b11100100_01000011 : OUT <= 3;  //228 / 67 = 3
    16'b11100100_01000100 : OUT <= 3;  //228 / 68 = 3
    16'b11100100_01000101 : OUT <= 3;  //228 / 69 = 3
    16'b11100100_01000110 : OUT <= 3;  //228 / 70 = 3
    16'b11100100_01000111 : OUT <= 3;  //228 / 71 = 3
    16'b11100100_01001000 : OUT <= 3;  //228 / 72 = 3
    16'b11100100_01001001 : OUT <= 3;  //228 / 73 = 3
    16'b11100100_01001010 : OUT <= 3;  //228 / 74 = 3
    16'b11100100_01001011 : OUT <= 3;  //228 / 75 = 3
    16'b11100100_01001100 : OUT <= 3;  //228 / 76 = 3
    16'b11100100_01001101 : OUT <= 2;  //228 / 77 = 2
    16'b11100100_01001110 : OUT <= 2;  //228 / 78 = 2
    16'b11100100_01001111 : OUT <= 2;  //228 / 79 = 2
    16'b11100100_01010000 : OUT <= 2;  //228 / 80 = 2
    16'b11100100_01010001 : OUT <= 2;  //228 / 81 = 2
    16'b11100100_01010010 : OUT <= 2;  //228 / 82 = 2
    16'b11100100_01010011 : OUT <= 2;  //228 / 83 = 2
    16'b11100100_01010100 : OUT <= 2;  //228 / 84 = 2
    16'b11100100_01010101 : OUT <= 2;  //228 / 85 = 2
    16'b11100100_01010110 : OUT <= 2;  //228 / 86 = 2
    16'b11100100_01010111 : OUT <= 2;  //228 / 87 = 2
    16'b11100100_01011000 : OUT <= 2;  //228 / 88 = 2
    16'b11100100_01011001 : OUT <= 2;  //228 / 89 = 2
    16'b11100100_01011010 : OUT <= 2;  //228 / 90 = 2
    16'b11100100_01011011 : OUT <= 2;  //228 / 91 = 2
    16'b11100100_01011100 : OUT <= 2;  //228 / 92 = 2
    16'b11100100_01011101 : OUT <= 2;  //228 / 93 = 2
    16'b11100100_01011110 : OUT <= 2;  //228 / 94 = 2
    16'b11100100_01011111 : OUT <= 2;  //228 / 95 = 2
    16'b11100100_01100000 : OUT <= 2;  //228 / 96 = 2
    16'b11100100_01100001 : OUT <= 2;  //228 / 97 = 2
    16'b11100100_01100010 : OUT <= 2;  //228 / 98 = 2
    16'b11100100_01100011 : OUT <= 2;  //228 / 99 = 2
    16'b11100100_01100100 : OUT <= 2;  //228 / 100 = 2
    16'b11100100_01100101 : OUT <= 2;  //228 / 101 = 2
    16'b11100100_01100110 : OUT <= 2;  //228 / 102 = 2
    16'b11100100_01100111 : OUT <= 2;  //228 / 103 = 2
    16'b11100100_01101000 : OUT <= 2;  //228 / 104 = 2
    16'b11100100_01101001 : OUT <= 2;  //228 / 105 = 2
    16'b11100100_01101010 : OUT <= 2;  //228 / 106 = 2
    16'b11100100_01101011 : OUT <= 2;  //228 / 107 = 2
    16'b11100100_01101100 : OUT <= 2;  //228 / 108 = 2
    16'b11100100_01101101 : OUT <= 2;  //228 / 109 = 2
    16'b11100100_01101110 : OUT <= 2;  //228 / 110 = 2
    16'b11100100_01101111 : OUT <= 2;  //228 / 111 = 2
    16'b11100100_01110000 : OUT <= 2;  //228 / 112 = 2
    16'b11100100_01110001 : OUT <= 2;  //228 / 113 = 2
    16'b11100100_01110010 : OUT <= 2;  //228 / 114 = 2
    16'b11100100_01110011 : OUT <= 1;  //228 / 115 = 1
    16'b11100100_01110100 : OUT <= 1;  //228 / 116 = 1
    16'b11100100_01110101 : OUT <= 1;  //228 / 117 = 1
    16'b11100100_01110110 : OUT <= 1;  //228 / 118 = 1
    16'b11100100_01110111 : OUT <= 1;  //228 / 119 = 1
    16'b11100100_01111000 : OUT <= 1;  //228 / 120 = 1
    16'b11100100_01111001 : OUT <= 1;  //228 / 121 = 1
    16'b11100100_01111010 : OUT <= 1;  //228 / 122 = 1
    16'b11100100_01111011 : OUT <= 1;  //228 / 123 = 1
    16'b11100100_01111100 : OUT <= 1;  //228 / 124 = 1
    16'b11100100_01111101 : OUT <= 1;  //228 / 125 = 1
    16'b11100100_01111110 : OUT <= 1;  //228 / 126 = 1
    16'b11100100_01111111 : OUT <= 1;  //228 / 127 = 1
    16'b11100100_10000000 : OUT <= 1;  //228 / 128 = 1
    16'b11100100_10000001 : OUT <= 1;  //228 / 129 = 1
    16'b11100100_10000010 : OUT <= 1;  //228 / 130 = 1
    16'b11100100_10000011 : OUT <= 1;  //228 / 131 = 1
    16'b11100100_10000100 : OUT <= 1;  //228 / 132 = 1
    16'b11100100_10000101 : OUT <= 1;  //228 / 133 = 1
    16'b11100100_10000110 : OUT <= 1;  //228 / 134 = 1
    16'b11100100_10000111 : OUT <= 1;  //228 / 135 = 1
    16'b11100100_10001000 : OUT <= 1;  //228 / 136 = 1
    16'b11100100_10001001 : OUT <= 1;  //228 / 137 = 1
    16'b11100100_10001010 : OUT <= 1;  //228 / 138 = 1
    16'b11100100_10001011 : OUT <= 1;  //228 / 139 = 1
    16'b11100100_10001100 : OUT <= 1;  //228 / 140 = 1
    16'b11100100_10001101 : OUT <= 1;  //228 / 141 = 1
    16'b11100100_10001110 : OUT <= 1;  //228 / 142 = 1
    16'b11100100_10001111 : OUT <= 1;  //228 / 143 = 1
    16'b11100100_10010000 : OUT <= 1;  //228 / 144 = 1
    16'b11100100_10010001 : OUT <= 1;  //228 / 145 = 1
    16'b11100100_10010010 : OUT <= 1;  //228 / 146 = 1
    16'b11100100_10010011 : OUT <= 1;  //228 / 147 = 1
    16'b11100100_10010100 : OUT <= 1;  //228 / 148 = 1
    16'b11100100_10010101 : OUT <= 1;  //228 / 149 = 1
    16'b11100100_10010110 : OUT <= 1;  //228 / 150 = 1
    16'b11100100_10010111 : OUT <= 1;  //228 / 151 = 1
    16'b11100100_10011000 : OUT <= 1;  //228 / 152 = 1
    16'b11100100_10011001 : OUT <= 1;  //228 / 153 = 1
    16'b11100100_10011010 : OUT <= 1;  //228 / 154 = 1
    16'b11100100_10011011 : OUT <= 1;  //228 / 155 = 1
    16'b11100100_10011100 : OUT <= 1;  //228 / 156 = 1
    16'b11100100_10011101 : OUT <= 1;  //228 / 157 = 1
    16'b11100100_10011110 : OUT <= 1;  //228 / 158 = 1
    16'b11100100_10011111 : OUT <= 1;  //228 / 159 = 1
    16'b11100100_10100000 : OUT <= 1;  //228 / 160 = 1
    16'b11100100_10100001 : OUT <= 1;  //228 / 161 = 1
    16'b11100100_10100010 : OUT <= 1;  //228 / 162 = 1
    16'b11100100_10100011 : OUT <= 1;  //228 / 163 = 1
    16'b11100100_10100100 : OUT <= 1;  //228 / 164 = 1
    16'b11100100_10100101 : OUT <= 1;  //228 / 165 = 1
    16'b11100100_10100110 : OUT <= 1;  //228 / 166 = 1
    16'b11100100_10100111 : OUT <= 1;  //228 / 167 = 1
    16'b11100100_10101000 : OUT <= 1;  //228 / 168 = 1
    16'b11100100_10101001 : OUT <= 1;  //228 / 169 = 1
    16'b11100100_10101010 : OUT <= 1;  //228 / 170 = 1
    16'b11100100_10101011 : OUT <= 1;  //228 / 171 = 1
    16'b11100100_10101100 : OUT <= 1;  //228 / 172 = 1
    16'b11100100_10101101 : OUT <= 1;  //228 / 173 = 1
    16'b11100100_10101110 : OUT <= 1;  //228 / 174 = 1
    16'b11100100_10101111 : OUT <= 1;  //228 / 175 = 1
    16'b11100100_10110000 : OUT <= 1;  //228 / 176 = 1
    16'b11100100_10110001 : OUT <= 1;  //228 / 177 = 1
    16'b11100100_10110010 : OUT <= 1;  //228 / 178 = 1
    16'b11100100_10110011 : OUT <= 1;  //228 / 179 = 1
    16'b11100100_10110100 : OUT <= 1;  //228 / 180 = 1
    16'b11100100_10110101 : OUT <= 1;  //228 / 181 = 1
    16'b11100100_10110110 : OUT <= 1;  //228 / 182 = 1
    16'b11100100_10110111 : OUT <= 1;  //228 / 183 = 1
    16'b11100100_10111000 : OUT <= 1;  //228 / 184 = 1
    16'b11100100_10111001 : OUT <= 1;  //228 / 185 = 1
    16'b11100100_10111010 : OUT <= 1;  //228 / 186 = 1
    16'b11100100_10111011 : OUT <= 1;  //228 / 187 = 1
    16'b11100100_10111100 : OUT <= 1;  //228 / 188 = 1
    16'b11100100_10111101 : OUT <= 1;  //228 / 189 = 1
    16'b11100100_10111110 : OUT <= 1;  //228 / 190 = 1
    16'b11100100_10111111 : OUT <= 1;  //228 / 191 = 1
    16'b11100100_11000000 : OUT <= 1;  //228 / 192 = 1
    16'b11100100_11000001 : OUT <= 1;  //228 / 193 = 1
    16'b11100100_11000010 : OUT <= 1;  //228 / 194 = 1
    16'b11100100_11000011 : OUT <= 1;  //228 / 195 = 1
    16'b11100100_11000100 : OUT <= 1;  //228 / 196 = 1
    16'b11100100_11000101 : OUT <= 1;  //228 / 197 = 1
    16'b11100100_11000110 : OUT <= 1;  //228 / 198 = 1
    16'b11100100_11000111 : OUT <= 1;  //228 / 199 = 1
    16'b11100100_11001000 : OUT <= 1;  //228 / 200 = 1
    16'b11100100_11001001 : OUT <= 1;  //228 / 201 = 1
    16'b11100100_11001010 : OUT <= 1;  //228 / 202 = 1
    16'b11100100_11001011 : OUT <= 1;  //228 / 203 = 1
    16'b11100100_11001100 : OUT <= 1;  //228 / 204 = 1
    16'b11100100_11001101 : OUT <= 1;  //228 / 205 = 1
    16'b11100100_11001110 : OUT <= 1;  //228 / 206 = 1
    16'b11100100_11001111 : OUT <= 1;  //228 / 207 = 1
    16'b11100100_11010000 : OUT <= 1;  //228 / 208 = 1
    16'b11100100_11010001 : OUT <= 1;  //228 / 209 = 1
    16'b11100100_11010010 : OUT <= 1;  //228 / 210 = 1
    16'b11100100_11010011 : OUT <= 1;  //228 / 211 = 1
    16'b11100100_11010100 : OUT <= 1;  //228 / 212 = 1
    16'b11100100_11010101 : OUT <= 1;  //228 / 213 = 1
    16'b11100100_11010110 : OUT <= 1;  //228 / 214 = 1
    16'b11100100_11010111 : OUT <= 1;  //228 / 215 = 1
    16'b11100100_11011000 : OUT <= 1;  //228 / 216 = 1
    16'b11100100_11011001 : OUT <= 1;  //228 / 217 = 1
    16'b11100100_11011010 : OUT <= 1;  //228 / 218 = 1
    16'b11100100_11011011 : OUT <= 1;  //228 / 219 = 1
    16'b11100100_11011100 : OUT <= 1;  //228 / 220 = 1
    16'b11100100_11011101 : OUT <= 1;  //228 / 221 = 1
    16'b11100100_11011110 : OUT <= 1;  //228 / 222 = 1
    16'b11100100_11011111 : OUT <= 1;  //228 / 223 = 1
    16'b11100100_11100000 : OUT <= 1;  //228 / 224 = 1
    16'b11100100_11100001 : OUT <= 1;  //228 / 225 = 1
    16'b11100100_11100010 : OUT <= 1;  //228 / 226 = 1
    16'b11100100_11100011 : OUT <= 1;  //228 / 227 = 1
    16'b11100100_11100100 : OUT <= 1;  //228 / 228 = 1
    16'b11100100_11100101 : OUT <= 0;  //228 / 229 = 0
    16'b11100100_11100110 : OUT <= 0;  //228 / 230 = 0
    16'b11100100_11100111 : OUT <= 0;  //228 / 231 = 0
    16'b11100100_11101000 : OUT <= 0;  //228 / 232 = 0
    16'b11100100_11101001 : OUT <= 0;  //228 / 233 = 0
    16'b11100100_11101010 : OUT <= 0;  //228 / 234 = 0
    16'b11100100_11101011 : OUT <= 0;  //228 / 235 = 0
    16'b11100100_11101100 : OUT <= 0;  //228 / 236 = 0
    16'b11100100_11101101 : OUT <= 0;  //228 / 237 = 0
    16'b11100100_11101110 : OUT <= 0;  //228 / 238 = 0
    16'b11100100_11101111 : OUT <= 0;  //228 / 239 = 0
    16'b11100100_11110000 : OUT <= 0;  //228 / 240 = 0
    16'b11100100_11110001 : OUT <= 0;  //228 / 241 = 0
    16'b11100100_11110010 : OUT <= 0;  //228 / 242 = 0
    16'b11100100_11110011 : OUT <= 0;  //228 / 243 = 0
    16'b11100100_11110100 : OUT <= 0;  //228 / 244 = 0
    16'b11100100_11110101 : OUT <= 0;  //228 / 245 = 0
    16'b11100100_11110110 : OUT <= 0;  //228 / 246 = 0
    16'b11100100_11110111 : OUT <= 0;  //228 / 247 = 0
    16'b11100100_11111000 : OUT <= 0;  //228 / 248 = 0
    16'b11100100_11111001 : OUT <= 0;  //228 / 249 = 0
    16'b11100100_11111010 : OUT <= 0;  //228 / 250 = 0
    16'b11100100_11111011 : OUT <= 0;  //228 / 251 = 0
    16'b11100100_11111100 : OUT <= 0;  //228 / 252 = 0
    16'b11100100_11111101 : OUT <= 0;  //228 / 253 = 0
    16'b11100100_11111110 : OUT <= 0;  //228 / 254 = 0
    16'b11100100_11111111 : OUT <= 0;  //228 / 255 = 0
    16'b11100101_00000000 : OUT <= 0;  //229 / 0 = 0
    16'b11100101_00000001 : OUT <= 229;  //229 / 1 = 229
    16'b11100101_00000010 : OUT <= 114;  //229 / 2 = 114
    16'b11100101_00000011 : OUT <= 76;  //229 / 3 = 76
    16'b11100101_00000100 : OUT <= 57;  //229 / 4 = 57
    16'b11100101_00000101 : OUT <= 45;  //229 / 5 = 45
    16'b11100101_00000110 : OUT <= 38;  //229 / 6 = 38
    16'b11100101_00000111 : OUT <= 32;  //229 / 7 = 32
    16'b11100101_00001000 : OUT <= 28;  //229 / 8 = 28
    16'b11100101_00001001 : OUT <= 25;  //229 / 9 = 25
    16'b11100101_00001010 : OUT <= 22;  //229 / 10 = 22
    16'b11100101_00001011 : OUT <= 20;  //229 / 11 = 20
    16'b11100101_00001100 : OUT <= 19;  //229 / 12 = 19
    16'b11100101_00001101 : OUT <= 17;  //229 / 13 = 17
    16'b11100101_00001110 : OUT <= 16;  //229 / 14 = 16
    16'b11100101_00001111 : OUT <= 15;  //229 / 15 = 15
    16'b11100101_00010000 : OUT <= 14;  //229 / 16 = 14
    16'b11100101_00010001 : OUT <= 13;  //229 / 17 = 13
    16'b11100101_00010010 : OUT <= 12;  //229 / 18 = 12
    16'b11100101_00010011 : OUT <= 12;  //229 / 19 = 12
    16'b11100101_00010100 : OUT <= 11;  //229 / 20 = 11
    16'b11100101_00010101 : OUT <= 10;  //229 / 21 = 10
    16'b11100101_00010110 : OUT <= 10;  //229 / 22 = 10
    16'b11100101_00010111 : OUT <= 9;  //229 / 23 = 9
    16'b11100101_00011000 : OUT <= 9;  //229 / 24 = 9
    16'b11100101_00011001 : OUT <= 9;  //229 / 25 = 9
    16'b11100101_00011010 : OUT <= 8;  //229 / 26 = 8
    16'b11100101_00011011 : OUT <= 8;  //229 / 27 = 8
    16'b11100101_00011100 : OUT <= 8;  //229 / 28 = 8
    16'b11100101_00011101 : OUT <= 7;  //229 / 29 = 7
    16'b11100101_00011110 : OUT <= 7;  //229 / 30 = 7
    16'b11100101_00011111 : OUT <= 7;  //229 / 31 = 7
    16'b11100101_00100000 : OUT <= 7;  //229 / 32 = 7
    16'b11100101_00100001 : OUT <= 6;  //229 / 33 = 6
    16'b11100101_00100010 : OUT <= 6;  //229 / 34 = 6
    16'b11100101_00100011 : OUT <= 6;  //229 / 35 = 6
    16'b11100101_00100100 : OUT <= 6;  //229 / 36 = 6
    16'b11100101_00100101 : OUT <= 6;  //229 / 37 = 6
    16'b11100101_00100110 : OUT <= 6;  //229 / 38 = 6
    16'b11100101_00100111 : OUT <= 5;  //229 / 39 = 5
    16'b11100101_00101000 : OUT <= 5;  //229 / 40 = 5
    16'b11100101_00101001 : OUT <= 5;  //229 / 41 = 5
    16'b11100101_00101010 : OUT <= 5;  //229 / 42 = 5
    16'b11100101_00101011 : OUT <= 5;  //229 / 43 = 5
    16'b11100101_00101100 : OUT <= 5;  //229 / 44 = 5
    16'b11100101_00101101 : OUT <= 5;  //229 / 45 = 5
    16'b11100101_00101110 : OUT <= 4;  //229 / 46 = 4
    16'b11100101_00101111 : OUT <= 4;  //229 / 47 = 4
    16'b11100101_00110000 : OUT <= 4;  //229 / 48 = 4
    16'b11100101_00110001 : OUT <= 4;  //229 / 49 = 4
    16'b11100101_00110010 : OUT <= 4;  //229 / 50 = 4
    16'b11100101_00110011 : OUT <= 4;  //229 / 51 = 4
    16'b11100101_00110100 : OUT <= 4;  //229 / 52 = 4
    16'b11100101_00110101 : OUT <= 4;  //229 / 53 = 4
    16'b11100101_00110110 : OUT <= 4;  //229 / 54 = 4
    16'b11100101_00110111 : OUT <= 4;  //229 / 55 = 4
    16'b11100101_00111000 : OUT <= 4;  //229 / 56 = 4
    16'b11100101_00111001 : OUT <= 4;  //229 / 57 = 4
    16'b11100101_00111010 : OUT <= 3;  //229 / 58 = 3
    16'b11100101_00111011 : OUT <= 3;  //229 / 59 = 3
    16'b11100101_00111100 : OUT <= 3;  //229 / 60 = 3
    16'b11100101_00111101 : OUT <= 3;  //229 / 61 = 3
    16'b11100101_00111110 : OUT <= 3;  //229 / 62 = 3
    16'b11100101_00111111 : OUT <= 3;  //229 / 63 = 3
    16'b11100101_01000000 : OUT <= 3;  //229 / 64 = 3
    16'b11100101_01000001 : OUT <= 3;  //229 / 65 = 3
    16'b11100101_01000010 : OUT <= 3;  //229 / 66 = 3
    16'b11100101_01000011 : OUT <= 3;  //229 / 67 = 3
    16'b11100101_01000100 : OUT <= 3;  //229 / 68 = 3
    16'b11100101_01000101 : OUT <= 3;  //229 / 69 = 3
    16'b11100101_01000110 : OUT <= 3;  //229 / 70 = 3
    16'b11100101_01000111 : OUT <= 3;  //229 / 71 = 3
    16'b11100101_01001000 : OUT <= 3;  //229 / 72 = 3
    16'b11100101_01001001 : OUT <= 3;  //229 / 73 = 3
    16'b11100101_01001010 : OUT <= 3;  //229 / 74 = 3
    16'b11100101_01001011 : OUT <= 3;  //229 / 75 = 3
    16'b11100101_01001100 : OUT <= 3;  //229 / 76 = 3
    16'b11100101_01001101 : OUT <= 2;  //229 / 77 = 2
    16'b11100101_01001110 : OUT <= 2;  //229 / 78 = 2
    16'b11100101_01001111 : OUT <= 2;  //229 / 79 = 2
    16'b11100101_01010000 : OUT <= 2;  //229 / 80 = 2
    16'b11100101_01010001 : OUT <= 2;  //229 / 81 = 2
    16'b11100101_01010010 : OUT <= 2;  //229 / 82 = 2
    16'b11100101_01010011 : OUT <= 2;  //229 / 83 = 2
    16'b11100101_01010100 : OUT <= 2;  //229 / 84 = 2
    16'b11100101_01010101 : OUT <= 2;  //229 / 85 = 2
    16'b11100101_01010110 : OUT <= 2;  //229 / 86 = 2
    16'b11100101_01010111 : OUT <= 2;  //229 / 87 = 2
    16'b11100101_01011000 : OUT <= 2;  //229 / 88 = 2
    16'b11100101_01011001 : OUT <= 2;  //229 / 89 = 2
    16'b11100101_01011010 : OUT <= 2;  //229 / 90 = 2
    16'b11100101_01011011 : OUT <= 2;  //229 / 91 = 2
    16'b11100101_01011100 : OUT <= 2;  //229 / 92 = 2
    16'b11100101_01011101 : OUT <= 2;  //229 / 93 = 2
    16'b11100101_01011110 : OUT <= 2;  //229 / 94 = 2
    16'b11100101_01011111 : OUT <= 2;  //229 / 95 = 2
    16'b11100101_01100000 : OUT <= 2;  //229 / 96 = 2
    16'b11100101_01100001 : OUT <= 2;  //229 / 97 = 2
    16'b11100101_01100010 : OUT <= 2;  //229 / 98 = 2
    16'b11100101_01100011 : OUT <= 2;  //229 / 99 = 2
    16'b11100101_01100100 : OUT <= 2;  //229 / 100 = 2
    16'b11100101_01100101 : OUT <= 2;  //229 / 101 = 2
    16'b11100101_01100110 : OUT <= 2;  //229 / 102 = 2
    16'b11100101_01100111 : OUT <= 2;  //229 / 103 = 2
    16'b11100101_01101000 : OUT <= 2;  //229 / 104 = 2
    16'b11100101_01101001 : OUT <= 2;  //229 / 105 = 2
    16'b11100101_01101010 : OUT <= 2;  //229 / 106 = 2
    16'b11100101_01101011 : OUT <= 2;  //229 / 107 = 2
    16'b11100101_01101100 : OUT <= 2;  //229 / 108 = 2
    16'b11100101_01101101 : OUT <= 2;  //229 / 109 = 2
    16'b11100101_01101110 : OUT <= 2;  //229 / 110 = 2
    16'b11100101_01101111 : OUT <= 2;  //229 / 111 = 2
    16'b11100101_01110000 : OUT <= 2;  //229 / 112 = 2
    16'b11100101_01110001 : OUT <= 2;  //229 / 113 = 2
    16'b11100101_01110010 : OUT <= 2;  //229 / 114 = 2
    16'b11100101_01110011 : OUT <= 1;  //229 / 115 = 1
    16'b11100101_01110100 : OUT <= 1;  //229 / 116 = 1
    16'b11100101_01110101 : OUT <= 1;  //229 / 117 = 1
    16'b11100101_01110110 : OUT <= 1;  //229 / 118 = 1
    16'b11100101_01110111 : OUT <= 1;  //229 / 119 = 1
    16'b11100101_01111000 : OUT <= 1;  //229 / 120 = 1
    16'b11100101_01111001 : OUT <= 1;  //229 / 121 = 1
    16'b11100101_01111010 : OUT <= 1;  //229 / 122 = 1
    16'b11100101_01111011 : OUT <= 1;  //229 / 123 = 1
    16'b11100101_01111100 : OUT <= 1;  //229 / 124 = 1
    16'b11100101_01111101 : OUT <= 1;  //229 / 125 = 1
    16'b11100101_01111110 : OUT <= 1;  //229 / 126 = 1
    16'b11100101_01111111 : OUT <= 1;  //229 / 127 = 1
    16'b11100101_10000000 : OUT <= 1;  //229 / 128 = 1
    16'b11100101_10000001 : OUT <= 1;  //229 / 129 = 1
    16'b11100101_10000010 : OUT <= 1;  //229 / 130 = 1
    16'b11100101_10000011 : OUT <= 1;  //229 / 131 = 1
    16'b11100101_10000100 : OUT <= 1;  //229 / 132 = 1
    16'b11100101_10000101 : OUT <= 1;  //229 / 133 = 1
    16'b11100101_10000110 : OUT <= 1;  //229 / 134 = 1
    16'b11100101_10000111 : OUT <= 1;  //229 / 135 = 1
    16'b11100101_10001000 : OUT <= 1;  //229 / 136 = 1
    16'b11100101_10001001 : OUT <= 1;  //229 / 137 = 1
    16'b11100101_10001010 : OUT <= 1;  //229 / 138 = 1
    16'b11100101_10001011 : OUT <= 1;  //229 / 139 = 1
    16'b11100101_10001100 : OUT <= 1;  //229 / 140 = 1
    16'b11100101_10001101 : OUT <= 1;  //229 / 141 = 1
    16'b11100101_10001110 : OUT <= 1;  //229 / 142 = 1
    16'b11100101_10001111 : OUT <= 1;  //229 / 143 = 1
    16'b11100101_10010000 : OUT <= 1;  //229 / 144 = 1
    16'b11100101_10010001 : OUT <= 1;  //229 / 145 = 1
    16'b11100101_10010010 : OUT <= 1;  //229 / 146 = 1
    16'b11100101_10010011 : OUT <= 1;  //229 / 147 = 1
    16'b11100101_10010100 : OUT <= 1;  //229 / 148 = 1
    16'b11100101_10010101 : OUT <= 1;  //229 / 149 = 1
    16'b11100101_10010110 : OUT <= 1;  //229 / 150 = 1
    16'b11100101_10010111 : OUT <= 1;  //229 / 151 = 1
    16'b11100101_10011000 : OUT <= 1;  //229 / 152 = 1
    16'b11100101_10011001 : OUT <= 1;  //229 / 153 = 1
    16'b11100101_10011010 : OUT <= 1;  //229 / 154 = 1
    16'b11100101_10011011 : OUT <= 1;  //229 / 155 = 1
    16'b11100101_10011100 : OUT <= 1;  //229 / 156 = 1
    16'b11100101_10011101 : OUT <= 1;  //229 / 157 = 1
    16'b11100101_10011110 : OUT <= 1;  //229 / 158 = 1
    16'b11100101_10011111 : OUT <= 1;  //229 / 159 = 1
    16'b11100101_10100000 : OUT <= 1;  //229 / 160 = 1
    16'b11100101_10100001 : OUT <= 1;  //229 / 161 = 1
    16'b11100101_10100010 : OUT <= 1;  //229 / 162 = 1
    16'b11100101_10100011 : OUT <= 1;  //229 / 163 = 1
    16'b11100101_10100100 : OUT <= 1;  //229 / 164 = 1
    16'b11100101_10100101 : OUT <= 1;  //229 / 165 = 1
    16'b11100101_10100110 : OUT <= 1;  //229 / 166 = 1
    16'b11100101_10100111 : OUT <= 1;  //229 / 167 = 1
    16'b11100101_10101000 : OUT <= 1;  //229 / 168 = 1
    16'b11100101_10101001 : OUT <= 1;  //229 / 169 = 1
    16'b11100101_10101010 : OUT <= 1;  //229 / 170 = 1
    16'b11100101_10101011 : OUT <= 1;  //229 / 171 = 1
    16'b11100101_10101100 : OUT <= 1;  //229 / 172 = 1
    16'b11100101_10101101 : OUT <= 1;  //229 / 173 = 1
    16'b11100101_10101110 : OUT <= 1;  //229 / 174 = 1
    16'b11100101_10101111 : OUT <= 1;  //229 / 175 = 1
    16'b11100101_10110000 : OUT <= 1;  //229 / 176 = 1
    16'b11100101_10110001 : OUT <= 1;  //229 / 177 = 1
    16'b11100101_10110010 : OUT <= 1;  //229 / 178 = 1
    16'b11100101_10110011 : OUT <= 1;  //229 / 179 = 1
    16'b11100101_10110100 : OUT <= 1;  //229 / 180 = 1
    16'b11100101_10110101 : OUT <= 1;  //229 / 181 = 1
    16'b11100101_10110110 : OUT <= 1;  //229 / 182 = 1
    16'b11100101_10110111 : OUT <= 1;  //229 / 183 = 1
    16'b11100101_10111000 : OUT <= 1;  //229 / 184 = 1
    16'b11100101_10111001 : OUT <= 1;  //229 / 185 = 1
    16'b11100101_10111010 : OUT <= 1;  //229 / 186 = 1
    16'b11100101_10111011 : OUT <= 1;  //229 / 187 = 1
    16'b11100101_10111100 : OUT <= 1;  //229 / 188 = 1
    16'b11100101_10111101 : OUT <= 1;  //229 / 189 = 1
    16'b11100101_10111110 : OUT <= 1;  //229 / 190 = 1
    16'b11100101_10111111 : OUT <= 1;  //229 / 191 = 1
    16'b11100101_11000000 : OUT <= 1;  //229 / 192 = 1
    16'b11100101_11000001 : OUT <= 1;  //229 / 193 = 1
    16'b11100101_11000010 : OUT <= 1;  //229 / 194 = 1
    16'b11100101_11000011 : OUT <= 1;  //229 / 195 = 1
    16'b11100101_11000100 : OUT <= 1;  //229 / 196 = 1
    16'b11100101_11000101 : OUT <= 1;  //229 / 197 = 1
    16'b11100101_11000110 : OUT <= 1;  //229 / 198 = 1
    16'b11100101_11000111 : OUT <= 1;  //229 / 199 = 1
    16'b11100101_11001000 : OUT <= 1;  //229 / 200 = 1
    16'b11100101_11001001 : OUT <= 1;  //229 / 201 = 1
    16'b11100101_11001010 : OUT <= 1;  //229 / 202 = 1
    16'b11100101_11001011 : OUT <= 1;  //229 / 203 = 1
    16'b11100101_11001100 : OUT <= 1;  //229 / 204 = 1
    16'b11100101_11001101 : OUT <= 1;  //229 / 205 = 1
    16'b11100101_11001110 : OUT <= 1;  //229 / 206 = 1
    16'b11100101_11001111 : OUT <= 1;  //229 / 207 = 1
    16'b11100101_11010000 : OUT <= 1;  //229 / 208 = 1
    16'b11100101_11010001 : OUT <= 1;  //229 / 209 = 1
    16'b11100101_11010010 : OUT <= 1;  //229 / 210 = 1
    16'b11100101_11010011 : OUT <= 1;  //229 / 211 = 1
    16'b11100101_11010100 : OUT <= 1;  //229 / 212 = 1
    16'b11100101_11010101 : OUT <= 1;  //229 / 213 = 1
    16'b11100101_11010110 : OUT <= 1;  //229 / 214 = 1
    16'b11100101_11010111 : OUT <= 1;  //229 / 215 = 1
    16'b11100101_11011000 : OUT <= 1;  //229 / 216 = 1
    16'b11100101_11011001 : OUT <= 1;  //229 / 217 = 1
    16'b11100101_11011010 : OUT <= 1;  //229 / 218 = 1
    16'b11100101_11011011 : OUT <= 1;  //229 / 219 = 1
    16'b11100101_11011100 : OUT <= 1;  //229 / 220 = 1
    16'b11100101_11011101 : OUT <= 1;  //229 / 221 = 1
    16'b11100101_11011110 : OUT <= 1;  //229 / 222 = 1
    16'b11100101_11011111 : OUT <= 1;  //229 / 223 = 1
    16'b11100101_11100000 : OUT <= 1;  //229 / 224 = 1
    16'b11100101_11100001 : OUT <= 1;  //229 / 225 = 1
    16'b11100101_11100010 : OUT <= 1;  //229 / 226 = 1
    16'b11100101_11100011 : OUT <= 1;  //229 / 227 = 1
    16'b11100101_11100100 : OUT <= 1;  //229 / 228 = 1
    16'b11100101_11100101 : OUT <= 1;  //229 / 229 = 1
    16'b11100101_11100110 : OUT <= 0;  //229 / 230 = 0
    16'b11100101_11100111 : OUT <= 0;  //229 / 231 = 0
    16'b11100101_11101000 : OUT <= 0;  //229 / 232 = 0
    16'b11100101_11101001 : OUT <= 0;  //229 / 233 = 0
    16'b11100101_11101010 : OUT <= 0;  //229 / 234 = 0
    16'b11100101_11101011 : OUT <= 0;  //229 / 235 = 0
    16'b11100101_11101100 : OUT <= 0;  //229 / 236 = 0
    16'b11100101_11101101 : OUT <= 0;  //229 / 237 = 0
    16'b11100101_11101110 : OUT <= 0;  //229 / 238 = 0
    16'b11100101_11101111 : OUT <= 0;  //229 / 239 = 0
    16'b11100101_11110000 : OUT <= 0;  //229 / 240 = 0
    16'b11100101_11110001 : OUT <= 0;  //229 / 241 = 0
    16'b11100101_11110010 : OUT <= 0;  //229 / 242 = 0
    16'b11100101_11110011 : OUT <= 0;  //229 / 243 = 0
    16'b11100101_11110100 : OUT <= 0;  //229 / 244 = 0
    16'b11100101_11110101 : OUT <= 0;  //229 / 245 = 0
    16'b11100101_11110110 : OUT <= 0;  //229 / 246 = 0
    16'b11100101_11110111 : OUT <= 0;  //229 / 247 = 0
    16'b11100101_11111000 : OUT <= 0;  //229 / 248 = 0
    16'b11100101_11111001 : OUT <= 0;  //229 / 249 = 0
    16'b11100101_11111010 : OUT <= 0;  //229 / 250 = 0
    16'b11100101_11111011 : OUT <= 0;  //229 / 251 = 0
    16'b11100101_11111100 : OUT <= 0;  //229 / 252 = 0
    16'b11100101_11111101 : OUT <= 0;  //229 / 253 = 0
    16'b11100101_11111110 : OUT <= 0;  //229 / 254 = 0
    16'b11100101_11111111 : OUT <= 0;  //229 / 255 = 0
    16'b11100110_00000000 : OUT <= 0;  //230 / 0 = 0
    16'b11100110_00000001 : OUT <= 230;  //230 / 1 = 230
    16'b11100110_00000010 : OUT <= 115;  //230 / 2 = 115
    16'b11100110_00000011 : OUT <= 76;  //230 / 3 = 76
    16'b11100110_00000100 : OUT <= 57;  //230 / 4 = 57
    16'b11100110_00000101 : OUT <= 46;  //230 / 5 = 46
    16'b11100110_00000110 : OUT <= 38;  //230 / 6 = 38
    16'b11100110_00000111 : OUT <= 32;  //230 / 7 = 32
    16'b11100110_00001000 : OUT <= 28;  //230 / 8 = 28
    16'b11100110_00001001 : OUT <= 25;  //230 / 9 = 25
    16'b11100110_00001010 : OUT <= 23;  //230 / 10 = 23
    16'b11100110_00001011 : OUT <= 20;  //230 / 11 = 20
    16'b11100110_00001100 : OUT <= 19;  //230 / 12 = 19
    16'b11100110_00001101 : OUT <= 17;  //230 / 13 = 17
    16'b11100110_00001110 : OUT <= 16;  //230 / 14 = 16
    16'b11100110_00001111 : OUT <= 15;  //230 / 15 = 15
    16'b11100110_00010000 : OUT <= 14;  //230 / 16 = 14
    16'b11100110_00010001 : OUT <= 13;  //230 / 17 = 13
    16'b11100110_00010010 : OUT <= 12;  //230 / 18 = 12
    16'b11100110_00010011 : OUT <= 12;  //230 / 19 = 12
    16'b11100110_00010100 : OUT <= 11;  //230 / 20 = 11
    16'b11100110_00010101 : OUT <= 10;  //230 / 21 = 10
    16'b11100110_00010110 : OUT <= 10;  //230 / 22 = 10
    16'b11100110_00010111 : OUT <= 10;  //230 / 23 = 10
    16'b11100110_00011000 : OUT <= 9;  //230 / 24 = 9
    16'b11100110_00011001 : OUT <= 9;  //230 / 25 = 9
    16'b11100110_00011010 : OUT <= 8;  //230 / 26 = 8
    16'b11100110_00011011 : OUT <= 8;  //230 / 27 = 8
    16'b11100110_00011100 : OUT <= 8;  //230 / 28 = 8
    16'b11100110_00011101 : OUT <= 7;  //230 / 29 = 7
    16'b11100110_00011110 : OUT <= 7;  //230 / 30 = 7
    16'b11100110_00011111 : OUT <= 7;  //230 / 31 = 7
    16'b11100110_00100000 : OUT <= 7;  //230 / 32 = 7
    16'b11100110_00100001 : OUT <= 6;  //230 / 33 = 6
    16'b11100110_00100010 : OUT <= 6;  //230 / 34 = 6
    16'b11100110_00100011 : OUT <= 6;  //230 / 35 = 6
    16'b11100110_00100100 : OUT <= 6;  //230 / 36 = 6
    16'b11100110_00100101 : OUT <= 6;  //230 / 37 = 6
    16'b11100110_00100110 : OUT <= 6;  //230 / 38 = 6
    16'b11100110_00100111 : OUT <= 5;  //230 / 39 = 5
    16'b11100110_00101000 : OUT <= 5;  //230 / 40 = 5
    16'b11100110_00101001 : OUT <= 5;  //230 / 41 = 5
    16'b11100110_00101010 : OUT <= 5;  //230 / 42 = 5
    16'b11100110_00101011 : OUT <= 5;  //230 / 43 = 5
    16'b11100110_00101100 : OUT <= 5;  //230 / 44 = 5
    16'b11100110_00101101 : OUT <= 5;  //230 / 45 = 5
    16'b11100110_00101110 : OUT <= 5;  //230 / 46 = 5
    16'b11100110_00101111 : OUT <= 4;  //230 / 47 = 4
    16'b11100110_00110000 : OUT <= 4;  //230 / 48 = 4
    16'b11100110_00110001 : OUT <= 4;  //230 / 49 = 4
    16'b11100110_00110010 : OUT <= 4;  //230 / 50 = 4
    16'b11100110_00110011 : OUT <= 4;  //230 / 51 = 4
    16'b11100110_00110100 : OUT <= 4;  //230 / 52 = 4
    16'b11100110_00110101 : OUT <= 4;  //230 / 53 = 4
    16'b11100110_00110110 : OUT <= 4;  //230 / 54 = 4
    16'b11100110_00110111 : OUT <= 4;  //230 / 55 = 4
    16'b11100110_00111000 : OUT <= 4;  //230 / 56 = 4
    16'b11100110_00111001 : OUT <= 4;  //230 / 57 = 4
    16'b11100110_00111010 : OUT <= 3;  //230 / 58 = 3
    16'b11100110_00111011 : OUT <= 3;  //230 / 59 = 3
    16'b11100110_00111100 : OUT <= 3;  //230 / 60 = 3
    16'b11100110_00111101 : OUT <= 3;  //230 / 61 = 3
    16'b11100110_00111110 : OUT <= 3;  //230 / 62 = 3
    16'b11100110_00111111 : OUT <= 3;  //230 / 63 = 3
    16'b11100110_01000000 : OUT <= 3;  //230 / 64 = 3
    16'b11100110_01000001 : OUT <= 3;  //230 / 65 = 3
    16'b11100110_01000010 : OUT <= 3;  //230 / 66 = 3
    16'b11100110_01000011 : OUT <= 3;  //230 / 67 = 3
    16'b11100110_01000100 : OUT <= 3;  //230 / 68 = 3
    16'b11100110_01000101 : OUT <= 3;  //230 / 69 = 3
    16'b11100110_01000110 : OUT <= 3;  //230 / 70 = 3
    16'b11100110_01000111 : OUT <= 3;  //230 / 71 = 3
    16'b11100110_01001000 : OUT <= 3;  //230 / 72 = 3
    16'b11100110_01001001 : OUT <= 3;  //230 / 73 = 3
    16'b11100110_01001010 : OUT <= 3;  //230 / 74 = 3
    16'b11100110_01001011 : OUT <= 3;  //230 / 75 = 3
    16'b11100110_01001100 : OUT <= 3;  //230 / 76 = 3
    16'b11100110_01001101 : OUT <= 2;  //230 / 77 = 2
    16'b11100110_01001110 : OUT <= 2;  //230 / 78 = 2
    16'b11100110_01001111 : OUT <= 2;  //230 / 79 = 2
    16'b11100110_01010000 : OUT <= 2;  //230 / 80 = 2
    16'b11100110_01010001 : OUT <= 2;  //230 / 81 = 2
    16'b11100110_01010010 : OUT <= 2;  //230 / 82 = 2
    16'b11100110_01010011 : OUT <= 2;  //230 / 83 = 2
    16'b11100110_01010100 : OUT <= 2;  //230 / 84 = 2
    16'b11100110_01010101 : OUT <= 2;  //230 / 85 = 2
    16'b11100110_01010110 : OUT <= 2;  //230 / 86 = 2
    16'b11100110_01010111 : OUT <= 2;  //230 / 87 = 2
    16'b11100110_01011000 : OUT <= 2;  //230 / 88 = 2
    16'b11100110_01011001 : OUT <= 2;  //230 / 89 = 2
    16'b11100110_01011010 : OUT <= 2;  //230 / 90 = 2
    16'b11100110_01011011 : OUT <= 2;  //230 / 91 = 2
    16'b11100110_01011100 : OUT <= 2;  //230 / 92 = 2
    16'b11100110_01011101 : OUT <= 2;  //230 / 93 = 2
    16'b11100110_01011110 : OUT <= 2;  //230 / 94 = 2
    16'b11100110_01011111 : OUT <= 2;  //230 / 95 = 2
    16'b11100110_01100000 : OUT <= 2;  //230 / 96 = 2
    16'b11100110_01100001 : OUT <= 2;  //230 / 97 = 2
    16'b11100110_01100010 : OUT <= 2;  //230 / 98 = 2
    16'b11100110_01100011 : OUT <= 2;  //230 / 99 = 2
    16'b11100110_01100100 : OUT <= 2;  //230 / 100 = 2
    16'b11100110_01100101 : OUT <= 2;  //230 / 101 = 2
    16'b11100110_01100110 : OUT <= 2;  //230 / 102 = 2
    16'b11100110_01100111 : OUT <= 2;  //230 / 103 = 2
    16'b11100110_01101000 : OUT <= 2;  //230 / 104 = 2
    16'b11100110_01101001 : OUT <= 2;  //230 / 105 = 2
    16'b11100110_01101010 : OUT <= 2;  //230 / 106 = 2
    16'b11100110_01101011 : OUT <= 2;  //230 / 107 = 2
    16'b11100110_01101100 : OUT <= 2;  //230 / 108 = 2
    16'b11100110_01101101 : OUT <= 2;  //230 / 109 = 2
    16'b11100110_01101110 : OUT <= 2;  //230 / 110 = 2
    16'b11100110_01101111 : OUT <= 2;  //230 / 111 = 2
    16'b11100110_01110000 : OUT <= 2;  //230 / 112 = 2
    16'b11100110_01110001 : OUT <= 2;  //230 / 113 = 2
    16'b11100110_01110010 : OUT <= 2;  //230 / 114 = 2
    16'b11100110_01110011 : OUT <= 2;  //230 / 115 = 2
    16'b11100110_01110100 : OUT <= 1;  //230 / 116 = 1
    16'b11100110_01110101 : OUT <= 1;  //230 / 117 = 1
    16'b11100110_01110110 : OUT <= 1;  //230 / 118 = 1
    16'b11100110_01110111 : OUT <= 1;  //230 / 119 = 1
    16'b11100110_01111000 : OUT <= 1;  //230 / 120 = 1
    16'b11100110_01111001 : OUT <= 1;  //230 / 121 = 1
    16'b11100110_01111010 : OUT <= 1;  //230 / 122 = 1
    16'b11100110_01111011 : OUT <= 1;  //230 / 123 = 1
    16'b11100110_01111100 : OUT <= 1;  //230 / 124 = 1
    16'b11100110_01111101 : OUT <= 1;  //230 / 125 = 1
    16'b11100110_01111110 : OUT <= 1;  //230 / 126 = 1
    16'b11100110_01111111 : OUT <= 1;  //230 / 127 = 1
    16'b11100110_10000000 : OUT <= 1;  //230 / 128 = 1
    16'b11100110_10000001 : OUT <= 1;  //230 / 129 = 1
    16'b11100110_10000010 : OUT <= 1;  //230 / 130 = 1
    16'b11100110_10000011 : OUT <= 1;  //230 / 131 = 1
    16'b11100110_10000100 : OUT <= 1;  //230 / 132 = 1
    16'b11100110_10000101 : OUT <= 1;  //230 / 133 = 1
    16'b11100110_10000110 : OUT <= 1;  //230 / 134 = 1
    16'b11100110_10000111 : OUT <= 1;  //230 / 135 = 1
    16'b11100110_10001000 : OUT <= 1;  //230 / 136 = 1
    16'b11100110_10001001 : OUT <= 1;  //230 / 137 = 1
    16'b11100110_10001010 : OUT <= 1;  //230 / 138 = 1
    16'b11100110_10001011 : OUT <= 1;  //230 / 139 = 1
    16'b11100110_10001100 : OUT <= 1;  //230 / 140 = 1
    16'b11100110_10001101 : OUT <= 1;  //230 / 141 = 1
    16'b11100110_10001110 : OUT <= 1;  //230 / 142 = 1
    16'b11100110_10001111 : OUT <= 1;  //230 / 143 = 1
    16'b11100110_10010000 : OUT <= 1;  //230 / 144 = 1
    16'b11100110_10010001 : OUT <= 1;  //230 / 145 = 1
    16'b11100110_10010010 : OUT <= 1;  //230 / 146 = 1
    16'b11100110_10010011 : OUT <= 1;  //230 / 147 = 1
    16'b11100110_10010100 : OUT <= 1;  //230 / 148 = 1
    16'b11100110_10010101 : OUT <= 1;  //230 / 149 = 1
    16'b11100110_10010110 : OUT <= 1;  //230 / 150 = 1
    16'b11100110_10010111 : OUT <= 1;  //230 / 151 = 1
    16'b11100110_10011000 : OUT <= 1;  //230 / 152 = 1
    16'b11100110_10011001 : OUT <= 1;  //230 / 153 = 1
    16'b11100110_10011010 : OUT <= 1;  //230 / 154 = 1
    16'b11100110_10011011 : OUT <= 1;  //230 / 155 = 1
    16'b11100110_10011100 : OUT <= 1;  //230 / 156 = 1
    16'b11100110_10011101 : OUT <= 1;  //230 / 157 = 1
    16'b11100110_10011110 : OUT <= 1;  //230 / 158 = 1
    16'b11100110_10011111 : OUT <= 1;  //230 / 159 = 1
    16'b11100110_10100000 : OUT <= 1;  //230 / 160 = 1
    16'b11100110_10100001 : OUT <= 1;  //230 / 161 = 1
    16'b11100110_10100010 : OUT <= 1;  //230 / 162 = 1
    16'b11100110_10100011 : OUT <= 1;  //230 / 163 = 1
    16'b11100110_10100100 : OUT <= 1;  //230 / 164 = 1
    16'b11100110_10100101 : OUT <= 1;  //230 / 165 = 1
    16'b11100110_10100110 : OUT <= 1;  //230 / 166 = 1
    16'b11100110_10100111 : OUT <= 1;  //230 / 167 = 1
    16'b11100110_10101000 : OUT <= 1;  //230 / 168 = 1
    16'b11100110_10101001 : OUT <= 1;  //230 / 169 = 1
    16'b11100110_10101010 : OUT <= 1;  //230 / 170 = 1
    16'b11100110_10101011 : OUT <= 1;  //230 / 171 = 1
    16'b11100110_10101100 : OUT <= 1;  //230 / 172 = 1
    16'b11100110_10101101 : OUT <= 1;  //230 / 173 = 1
    16'b11100110_10101110 : OUT <= 1;  //230 / 174 = 1
    16'b11100110_10101111 : OUT <= 1;  //230 / 175 = 1
    16'b11100110_10110000 : OUT <= 1;  //230 / 176 = 1
    16'b11100110_10110001 : OUT <= 1;  //230 / 177 = 1
    16'b11100110_10110010 : OUT <= 1;  //230 / 178 = 1
    16'b11100110_10110011 : OUT <= 1;  //230 / 179 = 1
    16'b11100110_10110100 : OUT <= 1;  //230 / 180 = 1
    16'b11100110_10110101 : OUT <= 1;  //230 / 181 = 1
    16'b11100110_10110110 : OUT <= 1;  //230 / 182 = 1
    16'b11100110_10110111 : OUT <= 1;  //230 / 183 = 1
    16'b11100110_10111000 : OUT <= 1;  //230 / 184 = 1
    16'b11100110_10111001 : OUT <= 1;  //230 / 185 = 1
    16'b11100110_10111010 : OUT <= 1;  //230 / 186 = 1
    16'b11100110_10111011 : OUT <= 1;  //230 / 187 = 1
    16'b11100110_10111100 : OUT <= 1;  //230 / 188 = 1
    16'b11100110_10111101 : OUT <= 1;  //230 / 189 = 1
    16'b11100110_10111110 : OUT <= 1;  //230 / 190 = 1
    16'b11100110_10111111 : OUT <= 1;  //230 / 191 = 1
    16'b11100110_11000000 : OUT <= 1;  //230 / 192 = 1
    16'b11100110_11000001 : OUT <= 1;  //230 / 193 = 1
    16'b11100110_11000010 : OUT <= 1;  //230 / 194 = 1
    16'b11100110_11000011 : OUT <= 1;  //230 / 195 = 1
    16'b11100110_11000100 : OUT <= 1;  //230 / 196 = 1
    16'b11100110_11000101 : OUT <= 1;  //230 / 197 = 1
    16'b11100110_11000110 : OUT <= 1;  //230 / 198 = 1
    16'b11100110_11000111 : OUT <= 1;  //230 / 199 = 1
    16'b11100110_11001000 : OUT <= 1;  //230 / 200 = 1
    16'b11100110_11001001 : OUT <= 1;  //230 / 201 = 1
    16'b11100110_11001010 : OUT <= 1;  //230 / 202 = 1
    16'b11100110_11001011 : OUT <= 1;  //230 / 203 = 1
    16'b11100110_11001100 : OUT <= 1;  //230 / 204 = 1
    16'b11100110_11001101 : OUT <= 1;  //230 / 205 = 1
    16'b11100110_11001110 : OUT <= 1;  //230 / 206 = 1
    16'b11100110_11001111 : OUT <= 1;  //230 / 207 = 1
    16'b11100110_11010000 : OUT <= 1;  //230 / 208 = 1
    16'b11100110_11010001 : OUT <= 1;  //230 / 209 = 1
    16'b11100110_11010010 : OUT <= 1;  //230 / 210 = 1
    16'b11100110_11010011 : OUT <= 1;  //230 / 211 = 1
    16'b11100110_11010100 : OUT <= 1;  //230 / 212 = 1
    16'b11100110_11010101 : OUT <= 1;  //230 / 213 = 1
    16'b11100110_11010110 : OUT <= 1;  //230 / 214 = 1
    16'b11100110_11010111 : OUT <= 1;  //230 / 215 = 1
    16'b11100110_11011000 : OUT <= 1;  //230 / 216 = 1
    16'b11100110_11011001 : OUT <= 1;  //230 / 217 = 1
    16'b11100110_11011010 : OUT <= 1;  //230 / 218 = 1
    16'b11100110_11011011 : OUT <= 1;  //230 / 219 = 1
    16'b11100110_11011100 : OUT <= 1;  //230 / 220 = 1
    16'b11100110_11011101 : OUT <= 1;  //230 / 221 = 1
    16'b11100110_11011110 : OUT <= 1;  //230 / 222 = 1
    16'b11100110_11011111 : OUT <= 1;  //230 / 223 = 1
    16'b11100110_11100000 : OUT <= 1;  //230 / 224 = 1
    16'b11100110_11100001 : OUT <= 1;  //230 / 225 = 1
    16'b11100110_11100010 : OUT <= 1;  //230 / 226 = 1
    16'b11100110_11100011 : OUT <= 1;  //230 / 227 = 1
    16'b11100110_11100100 : OUT <= 1;  //230 / 228 = 1
    16'b11100110_11100101 : OUT <= 1;  //230 / 229 = 1
    16'b11100110_11100110 : OUT <= 1;  //230 / 230 = 1
    16'b11100110_11100111 : OUT <= 0;  //230 / 231 = 0
    16'b11100110_11101000 : OUT <= 0;  //230 / 232 = 0
    16'b11100110_11101001 : OUT <= 0;  //230 / 233 = 0
    16'b11100110_11101010 : OUT <= 0;  //230 / 234 = 0
    16'b11100110_11101011 : OUT <= 0;  //230 / 235 = 0
    16'b11100110_11101100 : OUT <= 0;  //230 / 236 = 0
    16'b11100110_11101101 : OUT <= 0;  //230 / 237 = 0
    16'b11100110_11101110 : OUT <= 0;  //230 / 238 = 0
    16'b11100110_11101111 : OUT <= 0;  //230 / 239 = 0
    16'b11100110_11110000 : OUT <= 0;  //230 / 240 = 0
    16'b11100110_11110001 : OUT <= 0;  //230 / 241 = 0
    16'b11100110_11110010 : OUT <= 0;  //230 / 242 = 0
    16'b11100110_11110011 : OUT <= 0;  //230 / 243 = 0
    16'b11100110_11110100 : OUT <= 0;  //230 / 244 = 0
    16'b11100110_11110101 : OUT <= 0;  //230 / 245 = 0
    16'b11100110_11110110 : OUT <= 0;  //230 / 246 = 0
    16'b11100110_11110111 : OUT <= 0;  //230 / 247 = 0
    16'b11100110_11111000 : OUT <= 0;  //230 / 248 = 0
    16'b11100110_11111001 : OUT <= 0;  //230 / 249 = 0
    16'b11100110_11111010 : OUT <= 0;  //230 / 250 = 0
    16'b11100110_11111011 : OUT <= 0;  //230 / 251 = 0
    16'b11100110_11111100 : OUT <= 0;  //230 / 252 = 0
    16'b11100110_11111101 : OUT <= 0;  //230 / 253 = 0
    16'b11100110_11111110 : OUT <= 0;  //230 / 254 = 0
    16'b11100110_11111111 : OUT <= 0;  //230 / 255 = 0
    16'b11100111_00000000 : OUT <= 0;  //231 / 0 = 0
    16'b11100111_00000001 : OUT <= 231;  //231 / 1 = 231
    16'b11100111_00000010 : OUT <= 115;  //231 / 2 = 115
    16'b11100111_00000011 : OUT <= 77;  //231 / 3 = 77
    16'b11100111_00000100 : OUT <= 57;  //231 / 4 = 57
    16'b11100111_00000101 : OUT <= 46;  //231 / 5 = 46
    16'b11100111_00000110 : OUT <= 38;  //231 / 6 = 38
    16'b11100111_00000111 : OUT <= 33;  //231 / 7 = 33
    16'b11100111_00001000 : OUT <= 28;  //231 / 8 = 28
    16'b11100111_00001001 : OUT <= 25;  //231 / 9 = 25
    16'b11100111_00001010 : OUT <= 23;  //231 / 10 = 23
    16'b11100111_00001011 : OUT <= 21;  //231 / 11 = 21
    16'b11100111_00001100 : OUT <= 19;  //231 / 12 = 19
    16'b11100111_00001101 : OUT <= 17;  //231 / 13 = 17
    16'b11100111_00001110 : OUT <= 16;  //231 / 14 = 16
    16'b11100111_00001111 : OUT <= 15;  //231 / 15 = 15
    16'b11100111_00010000 : OUT <= 14;  //231 / 16 = 14
    16'b11100111_00010001 : OUT <= 13;  //231 / 17 = 13
    16'b11100111_00010010 : OUT <= 12;  //231 / 18 = 12
    16'b11100111_00010011 : OUT <= 12;  //231 / 19 = 12
    16'b11100111_00010100 : OUT <= 11;  //231 / 20 = 11
    16'b11100111_00010101 : OUT <= 11;  //231 / 21 = 11
    16'b11100111_00010110 : OUT <= 10;  //231 / 22 = 10
    16'b11100111_00010111 : OUT <= 10;  //231 / 23 = 10
    16'b11100111_00011000 : OUT <= 9;  //231 / 24 = 9
    16'b11100111_00011001 : OUT <= 9;  //231 / 25 = 9
    16'b11100111_00011010 : OUT <= 8;  //231 / 26 = 8
    16'b11100111_00011011 : OUT <= 8;  //231 / 27 = 8
    16'b11100111_00011100 : OUT <= 8;  //231 / 28 = 8
    16'b11100111_00011101 : OUT <= 7;  //231 / 29 = 7
    16'b11100111_00011110 : OUT <= 7;  //231 / 30 = 7
    16'b11100111_00011111 : OUT <= 7;  //231 / 31 = 7
    16'b11100111_00100000 : OUT <= 7;  //231 / 32 = 7
    16'b11100111_00100001 : OUT <= 7;  //231 / 33 = 7
    16'b11100111_00100010 : OUT <= 6;  //231 / 34 = 6
    16'b11100111_00100011 : OUT <= 6;  //231 / 35 = 6
    16'b11100111_00100100 : OUT <= 6;  //231 / 36 = 6
    16'b11100111_00100101 : OUT <= 6;  //231 / 37 = 6
    16'b11100111_00100110 : OUT <= 6;  //231 / 38 = 6
    16'b11100111_00100111 : OUT <= 5;  //231 / 39 = 5
    16'b11100111_00101000 : OUT <= 5;  //231 / 40 = 5
    16'b11100111_00101001 : OUT <= 5;  //231 / 41 = 5
    16'b11100111_00101010 : OUT <= 5;  //231 / 42 = 5
    16'b11100111_00101011 : OUT <= 5;  //231 / 43 = 5
    16'b11100111_00101100 : OUT <= 5;  //231 / 44 = 5
    16'b11100111_00101101 : OUT <= 5;  //231 / 45 = 5
    16'b11100111_00101110 : OUT <= 5;  //231 / 46 = 5
    16'b11100111_00101111 : OUT <= 4;  //231 / 47 = 4
    16'b11100111_00110000 : OUT <= 4;  //231 / 48 = 4
    16'b11100111_00110001 : OUT <= 4;  //231 / 49 = 4
    16'b11100111_00110010 : OUT <= 4;  //231 / 50 = 4
    16'b11100111_00110011 : OUT <= 4;  //231 / 51 = 4
    16'b11100111_00110100 : OUT <= 4;  //231 / 52 = 4
    16'b11100111_00110101 : OUT <= 4;  //231 / 53 = 4
    16'b11100111_00110110 : OUT <= 4;  //231 / 54 = 4
    16'b11100111_00110111 : OUT <= 4;  //231 / 55 = 4
    16'b11100111_00111000 : OUT <= 4;  //231 / 56 = 4
    16'b11100111_00111001 : OUT <= 4;  //231 / 57 = 4
    16'b11100111_00111010 : OUT <= 3;  //231 / 58 = 3
    16'b11100111_00111011 : OUT <= 3;  //231 / 59 = 3
    16'b11100111_00111100 : OUT <= 3;  //231 / 60 = 3
    16'b11100111_00111101 : OUT <= 3;  //231 / 61 = 3
    16'b11100111_00111110 : OUT <= 3;  //231 / 62 = 3
    16'b11100111_00111111 : OUT <= 3;  //231 / 63 = 3
    16'b11100111_01000000 : OUT <= 3;  //231 / 64 = 3
    16'b11100111_01000001 : OUT <= 3;  //231 / 65 = 3
    16'b11100111_01000010 : OUT <= 3;  //231 / 66 = 3
    16'b11100111_01000011 : OUT <= 3;  //231 / 67 = 3
    16'b11100111_01000100 : OUT <= 3;  //231 / 68 = 3
    16'b11100111_01000101 : OUT <= 3;  //231 / 69 = 3
    16'b11100111_01000110 : OUT <= 3;  //231 / 70 = 3
    16'b11100111_01000111 : OUT <= 3;  //231 / 71 = 3
    16'b11100111_01001000 : OUT <= 3;  //231 / 72 = 3
    16'b11100111_01001001 : OUT <= 3;  //231 / 73 = 3
    16'b11100111_01001010 : OUT <= 3;  //231 / 74 = 3
    16'b11100111_01001011 : OUT <= 3;  //231 / 75 = 3
    16'b11100111_01001100 : OUT <= 3;  //231 / 76 = 3
    16'b11100111_01001101 : OUT <= 3;  //231 / 77 = 3
    16'b11100111_01001110 : OUT <= 2;  //231 / 78 = 2
    16'b11100111_01001111 : OUT <= 2;  //231 / 79 = 2
    16'b11100111_01010000 : OUT <= 2;  //231 / 80 = 2
    16'b11100111_01010001 : OUT <= 2;  //231 / 81 = 2
    16'b11100111_01010010 : OUT <= 2;  //231 / 82 = 2
    16'b11100111_01010011 : OUT <= 2;  //231 / 83 = 2
    16'b11100111_01010100 : OUT <= 2;  //231 / 84 = 2
    16'b11100111_01010101 : OUT <= 2;  //231 / 85 = 2
    16'b11100111_01010110 : OUT <= 2;  //231 / 86 = 2
    16'b11100111_01010111 : OUT <= 2;  //231 / 87 = 2
    16'b11100111_01011000 : OUT <= 2;  //231 / 88 = 2
    16'b11100111_01011001 : OUT <= 2;  //231 / 89 = 2
    16'b11100111_01011010 : OUT <= 2;  //231 / 90 = 2
    16'b11100111_01011011 : OUT <= 2;  //231 / 91 = 2
    16'b11100111_01011100 : OUT <= 2;  //231 / 92 = 2
    16'b11100111_01011101 : OUT <= 2;  //231 / 93 = 2
    16'b11100111_01011110 : OUT <= 2;  //231 / 94 = 2
    16'b11100111_01011111 : OUT <= 2;  //231 / 95 = 2
    16'b11100111_01100000 : OUT <= 2;  //231 / 96 = 2
    16'b11100111_01100001 : OUT <= 2;  //231 / 97 = 2
    16'b11100111_01100010 : OUT <= 2;  //231 / 98 = 2
    16'b11100111_01100011 : OUT <= 2;  //231 / 99 = 2
    16'b11100111_01100100 : OUT <= 2;  //231 / 100 = 2
    16'b11100111_01100101 : OUT <= 2;  //231 / 101 = 2
    16'b11100111_01100110 : OUT <= 2;  //231 / 102 = 2
    16'b11100111_01100111 : OUT <= 2;  //231 / 103 = 2
    16'b11100111_01101000 : OUT <= 2;  //231 / 104 = 2
    16'b11100111_01101001 : OUT <= 2;  //231 / 105 = 2
    16'b11100111_01101010 : OUT <= 2;  //231 / 106 = 2
    16'b11100111_01101011 : OUT <= 2;  //231 / 107 = 2
    16'b11100111_01101100 : OUT <= 2;  //231 / 108 = 2
    16'b11100111_01101101 : OUT <= 2;  //231 / 109 = 2
    16'b11100111_01101110 : OUT <= 2;  //231 / 110 = 2
    16'b11100111_01101111 : OUT <= 2;  //231 / 111 = 2
    16'b11100111_01110000 : OUT <= 2;  //231 / 112 = 2
    16'b11100111_01110001 : OUT <= 2;  //231 / 113 = 2
    16'b11100111_01110010 : OUT <= 2;  //231 / 114 = 2
    16'b11100111_01110011 : OUT <= 2;  //231 / 115 = 2
    16'b11100111_01110100 : OUT <= 1;  //231 / 116 = 1
    16'b11100111_01110101 : OUT <= 1;  //231 / 117 = 1
    16'b11100111_01110110 : OUT <= 1;  //231 / 118 = 1
    16'b11100111_01110111 : OUT <= 1;  //231 / 119 = 1
    16'b11100111_01111000 : OUT <= 1;  //231 / 120 = 1
    16'b11100111_01111001 : OUT <= 1;  //231 / 121 = 1
    16'b11100111_01111010 : OUT <= 1;  //231 / 122 = 1
    16'b11100111_01111011 : OUT <= 1;  //231 / 123 = 1
    16'b11100111_01111100 : OUT <= 1;  //231 / 124 = 1
    16'b11100111_01111101 : OUT <= 1;  //231 / 125 = 1
    16'b11100111_01111110 : OUT <= 1;  //231 / 126 = 1
    16'b11100111_01111111 : OUT <= 1;  //231 / 127 = 1
    16'b11100111_10000000 : OUT <= 1;  //231 / 128 = 1
    16'b11100111_10000001 : OUT <= 1;  //231 / 129 = 1
    16'b11100111_10000010 : OUT <= 1;  //231 / 130 = 1
    16'b11100111_10000011 : OUT <= 1;  //231 / 131 = 1
    16'b11100111_10000100 : OUT <= 1;  //231 / 132 = 1
    16'b11100111_10000101 : OUT <= 1;  //231 / 133 = 1
    16'b11100111_10000110 : OUT <= 1;  //231 / 134 = 1
    16'b11100111_10000111 : OUT <= 1;  //231 / 135 = 1
    16'b11100111_10001000 : OUT <= 1;  //231 / 136 = 1
    16'b11100111_10001001 : OUT <= 1;  //231 / 137 = 1
    16'b11100111_10001010 : OUT <= 1;  //231 / 138 = 1
    16'b11100111_10001011 : OUT <= 1;  //231 / 139 = 1
    16'b11100111_10001100 : OUT <= 1;  //231 / 140 = 1
    16'b11100111_10001101 : OUT <= 1;  //231 / 141 = 1
    16'b11100111_10001110 : OUT <= 1;  //231 / 142 = 1
    16'b11100111_10001111 : OUT <= 1;  //231 / 143 = 1
    16'b11100111_10010000 : OUT <= 1;  //231 / 144 = 1
    16'b11100111_10010001 : OUT <= 1;  //231 / 145 = 1
    16'b11100111_10010010 : OUT <= 1;  //231 / 146 = 1
    16'b11100111_10010011 : OUT <= 1;  //231 / 147 = 1
    16'b11100111_10010100 : OUT <= 1;  //231 / 148 = 1
    16'b11100111_10010101 : OUT <= 1;  //231 / 149 = 1
    16'b11100111_10010110 : OUT <= 1;  //231 / 150 = 1
    16'b11100111_10010111 : OUT <= 1;  //231 / 151 = 1
    16'b11100111_10011000 : OUT <= 1;  //231 / 152 = 1
    16'b11100111_10011001 : OUT <= 1;  //231 / 153 = 1
    16'b11100111_10011010 : OUT <= 1;  //231 / 154 = 1
    16'b11100111_10011011 : OUT <= 1;  //231 / 155 = 1
    16'b11100111_10011100 : OUT <= 1;  //231 / 156 = 1
    16'b11100111_10011101 : OUT <= 1;  //231 / 157 = 1
    16'b11100111_10011110 : OUT <= 1;  //231 / 158 = 1
    16'b11100111_10011111 : OUT <= 1;  //231 / 159 = 1
    16'b11100111_10100000 : OUT <= 1;  //231 / 160 = 1
    16'b11100111_10100001 : OUT <= 1;  //231 / 161 = 1
    16'b11100111_10100010 : OUT <= 1;  //231 / 162 = 1
    16'b11100111_10100011 : OUT <= 1;  //231 / 163 = 1
    16'b11100111_10100100 : OUT <= 1;  //231 / 164 = 1
    16'b11100111_10100101 : OUT <= 1;  //231 / 165 = 1
    16'b11100111_10100110 : OUT <= 1;  //231 / 166 = 1
    16'b11100111_10100111 : OUT <= 1;  //231 / 167 = 1
    16'b11100111_10101000 : OUT <= 1;  //231 / 168 = 1
    16'b11100111_10101001 : OUT <= 1;  //231 / 169 = 1
    16'b11100111_10101010 : OUT <= 1;  //231 / 170 = 1
    16'b11100111_10101011 : OUT <= 1;  //231 / 171 = 1
    16'b11100111_10101100 : OUT <= 1;  //231 / 172 = 1
    16'b11100111_10101101 : OUT <= 1;  //231 / 173 = 1
    16'b11100111_10101110 : OUT <= 1;  //231 / 174 = 1
    16'b11100111_10101111 : OUT <= 1;  //231 / 175 = 1
    16'b11100111_10110000 : OUT <= 1;  //231 / 176 = 1
    16'b11100111_10110001 : OUT <= 1;  //231 / 177 = 1
    16'b11100111_10110010 : OUT <= 1;  //231 / 178 = 1
    16'b11100111_10110011 : OUT <= 1;  //231 / 179 = 1
    16'b11100111_10110100 : OUT <= 1;  //231 / 180 = 1
    16'b11100111_10110101 : OUT <= 1;  //231 / 181 = 1
    16'b11100111_10110110 : OUT <= 1;  //231 / 182 = 1
    16'b11100111_10110111 : OUT <= 1;  //231 / 183 = 1
    16'b11100111_10111000 : OUT <= 1;  //231 / 184 = 1
    16'b11100111_10111001 : OUT <= 1;  //231 / 185 = 1
    16'b11100111_10111010 : OUT <= 1;  //231 / 186 = 1
    16'b11100111_10111011 : OUT <= 1;  //231 / 187 = 1
    16'b11100111_10111100 : OUT <= 1;  //231 / 188 = 1
    16'b11100111_10111101 : OUT <= 1;  //231 / 189 = 1
    16'b11100111_10111110 : OUT <= 1;  //231 / 190 = 1
    16'b11100111_10111111 : OUT <= 1;  //231 / 191 = 1
    16'b11100111_11000000 : OUT <= 1;  //231 / 192 = 1
    16'b11100111_11000001 : OUT <= 1;  //231 / 193 = 1
    16'b11100111_11000010 : OUT <= 1;  //231 / 194 = 1
    16'b11100111_11000011 : OUT <= 1;  //231 / 195 = 1
    16'b11100111_11000100 : OUT <= 1;  //231 / 196 = 1
    16'b11100111_11000101 : OUT <= 1;  //231 / 197 = 1
    16'b11100111_11000110 : OUT <= 1;  //231 / 198 = 1
    16'b11100111_11000111 : OUT <= 1;  //231 / 199 = 1
    16'b11100111_11001000 : OUT <= 1;  //231 / 200 = 1
    16'b11100111_11001001 : OUT <= 1;  //231 / 201 = 1
    16'b11100111_11001010 : OUT <= 1;  //231 / 202 = 1
    16'b11100111_11001011 : OUT <= 1;  //231 / 203 = 1
    16'b11100111_11001100 : OUT <= 1;  //231 / 204 = 1
    16'b11100111_11001101 : OUT <= 1;  //231 / 205 = 1
    16'b11100111_11001110 : OUT <= 1;  //231 / 206 = 1
    16'b11100111_11001111 : OUT <= 1;  //231 / 207 = 1
    16'b11100111_11010000 : OUT <= 1;  //231 / 208 = 1
    16'b11100111_11010001 : OUT <= 1;  //231 / 209 = 1
    16'b11100111_11010010 : OUT <= 1;  //231 / 210 = 1
    16'b11100111_11010011 : OUT <= 1;  //231 / 211 = 1
    16'b11100111_11010100 : OUT <= 1;  //231 / 212 = 1
    16'b11100111_11010101 : OUT <= 1;  //231 / 213 = 1
    16'b11100111_11010110 : OUT <= 1;  //231 / 214 = 1
    16'b11100111_11010111 : OUT <= 1;  //231 / 215 = 1
    16'b11100111_11011000 : OUT <= 1;  //231 / 216 = 1
    16'b11100111_11011001 : OUT <= 1;  //231 / 217 = 1
    16'b11100111_11011010 : OUT <= 1;  //231 / 218 = 1
    16'b11100111_11011011 : OUT <= 1;  //231 / 219 = 1
    16'b11100111_11011100 : OUT <= 1;  //231 / 220 = 1
    16'b11100111_11011101 : OUT <= 1;  //231 / 221 = 1
    16'b11100111_11011110 : OUT <= 1;  //231 / 222 = 1
    16'b11100111_11011111 : OUT <= 1;  //231 / 223 = 1
    16'b11100111_11100000 : OUT <= 1;  //231 / 224 = 1
    16'b11100111_11100001 : OUT <= 1;  //231 / 225 = 1
    16'b11100111_11100010 : OUT <= 1;  //231 / 226 = 1
    16'b11100111_11100011 : OUT <= 1;  //231 / 227 = 1
    16'b11100111_11100100 : OUT <= 1;  //231 / 228 = 1
    16'b11100111_11100101 : OUT <= 1;  //231 / 229 = 1
    16'b11100111_11100110 : OUT <= 1;  //231 / 230 = 1
    16'b11100111_11100111 : OUT <= 1;  //231 / 231 = 1
    16'b11100111_11101000 : OUT <= 0;  //231 / 232 = 0
    16'b11100111_11101001 : OUT <= 0;  //231 / 233 = 0
    16'b11100111_11101010 : OUT <= 0;  //231 / 234 = 0
    16'b11100111_11101011 : OUT <= 0;  //231 / 235 = 0
    16'b11100111_11101100 : OUT <= 0;  //231 / 236 = 0
    16'b11100111_11101101 : OUT <= 0;  //231 / 237 = 0
    16'b11100111_11101110 : OUT <= 0;  //231 / 238 = 0
    16'b11100111_11101111 : OUT <= 0;  //231 / 239 = 0
    16'b11100111_11110000 : OUT <= 0;  //231 / 240 = 0
    16'b11100111_11110001 : OUT <= 0;  //231 / 241 = 0
    16'b11100111_11110010 : OUT <= 0;  //231 / 242 = 0
    16'b11100111_11110011 : OUT <= 0;  //231 / 243 = 0
    16'b11100111_11110100 : OUT <= 0;  //231 / 244 = 0
    16'b11100111_11110101 : OUT <= 0;  //231 / 245 = 0
    16'b11100111_11110110 : OUT <= 0;  //231 / 246 = 0
    16'b11100111_11110111 : OUT <= 0;  //231 / 247 = 0
    16'b11100111_11111000 : OUT <= 0;  //231 / 248 = 0
    16'b11100111_11111001 : OUT <= 0;  //231 / 249 = 0
    16'b11100111_11111010 : OUT <= 0;  //231 / 250 = 0
    16'b11100111_11111011 : OUT <= 0;  //231 / 251 = 0
    16'b11100111_11111100 : OUT <= 0;  //231 / 252 = 0
    16'b11100111_11111101 : OUT <= 0;  //231 / 253 = 0
    16'b11100111_11111110 : OUT <= 0;  //231 / 254 = 0
    16'b11100111_11111111 : OUT <= 0;  //231 / 255 = 0
    16'b11101000_00000000 : OUT <= 0;  //232 / 0 = 0
    16'b11101000_00000001 : OUT <= 232;  //232 / 1 = 232
    16'b11101000_00000010 : OUT <= 116;  //232 / 2 = 116
    16'b11101000_00000011 : OUT <= 77;  //232 / 3 = 77
    16'b11101000_00000100 : OUT <= 58;  //232 / 4 = 58
    16'b11101000_00000101 : OUT <= 46;  //232 / 5 = 46
    16'b11101000_00000110 : OUT <= 38;  //232 / 6 = 38
    16'b11101000_00000111 : OUT <= 33;  //232 / 7 = 33
    16'b11101000_00001000 : OUT <= 29;  //232 / 8 = 29
    16'b11101000_00001001 : OUT <= 25;  //232 / 9 = 25
    16'b11101000_00001010 : OUT <= 23;  //232 / 10 = 23
    16'b11101000_00001011 : OUT <= 21;  //232 / 11 = 21
    16'b11101000_00001100 : OUT <= 19;  //232 / 12 = 19
    16'b11101000_00001101 : OUT <= 17;  //232 / 13 = 17
    16'b11101000_00001110 : OUT <= 16;  //232 / 14 = 16
    16'b11101000_00001111 : OUT <= 15;  //232 / 15 = 15
    16'b11101000_00010000 : OUT <= 14;  //232 / 16 = 14
    16'b11101000_00010001 : OUT <= 13;  //232 / 17 = 13
    16'b11101000_00010010 : OUT <= 12;  //232 / 18 = 12
    16'b11101000_00010011 : OUT <= 12;  //232 / 19 = 12
    16'b11101000_00010100 : OUT <= 11;  //232 / 20 = 11
    16'b11101000_00010101 : OUT <= 11;  //232 / 21 = 11
    16'b11101000_00010110 : OUT <= 10;  //232 / 22 = 10
    16'b11101000_00010111 : OUT <= 10;  //232 / 23 = 10
    16'b11101000_00011000 : OUT <= 9;  //232 / 24 = 9
    16'b11101000_00011001 : OUT <= 9;  //232 / 25 = 9
    16'b11101000_00011010 : OUT <= 8;  //232 / 26 = 8
    16'b11101000_00011011 : OUT <= 8;  //232 / 27 = 8
    16'b11101000_00011100 : OUT <= 8;  //232 / 28 = 8
    16'b11101000_00011101 : OUT <= 8;  //232 / 29 = 8
    16'b11101000_00011110 : OUT <= 7;  //232 / 30 = 7
    16'b11101000_00011111 : OUT <= 7;  //232 / 31 = 7
    16'b11101000_00100000 : OUT <= 7;  //232 / 32 = 7
    16'b11101000_00100001 : OUT <= 7;  //232 / 33 = 7
    16'b11101000_00100010 : OUT <= 6;  //232 / 34 = 6
    16'b11101000_00100011 : OUT <= 6;  //232 / 35 = 6
    16'b11101000_00100100 : OUT <= 6;  //232 / 36 = 6
    16'b11101000_00100101 : OUT <= 6;  //232 / 37 = 6
    16'b11101000_00100110 : OUT <= 6;  //232 / 38 = 6
    16'b11101000_00100111 : OUT <= 5;  //232 / 39 = 5
    16'b11101000_00101000 : OUT <= 5;  //232 / 40 = 5
    16'b11101000_00101001 : OUT <= 5;  //232 / 41 = 5
    16'b11101000_00101010 : OUT <= 5;  //232 / 42 = 5
    16'b11101000_00101011 : OUT <= 5;  //232 / 43 = 5
    16'b11101000_00101100 : OUT <= 5;  //232 / 44 = 5
    16'b11101000_00101101 : OUT <= 5;  //232 / 45 = 5
    16'b11101000_00101110 : OUT <= 5;  //232 / 46 = 5
    16'b11101000_00101111 : OUT <= 4;  //232 / 47 = 4
    16'b11101000_00110000 : OUT <= 4;  //232 / 48 = 4
    16'b11101000_00110001 : OUT <= 4;  //232 / 49 = 4
    16'b11101000_00110010 : OUT <= 4;  //232 / 50 = 4
    16'b11101000_00110011 : OUT <= 4;  //232 / 51 = 4
    16'b11101000_00110100 : OUT <= 4;  //232 / 52 = 4
    16'b11101000_00110101 : OUT <= 4;  //232 / 53 = 4
    16'b11101000_00110110 : OUT <= 4;  //232 / 54 = 4
    16'b11101000_00110111 : OUT <= 4;  //232 / 55 = 4
    16'b11101000_00111000 : OUT <= 4;  //232 / 56 = 4
    16'b11101000_00111001 : OUT <= 4;  //232 / 57 = 4
    16'b11101000_00111010 : OUT <= 4;  //232 / 58 = 4
    16'b11101000_00111011 : OUT <= 3;  //232 / 59 = 3
    16'b11101000_00111100 : OUT <= 3;  //232 / 60 = 3
    16'b11101000_00111101 : OUT <= 3;  //232 / 61 = 3
    16'b11101000_00111110 : OUT <= 3;  //232 / 62 = 3
    16'b11101000_00111111 : OUT <= 3;  //232 / 63 = 3
    16'b11101000_01000000 : OUT <= 3;  //232 / 64 = 3
    16'b11101000_01000001 : OUT <= 3;  //232 / 65 = 3
    16'b11101000_01000010 : OUT <= 3;  //232 / 66 = 3
    16'b11101000_01000011 : OUT <= 3;  //232 / 67 = 3
    16'b11101000_01000100 : OUT <= 3;  //232 / 68 = 3
    16'b11101000_01000101 : OUT <= 3;  //232 / 69 = 3
    16'b11101000_01000110 : OUT <= 3;  //232 / 70 = 3
    16'b11101000_01000111 : OUT <= 3;  //232 / 71 = 3
    16'b11101000_01001000 : OUT <= 3;  //232 / 72 = 3
    16'b11101000_01001001 : OUT <= 3;  //232 / 73 = 3
    16'b11101000_01001010 : OUT <= 3;  //232 / 74 = 3
    16'b11101000_01001011 : OUT <= 3;  //232 / 75 = 3
    16'b11101000_01001100 : OUT <= 3;  //232 / 76 = 3
    16'b11101000_01001101 : OUT <= 3;  //232 / 77 = 3
    16'b11101000_01001110 : OUT <= 2;  //232 / 78 = 2
    16'b11101000_01001111 : OUT <= 2;  //232 / 79 = 2
    16'b11101000_01010000 : OUT <= 2;  //232 / 80 = 2
    16'b11101000_01010001 : OUT <= 2;  //232 / 81 = 2
    16'b11101000_01010010 : OUT <= 2;  //232 / 82 = 2
    16'b11101000_01010011 : OUT <= 2;  //232 / 83 = 2
    16'b11101000_01010100 : OUT <= 2;  //232 / 84 = 2
    16'b11101000_01010101 : OUT <= 2;  //232 / 85 = 2
    16'b11101000_01010110 : OUT <= 2;  //232 / 86 = 2
    16'b11101000_01010111 : OUT <= 2;  //232 / 87 = 2
    16'b11101000_01011000 : OUT <= 2;  //232 / 88 = 2
    16'b11101000_01011001 : OUT <= 2;  //232 / 89 = 2
    16'b11101000_01011010 : OUT <= 2;  //232 / 90 = 2
    16'b11101000_01011011 : OUT <= 2;  //232 / 91 = 2
    16'b11101000_01011100 : OUT <= 2;  //232 / 92 = 2
    16'b11101000_01011101 : OUT <= 2;  //232 / 93 = 2
    16'b11101000_01011110 : OUT <= 2;  //232 / 94 = 2
    16'b11101000_01011111 : OUT <= 2;  //232 / 95 = 2
    16'b11101000_01100000 : OUT <= 2;  //232 / 96 = 2
    16'b11101000_01100001 : OUT <= 2;  //232 / 97 = 2
    16'b11101000_01100010 : OUT <= 2;  //232 / 98 = 2
    16'b11101000_01100011 : OUT <= 2;  //232 / 99 = 2
    16'b11101000_01100100 : OUT <= 2;  //232 / 100 = 2
    16'b11101000_01100101 : OUT <= 2;  //232 / 101 = 2
    16'b11101000_01100110 : OUT <= 2;  //232 / 102 = 2
    16'b11101000_01100111 : OUT <= 2;  //232 / 103 = 2
    16'b11101000_01101000 : OUT <= 2;  //232 / 104 = 2
    16'b11101000_01101001 : OUT <= 2;  //232 / 105 = 2
    16'b11101000_01101010 : OUT <= 2;  //232 / 106 = 2
    16'b11101000_01101011 : OUT <= 2;  //232 / 107 = 2
    16'b11101000_01101100 : OUT <= 2;  //232 / 108 = 2
    16'b11101000_01101101 : OUT <= 2;  //232 / 109 = 2
    16'b11101000_01101110 : OUT <= 2;  //232 / 110 = 2
    16'b11101000_01101111 : OUT <= 2;  //232 / 111 = 2
    16'b11101000_01110000 : OUT <= 2;  //232 / 112 = 2
    16'b11101000_01110001 : OUT <= 2;  //232 / 113 = 2
    16'b11101000_01110010 : OUT <= 2;  //232 / 114 = 2
    16'b11101000_01110011 : OUT <= 2;  //232 / 115 = 2
    16'b11101000_01110100 : OUT <= 2;  //232 / 116 = 2
    16'b11101000_01110101 : OUT <= 1;  //232 / 117 = 1
    16'b11101000_01110110 : OUT <= 1;  //232 / 118 = 1
    16'b11101000_01110111 : OUT <= 1;  //232 / 119 = 1
    16'b11101000_01111000 : OUT <= 1;  //232 / 120 = 1
    16'b11101000_01111001 : OUT <= 1;  //232 / 121 = 1
    16'b11101000_01111010 : OUT <= 1;  //232 / 122 = 1
    16'b11101000_01111011 : OUT <= 1;  //232 / 123 = 1
    16'b11101000_01111100 : OUT <= 1;  //232 / 124 = 1
    16'b11101000_01111101 : OUT <= 1;  //232 / 125 = 1
    16'b11101000_01111110 : OUT <= 1;  //232 / 126 = 1
    16'b11101000_01111111 : OUT <= 1;  //232 / 127 = 1
    16'b11101000_10000000 : OUT <= 1;  //232 / 128 = 1
    16'b11101000_10000001 : OUT <= 1;  //232 / 129 = 1
    16'b11101000_10000010 : OUT <= 1;  //232 / 130 = 1
    16'b11101000_10000011 : OUT <= 1;  //232 / 131 = 1
    16'b11101000_10000100 : OUT <= 1;  //232 / 132 = 1
    16'b11101000_10000101 : OUT <= 1;  //232 / 133 = 1
    16'b11101000_10000110 : OUT <= 1;  //232 / 134 = 1
    16'b11101000_10000111 : OUT <= 1;  //232 / 135 = 1
    16'b11101000_10001000 : OUT <= 1;  //232 / 136 = 1
    16'b11101000_10001001 : OUT <= 1;  //232 / 137 = 1
    16'b11101000_10001010 : OUT <= 1;  //232 / 138 = 1
    16'b11101000_10001011 : OUT <= 1;  //232 / 139 = 1
    16'b11101000_10001100 : OUT <= 1;  //232 / 140 = 1
    16'b11101000_10001101 : OUT <= 1;  //232 / 141 = 1
    16'b11101000_10001110 : OUT <= 1;  //232 / 142 = 1
    16'b11101000_10001111 : OUT <= 1;  //232 / 143 = 1
    16'b11101000_10010000 : OUT <= 1;  //232 / 144 = 1
    16'b11101000_10010001 : OUT <= 1;  //232 / 145 = 1
    16'b11101000_10010010 : OUT <= 1;  //232 / 146 = 1
    16'b11101000_10010011 : OUT <= 1;  //232 / 147 = 1
    16'b11101000_10010100 : OUT <= 1;  //232 / 148 = 1
    16'b11101000_10010101 : OUT <= 1;  //232 / 149 = 1
    16'b11101000_10010110 : OUT <= 1;  //232 / 150 = 1
    16'b11101000_10010111 : OUT <= 1;  //232 / 151 = 1
    16'b11101000_10011000 : OUT <= 1;  //232 / 152 = 1
    16'b11101000_10011001 : OUT <= 1;  //232 / 153 = 1
    16'b11101000_10011010 : OUT <= 1;  //232 / 154 = 1
    16'b11101000_10011011 : OUT <= 1;  //232 / 155 = 1
    16'b11101000_10011100 : OUT <= 1;  //232 / 156 = 1
    16'b11101000_10011101 : OUT <= 1;  //232 / 157 = 1
    16'b11101000_10011110 : OUT <= 1;  //232 / 158 = 1
    16'b11101000_10011111 : OUT <= 1;  //232 / 159 = 1
    16'b11101000_10100000 : OUT <= 1;  //232 / 160 = 1
    16'b11101000_10100001 : OUT <= 1;  //232 / 161 = 1
    16'b11101000_10100010 : OUT <= 1;  //232 / 162 = 1
    16'b11101000_10100011 : OUT <= 1;  //232 / 163 = 1
    16'b11101000_10100100 : OUT <= 1;  //232 / 164 = 1
    16'b11101000_10100101 : OUT <= 1;  //232 / 165 = 1
    16'b11101000_10100110 : OUT <= 1;  //232 / 166 = 1
    16'b11101000_10100111 : OUT <= 1;  //232 / 167 = 1
    16'b11101000_10101000 : OUT <= 1;  //232 / 168 = 1
    16'b11101000_10101001 : OUT <= 1;  //232 / 169 = 1
    16'b11101000_10101010 : OUT <= 1;  //232 / 170 = 1
    16'b11101000_10101011 : OUT <= 1;  //232 / 171 = 1
    16'b11101000_10101100 : OUT <= 1;  //232 / 172 = 1
    16'b11101000_10101101 : OUT <= 1;  //232 / 173 = 1
    16'b11101000_10101110 : OUT <= 1;  //232 / 174 = 1
    16'b11101000_10101111 : OUT <= 1;  //232 / 175 = 1
    16'b11101000_10110000 : OUT <= 1;  //232 / 176 = 1
    16'b11101000_10110001 : OUT <= 1;  //232 / 177 = 1
    16'b11101000_10110010 : OUT <= 1;  //232 / 178 = 1
    16'b11101000_10110011 : OUT <= 1;  //232 / 179 = 1
    16'b11101000_10110100 : OUT <= 1;  //232 / 180 = 1
    16'b11101000_10110101 : OUT <= 1;  //232 / 181 = 1
    16'b11101000_10110110 : OUT <= 1;  //232 / 182 = 1
    16'b11101000_10110111 : OUT <= 1;  //232 / 183 = 1
    16'b11101000_10111000 : OUT <= 1;  //232 / 184 = 1
    16'b11101000_10111001 : OUT <= 1;  //232 / 185 = 1
    16'b11101000_10111010 : OUT <= 1;  //232 / 186 = 1
    16'b11101000_10111011 : OUT <= 1;  //232 / 187 = 1
    16'b11101000_10111100 : OUT <= 1;  //232 / 188 = 1
    16'b11101000_10111101 : OUT <= 1;  //232 / 189 = 1
    16'b11101000_10111110 : OUT <= 1;  //232 / 190 = 1
    16'b11101000_10111111 : OUT <= 1;  //232 / 191 = 1
    16'b11101000_11000000 : OUT <= 1;  //232 / 192 = 1
    16'b11101000_11000001 : OUT <= 1;  //232 / 193 = 1
    16'b11101000_11000010 : OUT <= 1;  //232 / 194 = 1
    16'b11101000_11000011 : OUT <= 1;  //232 / 195 = 1
    16'b11101000_11000100 : OUT <= 1;  //232 / 196 = 1
    16'b11101000_11000101 : OUT <= 1;  //232 / 197 = 1
    16'b11101000_11000110 : OUT <= 1;  //232 / 198 = 1
    16'b11101000_11000111 : OUT <= 1;  //232 / 199 = 1
    16'b11101000_11001000 : OUT <= 1;  //232 / 200 = 1
    16'b11101000_11001001 : OUT <= 1;  //232 / 201 = 1
    16'b11101000_11001010 : OUT <= 1;  //232 / 202 = 1
    16'b11101000_11001011 : OUT <= 1;  //232 / 203 = 1
    16'b11101000_11001100 : OUT <= 1;  //232 / 204 = 1
    16'b11101000_11001101 : OUT <= 1;  //232 / 205 = 1
    16'b11101000_11001110 : OUT <= 1;  //232 / 206 = 1
    16'b11101000_11001111 : OUT <= 1;  //232 / 207 = 1
    16'b11101000_11010000 : OUT <= 1;  //232 / 208 = 1
    16'b11101000_11010001 : OUT <= 1;  //232 / 209 = 1
    16'b11101000_11010010 : OUT <= 1;  //232 / 210 = 1
    16'b11101000_11010011 : OUT <= 1;  //232 / 211 = 1
    16'b11101000_11010100 : OUT <= 1;  //232 / 212 = 1
    16'b11101000_11010101 : OUT <= 1;  //232 / 213 = 1
    16'b11101000_11010110 : OUT <= 1;  //232 / 214 = 1
    16'b11101000_11010111 : OUT <= 1;  //232 / 215 = 1
    16'b11101000_11011000 : OUT <= 1;  //232 / 216 = 1
    16'b11101000_11011001 : OUT <= 1;  //232 / 217 = 1
    16'b11101000_11011010 : OUT <= 1;  //232 / 218 = 1
    16'b11101000_11011011 : OUT <= 1;  //232 / 219 = 1
    16'b11101000_11011100 : OUT <= 1;  //232 / 220 = 1
    16'b11101000_11011101 : OUT <= 1;  //232 / 221 = 1
    16'b11101000_11011110 : OUT <= 1;  //232 / 222 = 1
    16'b11101000_11011111 : OUT <= 1;  //232 / 223 = 1
    16'b11101000_11100000 : OUT <= 1;  //232 / 224 = 1
    16'b11101000_11100001 : OUT <= 1;  //232 / 225 = 1
    16'b11101000_11100010 : OUT <= 1;  //232 / 226 = 1
    16'b11101000_11100011 : OUT <= 1;  //232 / 227 = 1
    16'b11101000_11100100 : OUT <= 1;  //232 / 228 = 1
    16'b11101000_11100101 : OUT <= 1;  //232 / 229 = 1
    16'b11101000_11100110 : OUT <= 1;  //232 / 230 = 1
    16'b11101000_11100111 : OUT <= 1;  //232 / 231 = 1
    16'b11101000_11101000 : OUT <= 1;  //232 / 232 = 1
    16'b11101000_11101001 : OUT <= 0;  //232 / 233 = 0
    16'b11101000_11101010 : OUT <= 0;  //232 / 234 = 0
    16'b11101000_11101011 : OUT <= 0;  //232 / 235 = 0
    16'b11101000_11101100 : OUT <= 0;  //232 / 236 = 0
    16'b11101000_11101101 : OUT <= 0;  //232 / 237 = 0
    16'b11101000_11101110 : OUT <= 0;  //232 / 238 = 0
    16'b11101000_11101111 : OUT <= 0;  //232 / 239 = 0
    16'b11101000_11110000 : OUT <= 0;  //232 / 240 = 0
    16'b11101000_11110001 : OUT <= 0;  //232 / 241 = 0
    16'b11101000_11110010 : OUT <= 0;  //232 / 242 = 0
    16'b11101000_11110011 : OUT <= 0;  //232 / 243 = 0
    16'b11101000_11110100 : OUT <= 0;  //232 / 244 = 0
    16'b11101000_11110101 : OUT <= 0;  //232 / 245 = 0
    16'b11101000_11110110 : OUT <= 0;  //232 / 246 = 0
    16'b11101000_11110111 : OUT <= 0;  //232 / 247 = 0
    16'b11101000_11111000 : OUT <= 0;  //232 / 248 = 0
    16'b11101000_11111001 : OUT <= 0;  //232 / 249 = 0
    16'b11101000_11111010 : OUT <= 0;  //232 / 250 = 0
    16'b11101000_11111011 : OUT <= 0;  //232 / 251 = 0
    16'b11101000_11111100 : OUT <= 0;  //232 / 252 = 0
    16'b11101000_11111101 : OUT <= 0;  //232 / 253 = 0
    16'b11101000_11111110 : OUT <= 0;  //232 / 254 = 0
    16'b11101000_11111111 : OUT <= 0;  //232 / 255 = 0
    16'b11101001_00000000 : OUT <= 0;  //233 / 0 = 0
    16'b11101001_00000001 : OUT <= 233;  //233 / 1 = 233
    16'b11101001_00000010 : OUT <= 116;  //233 / 2 = 116
    16'b11101001_00000011 : OUT <= 77;  //233 / 3 = 77
    16'b11101001_00000100 : OUT <= 58;  //233 / 4 = 58
    16'b11101001_00000101 : OUT <= 46;  //233 / 5 = 46
    16'b11101001_00000110 : OUT <= 38;  //233 / 6 = 38
    16'b11101001_00000111 : OUT <= 33;  //233 / 7 = 33
    16'b11101001_00001000 : OUT <= 29;  //233 / 8 = 29
    16'b11101001_00001001 : OUT <= 25;  //233 / 9 = 25
    16'b11101001_00001010 : OUT <= 23;  //233 / 10 = 23
    16'b11101001_00001011 : OUT <= 21;  //233 / 11 = 21
    16'b11101001_00001100 : OUT <= 19;  //233 / 12 = 19
    16'b11101001_00001101 : OUT <= 17;  //233 / 13 = 17
    16'b11101001_00001110 : OUT <= 16;  //233 / 14 = 16
    16'b11101001_00001111 : OUT <= 15;  //233 / 15 = 15
    16'b11101001_00010000 : OUT <= 14;  //233 / 16 = 14
    16'b11101001_00010001 : OUT <= 13;  //233 / 17 = 13
    16'b11101001_00010010 : OUT <= 12;  //233 / 18 = 12
    16'b11101001_00010011 : OUT <= 12;  //233 / 19 = 12
    16'b11101001_00010100 : OUT <= 11;  //233 / 20 = 11
    16'b11101001_00010101 : OUT <= 11;  //233 / 21 = 11
    16'b11101001_00010110 : OUT <= 10;  //233 / 22 = 10
    16'b11101001_00010111 : OUT <= 10;  //233 / 23 = 10
    16'b11101001_00011000 : OUT <= 9;  //233 / 24 = 9
    16'b11101001_00011001 : OUT <= 9;  //233 / 25 = 9
    16'b11101001_00011010 : OUT <= 8;  //233 / 26 = 8
    16'b11101001_00011011 : OUT <= 8;  //233 / 27 = 8
    16'b11101001_00011100 : OUT <= 8;  //233 / 28 = 8
    16'b11101001_00011101 : OUT <= 8;  //233 / 29 = 8
    16'b11101001_00011110 : OUT <= 7;  //233 / 30 = 7
    16'b11101001_00011111 : OUT <= 7;  //233 / 31 = 7
    16'b11101001_00100000 : OUT <= 7;  //233 / 32 = 7
    16'b11101001_00100001 : OUT <= 7;  //233 / 33 = 7
    16'b11101001_00100010 : OUT <= 6;  //233 / 34 = 6
    16'b11101001_00100011 : OUT <= 6;  //233 / 35 = 6
    16'b11101001_00100100 : OUT <= 6;  //233 / 36 = 6
    16'b11101001_00100101 : OUT <= 6;  //233 / 37 = 6
    16'b11101001_00100110 : OUT <= 6;  //233 / 38 = 6
    16'b11101001_00100111 : OUT <= 5;  //233 / 39 = 5
    16'b11101001_00101000 : OUT <= 5;  //233 / 40 = 5
    16'b11101001_00101001 : OUT <= 5;  //233 / 41 = 5
    16'b11101001_00101010 : OUT <= 5;  //233 / 42 = 5
    16'b11101001_00101011 : OUT <= 5;  //233 / 43 = 5
    16'b11101001_00101100 : OUT <= 5;  //233 / 44 = 5
    16'b11101001_00101101 : OUT <= 5;  //233 / 45 = 5
    16'b11101001_00101110 : OUT <= 5;  //233 / 46 = 5
    16'b11101001_00101111 : OUT <= 4;  //233 / 47 = 4
    16'b11101001_00110000 : OUT <= 4;  //233 / 48 = 4
    16'b11101001_00110001 : OUT <= 4;  //233 / 49 = 4
    16'b11101001_00110010 : OUT <= 4;  //233 / 50 = 4
    16'b11101001_00110011 : OUT <= 4;  //233 / 51 = 4
    16'b11101001_00110100 : OUT <= 4;  //233 / 52 = 4
    16'b11101001_00110101 : OUT <= 4;  //233 / 53 = 4
    16'b11101001_00110110 : OUT <= 4;  //233 / 54 = 4
    16'b11101001_00110111 : OUT <= 4;  //233 / 55 = 4
    16'b11101001_00111000 : OUT <= 4;  //233 / 56 = 4
    16'b11101001_00111001 : OUT <= 4;  //233 / 57 = 4
    16'b11101001_00111010 : OUT <= 4;  //233 / 58 = 4
    16'b11101001_00111011 : OUT <= 3;  //233 / 59 = 3
    16'b11101001_00111100 : OUT <= 3;  //233 / 60 = 3
    16'b11101001_00111101 : OUT <= 3;  //233 / 61 = 3
    16'b11101001_00111110 : OUT <= 3;  //233 / 62 = 3
    16'b11101001_00111111 : OUT <= 3;  //233 / 63 = 3
    16'b11101001_01000000 : OUT <= 3;  //233 / 64 = 3
    16'b11101001_01000001 : OUT <= 3;  //233 / 65 = 3
    16'b11101001_01000010 : OUT <= 3;  //233 / 66 = 3
    16'b11101001_01000011 : OUT <= 3;  //233 / 67 = 3
    16'b11101001_01000100 : OUT <= 3;  //233 / 68 = 3
    16'b11101001_01000101 : OUT <= 3;  //233 / 69 = 3
    16'b11101001_01000110 : OUT <= 3;  //233 / 70 = 3
    16'b11101001_01000111 : OUT <= 3;  //233 / 71 = 3
    16'b11101001_01001000 : OUT <= 3;  //233 / 72 = 3
    16'b11101001_01001001 : OUT <= 3;  //233 / 73 = 3
    16'b11101001_01001010 : OUT <= 3;  //233 / 74 = 3
    16'b11101001_01001011 : OUT <= 3;  //233 / 75 = 3
    16'b11101001_01001100 : OUT <= 3;  //233 / 76 = 3
    16'b11101001_01001101 : OUT <= 3;  //233 / 77 = 3
    16'b11101001_01001110 : OUT <= 2;  //233 / 78 = 2
    16'b11101001_01001111 : OUT <= 2;  //233 / 79 = 2
    16'b11101001_01010000 : OUT <= 2;  //233 / 80 = 2
    16'b11101001_01010001 : OUT <= 2;  //233 / 81 = 2
    16'b11101001_01010010 : OUT <= 2;  //233 / 82 = 2
    16'b11101001_01010011 : OUT <= 2;  //233 / 83 = 2
    16'b11101001_01010100 : OUT <= 2;  //233 / 84 = 2
    16'b11101001_01010101 : OUT <= 2;  //233 / 85 = 2
    16'b11101001_01010110 : OUT <= 2;  //233 / 86 = 2
    16'b11101001_01010111 : OUT <= 2;  //233 / 87 = 2
    16'b11101001_01011000 : OUT <= 2;  //233 / 88 = 2
    16'b11101001_01011001 : OUT <= 2;  //233 / 89 = 2
    16'b11101001_01011010 : OUT <= 2;  //233 / 90 = 2
    16'b11101001_01011011 : OUT <= 2;  //233 / 91 = 2
    16'b11101001_01011100 : OUT <= 2;  //233 / 92 = 2
    16'b11101001_01011101 : OUT <= 2;  //233 / 93 = 2
    16'b11101001_01011110 : OUT <= 2;  //233 / 94 = 2
    16'b11101001_01011111 : OUT <= 2;  //233 / 95 = 2
    16'b11101001_01100000 : OUT <= 2;  //233 / 96 = 2
    16'b11101001_01100001 : OUT <= 2;  //233 / 97 = 2
    16'b11101001_01100010 : OUT <= 2;  //233 / 98 = 2
    16'b11101001_01100011 : OUT <= 2;  //233 / 99 = 2
    16'b11101001_01100100 : OUT <= 2;  //233 / 100 = 2
    16'b11101001_01100101 : OUT <= 2;  //233 / 101 = 2
    16'b11101001_01100110 : OUT <= 2;  //233 / 102 = 2
    16'b11101001_01100111 : OUT <= 2;  //233 / 103 = 2
    16'b11101001_01101000 : OUT <= 2;  //233 / 104 = 2
    16'b11101001_01101001 : OUT <= 2;  //233 / 105 = 2
    16'b11101001_01101010 : OUT <= 2;  //233 / 106 = 2
    16'b11101001_01101011 : OUT <= 2;  //233 / 107 = 2
    16'b11101001_01101100 : OUT <= 2;  //233 / 108 = 2
    16'b11101001_01101101 : OUT <= 2;  //233 / 109 = 2
    16'b11101001_01101110 : OUT <= 2;  //233 / 110 = 2
    16'b11101001_01101111 : OUT <= 2;  //233 / 111 = 2
    16'b11101001_01110000 : OUT <= 2;  //233 / 112 = 2
    16'b11101001_01110001 : OUT <= 2;  //233 / 113 = 2
    16'b11101001_01110010 : OUT <= 2;  //233 / 114 = 2
    16'b11101001_01110011 : OUT <= 2;  //233 / 115 = 2
    16'b11101001_01110100 : OUT <= 2;  //233 / 116 = 2
    16'b11101001_01110101 : OUT <= 1;  //233 / 117 = 1
    16'b11101001_01110110 : OUT <= 1;  //233 / 118 = 1
    16'b11101001_01110111 : OUT <= 1;  //233 / 119 = 1
    16'b11101001_01111000 : OUT <= 1;  //233 / 120 = 1
    16'b11101001_01111001 : OUT <= 1;  //233 / 121 = 1
    16'b11101001_01111010 : OUT <= 1;  //233 / 122 = 1
    16'b11101001_01111011 : OUT <= 1;  //233 / 123 = 1
    16'b11101001_01111100 : OUT <= 1;  //233 / 124 = 1
    16'b11101001_01111101 : OUT <= 1;  //233 / 125 = 1
    16'b11101001_01111110 : OUT <= 1;  //233 / 126 = 1
    16'b11101001_01111111 : OUT <= 1;  //233 / 127 = 1
    16'b11101001_10000000 : OUT <= 1;  //233 / 128 = 1
    16'b11101001_10000001 : OUT <= 1;  //233 / 129 = 1
    16'b11101001_10000010 : OUT <= 1;  //233 / 130 = 1
    16'b11101001_10000011 : OUT <= 1;  //233 / 131 = 1
    16'b11101001_10000100 : OUT <= 1;  //233 / 132 = 1
    16'b11101001_10000101 : OUT <= 1;  //233 / 133 = 1
    16'b11101001_10000110 : OUT <= 1;  //233 / 134 = 1
    16'b11101001_10000111 : OUT <= 1;  //233 / 135 = 1
    16'b11101001_10001000 : OUT <= 1;  //233 / 136 = 1
    16'b11101001_10001001 : OUT <= 1;  //233 / 137 = 1
    16'b11101001_10001010 : OUT <= 1;  //233 / 138 = 1
    16'b11101001_10001011 : OUT <= 1;  //233 / 139 = 1
    16'b11101001_10001100 : OUT <= 1;  //233 / 140 = 1
    16'b11101001_10001101 : OUT <= 1;  //233 / 141 = 1
    16'b11101001_10001110 : OUT <= 1;  //233 / 142 = 1
    16'b11101001_10001111 : OUT <= 1;  //233 / 143 = 1
    16'b11101001_10010000 : OUT <= 1;  //233 / 144 = 1
    16'b11101001_10010001 : OUT <= 1;  //233 / 145 = 1
    16'b11101001_10010010 : OUT <= 1;  //233 / 146 = 1
    16'b11101001_10010011 : OUT <= 1;  //233 / 147 = 1
    16'b11101001_10010100 : OUT <= 1;  //233 / 148 = 1
    16'b11101001_10010101 : OUT <= 1;  //233 / 149 = 1
    16'b11101001_10010110 : OUT <= 1;  //233 / 150 = 1
    16'b11101001_10010111 : OUT <= 1;  //233 / 151 = 1
    16'b11101001_10011000 : OUT <= 1;  //233 / 152 = 1
    16'b11101001_10011001 : OUT <= 1;  //233 / 153 = 1
    16'b11101001_10011010 : OUT <= 1;  //233 / 154 = 1
    16'b11101001_10011011 : OUT <= 1;  //233 / 155 = 1
    16'b11101001_10011100 : OUT <= 1;  //233 / 156 = 1
    16'b11101001_10011101 : OUT <= 1;  //233 / 157 = 1
    16'b11101001_10011110 : OUT <= 1;  //233 / 158 = 1
    16'b11101001_10011111 : OUT <= 1;  //233 / 159 = 1
    16'b11101001_10100000 : OUT <= 1;  //233 / 160 = 1
    16'b11101001_10100001 : OUT <= 1;  //233 / 161 = 1
    16'b11101001_10100010 : OUT <= 1;  //233 / 162 = 1
    16'b11101001_10100011 : OUT <= 1;  //233 / 163 = 1
    16'b11101001_10100100 : OUT <= 1;  //233 / 164 = 1
    16'b11101001_10100101 : OUT <= 1;  //233 / 165 = 1
    16'b11101001_10100110 : OUT <= 1;  //233 / 166 = 1
    16'b11101001_10100111 : OUT <= 1;  //233 / 167 = 1
    16'b11101001_10101000 : OUT <= 1;  //233 / 168 = 1
    16'b11101001_10101001 : OUT <= 1;  //233 / 169 = 1
    16'b11101001_10101010 : OUT <= 1;  //233 / 170 = 1
    16'b11101001_10101011 : OUT <= 1;  //233 / 171 = 1
    16'b11101001_10101100 : OUT <= 1;  //233 / 172 = 1
    16'b11101001_10101101 : OUT <= 1;  //233 / 173 = 1
    16'b11101001_10101110 : OUT <= 1;  //233 / 174 = 1
    16'b11101001_10101111 : OUT <= 1;  //233 / 175 = 1
    16'b11101001_10110000 : OUT <= 1;  //233 / 176 = 1
    16'b11101001_10110001 : OUT <= 1;  //233 / 177 = 1
    16'b11101001_10110010 : OUT <= 1;  //233 / 178 = 1
    16'b11101001_10110011 : OUT <= 1;  //233 / 179 = 1
    16'b11101001_10110100 : OUT <= 1;  //233 / 180 = 1
    16'b11101001_10110101 : OUT <= 1;  //233 / 181 = 1
    16'b11101001_10110110 : OUT <= 1;  //233 / 182 = 1
    16'b11101001_10110111 : OUT <= 1;  //233 / 183 = 1
    16'b11101001_10111000 : OUT <= 1;  //233 / 184 = 1
    16'b11101001_10111001 : OUT <= 1;  //233 / 185 = 1
    16'b11101001_10111010 : OUT <= 1;  //233 / 186 = 1
    16'b11101001_10111011 : OUT <= 1;  //233 / 187 = 1
    16'b11101001_10111100 : OUT <= 1;  //233 / 188 = 1
    16'b11101001_10111101 : OUT <= 1;  //233 / 189 = 1
    16'b11101001_10111110 : OUT <= 1;  //233 / 190 = 1
    16'b11101001_10111111 : OUT <= 1;  //233 / 191 = 1
    16'b11101001_11000000 : OUT <= 1;  //233 / 192 = 1
    16'b11101001_11000001 : OUT <= 1;  //233 / 193 = 1
    16'b11101001_11000010 : OUT <= 1;  //233 / 194 = 1
    16'b11101001_11000011 : OUT <= 1;  //233 / 195 = 1
    16'b11101001_11000100 : OUT <= 1;  //233 / 196 = 1
    16'b11101001_11000101 : OUT <= 1;  //233 / 197 = 1
    16'b11101001_11000110 : OUT <= 1;  //233 / 198 = 1
    16'b11101001_11000111 : OUT <= 1;  //233 / 199 = 1
    16'b11101001_11001000 : OUT <= 1;  //233 / 200 = 1
    16'b11101001_11001001 : OUT <= 1;  //233 / 201 = 1
    16'b11101001_11001010 : OUT <= 1;  //233 / 202 = 1
    16'b11101001_11001011 : OUT <= 1;  //233 / 203 = 1
    16'b11101001_11001100 : OUT <= 1;  //233 / 204 = 1
    16'b11101001_11001101 : OUT <= 1;  //233 / 205 = 1
    16'b11101001_11001110 : OUT <= 1;  //233 / 206 = 1
    16'b11101001_11001111 : OUT <= 1;  //233 / 207 = 1
    16'b11101001_11010000 : OUT <= 1;  //233 / 208 = 1
    16'b11101001_11010001 : OUT <= 1;  //233 / 209 = 1
    16'b11101001_11010010 : OUT <= 1;  //233 / 210 = 1
    16'b11101001_11010011 : OUT <= 1;  //233 / 211 = 1
    16'b11101001_11010100 : OUT <= 1;  //233 / 212 = 1
    16'b11101001_11010101 : OUT <= 1;  //233 / 213 = 1
    16'b11101001_11010110 : OUT <= 1;  //233 / 214 = 1
    16'b11101001_11010111 : OUT <= 1;  //233 / 215 = 1
    16'b11101001_11011000 : OUT <= 1;  //233 / 216 = 1
    16'b11101001_11011001 : OUT <= 1;  //233 / 217 = 1
    16'b11101001_11011010 : OUT <= 1;  //233 / 218 = 1
    16'b11101001_11011011 : OUT <= 1;  //233 / 219 = 1
    16'b11101001_11011100 : OUT <= 1;  //233 / 220 = 1
    16'b11101001_11011101 : OUT <= 1;  //233 / 221 = 1
    16'b11101001_11011110 : OUT <= 1;  //233 / 222 = 1
    16'b11101001_11011111 : OUT <= 1;  //233 / 223 = 1
    16'b11101001_11100000 : OUT <= 1;  //233 / 224 = 1
    16'b11101001_11100001 : OUT <= 1;  //233 / 225 = 1
    16'b11101001_11100010 : OUT <= 1;  //233 / 226 = 1
    16'b11101001_11100011 : OUT <= 1;  //233 / 227 = 1
    16'b11101001_11100100 : OUT <= 1;  //233 / 228 = 1
    16'b11101001_11100101 : OUT <= 1;  //233 / 229 = 1
    16'b11101001_11100110 : OUT <= 1;  //233 / 230 = 1
    16'b11101001_11100111 : OUT <= 1;  //233 / 231 = 1
    16'b11101001_11101000 : OUT <= 1;  //233 / 232 = 1
    16'b11101001_11101001 : OUT <= 1;  //233 / 233 = 1
    16'b11101001_11101010 : OUT <= 0;  //233 / 234 = 0
    16'b11101001_11101011 : OUT <= 0;  //233 / 235 = 0
    16'b11101001_11101100 : OUT <= 0;  //233 / 236 = 0
    16'b11101001_11101101 : OUT <= 0;  //233 / 237 = 0
    16'b11101001_11101110 : OUT <= 0;  //233 / 238 = 0
    16'b11101001_11101111 : OUT <= 0;  //233 / 239 = 0
    16'b11101001_11110000 : OUT <= 0;  //233 / 240 = 0
    16'b11101001_11110001 : OUT <= 0;  //233 / 241 = 0
    16'b11101001_11110010 : OUT <= 0;  //233 / 242 = 0
    16'b11101001_11110011 : OUT <= 0;  //233 / 243 = 0
    16'b11101001_11110100 : OUT <= 0;  //233 / 244 = 0
    16'b11101001_11110101 : OUT <= 0;  //233 / 245 = 0
    16'b11101001_11110110 : OUT <= 0;  //233 / 246 = 0
    16'b11101001_11110111 : OUT <= 0;  //233 / 247 = 0
    16'b11101001_11111000 : OUT <= 0;  //233 / 248 = 0
    16'b11101001_11111001 : OUT <= 0;  //233 / 249 = 0
    16'b11101001_11111010 : OUT <= 0;  //233 / 250 = 0
    16'b11101001_11111011 : OUT <= 0;  //233 / 251 = 0
    16'b11101001_11111100 : OUT <= 0;  //233 / 252 = 0
    16'b11101001_11111101 : OUT <= 0;  //233 / 253 = 0
    16'b11101001_11111110 : OUT <= 0;  //233 / 254 = 0
    16'b11101001_11111111 : OUT <= 0;  //233 / 255 = 0
    16'b11101010_00000000 : OUT <= 0;  //234 / 0 = 0
    16'b11101010_00000001 : OUT <= 234;  //234 / 1 = 234
    16'b11101010_00000010 : OUT <= 117;  //234 / 2 = 117
    16'b11101010_00000011 : OUT <= 78;  //234 / 3 = 78
    16'b11101010_00000100 : OUT <= 58;  //234 / 4 = 58
    16'b11101010_00000101 : OUT <= 46;  //234 / 5 = 46
    16'b11101010_00000110 : OUT <= 39;  //234 / 6 = 39
    16'b11101010_00000111 : OUT <= 33;  //234 / 7 = 33
    16'b11101010_00001000 : OUT <= 29;  //234 / 8 = 29
    16'b11101010_00001001 : OUT <= 26;  //234 / 9 = 26
    16'b11101010_00001010 : OUT <= 23;  //234 / 10 = 23
    16'b11101010_00001011 : OUT <= 21;  //234 / 11 = 21
    16'b11101010_00001100 : OUT <= 19;  //234 / 12 = 19
    16'b11101010_00001101 : OUT <= 18;  //234 / 13 = 18
    16'b11101010_00001110 : OUT <= 16;  //234 / 14 = 16
    16'b11101010_00001111 : OUT <= 15;  //234 / 15 = 15
    16'b11101010_00010000 : OUT <= 14;  //234 / 16 = 14
    16'b11101010_00010001 : OUT <= 13;  //234 / 17 = 13
    16'b11101010_00010010 : OUT <= 13;  //234 / 18 = 13
    16'b11101010_00010011 : OUT <= 12;  //234 / 19 = 12
    16'b11101010_00010100 : OUT <= 11;  //234 / 20 = 11
    16'b11101010_00010101 : OUT <= 11;  //234 / 21 = 11
    16'b11101010_00010110 : OUT <= 10;  //234 / 22 = 10
    16'b11101010_00010111 : OUT <= 10;  //234 / 23 = 10
    16'b11101010_00011000 : OUT <= 9;  //234 / 24 = 9
    16'b11101010_00011001 : OUT <= 9;  //234 / 25 = 9
    16'b11101010_00011010 : OUT <= 9;  //234 / 26 = 9
    16'b11101010_00011011 : OUT <= 8;  //234 / 27 = 8
    16'b11101010_00011100 : OUT <= 8;  //234 / 28 = 8
    16'b11101010_00011101 : OUT <= 8;  //234 / 29 = 8
    16'b11101010_00011110 : OUT <= 7;  //234 / 30 = 7
    16'b11101010_00011111 : OUT <= 7;  //234 / 31 = 7
    16'b11101010_00100000 : OUT <= 7;  //234 / 32 = 7
    16'b11101010_00100001 : OUT <= 7;  //234 / 33 = 7
    16'b11101010_00100010 : OUT <= 6;  //234 / 34 = 6
    16'b11101010_00100011 : OUT <= 6;  //234 / 35 = 6
    16'b11101010_00100100 : OUT <= 6;  //234 / 36 = 6
    16'b11101010_00100101 : OUT <= 6;  //234 / 37 = 6
    16'b11101010_00100110 : OUT <= 6;  //234 / 38 = 6
    16'b11101010_00100111 : OUT <= 6;  //234 / 39 = 6
    16'b11101010_00101000 : OUT <= 5;  //234 / 40 = 5
    16'b11101010_00101001 : OUT <= 5;  //234 / 41 = 5
    16'b11101010_00101010 : OUT <= 5;  //234 / 42 = 5
    16'b11101010_00101011 : OUT <= 5;  //234 / 43 = 5
    16'b11101010_00101100 : OUT <= 5;  //234 / 44 = 5
    16'b11101010_00101101 : OUT <= 5;  //234 / 45 = 5
    16'b11101010_00101110 : OUT <= 5;  //234 / 46 = 5
    16'b11101010_00101111 : OUT <= 4;  //234 / 47 = 4
    16'b11101010_00110000 : OUT <= 4;  //234 / 48 = 4
    16'b11101010_00110001 : OUT <= 4;  //234 / 49 = 4
    16'b11101010_00110010 : OUT <= 4;  //234 / 50 = 4
    16'b11101010_00110011 : OUT <= 4;  //234 / 51 = 4
    16'b11101010_00110100 : OUT <= 4;  //234 / 52 = 4
    16'b11101010_00110101 : OUT <= 4;  //234 / 53 = 4
    16'b11101010_00110110 : OUT <= 4;  //234 / 54 = 4
    16'b11101010_00110111 : OUT <= 4;  //234 / 55 = 4
    16'b11101010_00111000 : OUT <= 4;  //234 / 56 = 4
    16'b11101010_00111001 : OUT <= 4;  //234 / 57 = 4
    16'b11101010_00111010 : OUT <= 4;  //234 / 58 = 4
    16'b11101010_00111011 : OUT <= 3;  //234 / 59 = 3
    16'b11101010_00111100 : OUT <= 3;  //234 / 60 = 3
    16'b11101010_00111101 : OUT <= 3;  //234 / 61 = 3
    16'b11101010_00111110 : OUT <= 3;  //234 / 62 = 3
    16'b11101010_00111111 : OUT <= 3;  //234 / 63 = 3
    16'b11101010_01000000 : OUT <= 3;  //234 / 64 = 3
    16'b11101010_01000001 : OUT <= 3;  //234 / 65 = 3
    16'b11101010_01000010 : OUT <= 3;  //234 / 66 = 3
    16'b11101010_01000011 : OUT <= 3;  //234 / 67 = 3
    16'b11101010_01000100 : OUT <= 3;  //234 / 68 = 3
    16'b11101010_01000101 : OUT <= 3;  //234 / 69 = 3
    16'b11101010_01000110 : OUT <= 3;  //234 / 70 = 3
    16'b11101010_01000111 : OUT <= 3;  //234 / 71 = 3
    16'b11101010_01001000 : OUT <= 3;  //234 / 72 = 3
    16'b11101010_01001001 : OUT <= 3;  //234 / 73 = 3
    16'b11101010_01001010 : OUT <= 3;  //234 / 74 = 3
    16'b11101010_01001011 : OUT <= 3;  //234 / 75 = 3
    16'b11101010_01001100 : OUT <= 3;  //234 / 76 = 3
    16'b11101010_01001101 : OUT <= 3;  //234 / 77 = 3
    16'b11101010_01001110 : OUT <= 3;  //234 / 78 = 3
    16'b11101010_01001111 : OUT <= 2;  //234 / 79 = 2
    16'b11101010_01010000 : OUT <= 2;  //234 / 80 = 2
    16'b11101010_01010001 : OUT <= 2;  //234 / 81 = 2
    16'b11101010_01010010 : OUT <= 2;  //234 / 82 = 2
    16'b11101010_01010011 : OUT <= 2;  //234 / 83 = 2
    16'b11101010_01010100 : OUT <= 2;  //234 / 84 = 2
    16'b11101010_01010101 : OUT <= 2;  //234 / 85 = 2
    16'b11101010_01010110 : OUT <= 2;  //234 / 86 = 2
    16'b11101010_01010111 : OUT <= 2;  //234 / 87 = 2
    16'b11101010_01011000 : OUT <= 2;  //234 / 88 = 2
    16'b11101010_01011001 : OUT <= 2;  //234 / 89 = 2
    16'b11101010_01011010 : OUT <= 2;  //234 / 90 = 2
    16'b11101010_01011011 : OUT <= 2;  //234 / 91 = 2
    16'b11101010_01011100 : OUT <= 2;  //234 / 92 = 2
    16'b11101010_01011101 : OUT <= 2;  //234 / 93 = 2
    16'b11101010_01011110 : OUT <= 2;  //234 / 94 = 2
    16'b11101010_01011111 : OUT <= 2;  //234 / 95 = 2
    16'b11101010_01100000 : OUT <= 2;  //234 / 96 = 2
    16'b11101010_01100001 : OUT <= 2;  //234 / 97 = 2
    16'b11101010_01100010 : OUT <= 2;  //234 / 98 = 2
    16'b11101010_01100011 : OUT <= 2;  //234 / 99 = 2
    16'b11101010_01100100 : OUT <= 2;  //234 / 100 = 2
    16'b11101010_01100101 : OUT <= 2;  //234 / 101 = 2
    16'b11101010_01100110 : OUT <= 2;  //234 / 102 = 2
    16'b11101010_01100111 : OUT <= 2;  //234 / 103 = 2
    16'b11101010_01101000 : OUT <= 2;  //234 / 104 = 2
    16'b11101010_01101001 : OUT <= 2;  //234 / 105 = 2
    16'b11101010_01101010 : OUT <= 2;  //234 / 106 = 2
    16'b11101010_01101011 : OUT <= 2;  //234 / 107 = 2
    16'b11101010_01101100 : OUT <= 2;  //234 / 108 = 2
    16'b11101010_01101101 : OUT <= 2;  //234 / 109 = 2
    16'b11101010_01101110 : OUT <= 2;  //234 / 110 = 2
    16'b11101010_01101111 : OUT <= 2;  //234 / 111 = 2
    16'b11101010_01110000 : OUT <= 2;  //234 / 112 = 2
    16'b11101010_01110001 : OUT <= 2;  //234 / 113 = 2
    16'b11101010_01110010 : OUT <= 2;  //234 / 114 = 2
    16'b11101010_01110011 : OUT <= 2;  //234 / 115 = 2
    16'b11101010_01110100 : OUT <= 2;  //234 / 116 = 2
    16'b11101010_01110101 : OUT <= 2;  //234 / 117 = 2
    16'b11101010_01110110 : OUT <= 1;  //234 / 118 = 1
    16'b11101010_01110111 : OUT <= 1;  //234 / 119 = 1
    16'b11101010_01111000 : OUT <= 1;  //234 / 120 = 1
    16'b11101010_01111001 : OUT <= 1;  //234 / 121 = 1
    16'b11101010_01111010 : OUT <= 1;  //234 / 122 = 1
    16'b11101010_01111011 : OUT <= 1;  //234 / 123 = 1
    16'b11101010_01111100 : OUT <= 1;  //234 / 124 = 1
    16'b11101010_01111101 : OUT <= 1;  //234 / 125 = 1
    16'b11101010_01111110 : OUT <= 1;  //234 / 126 = 1
    16'b11101010_01111111 : OUT <= 1;  //234 / 127 = 1
    16'b11101010_10000000 : OUT <= 1;  //234 / 128 = 1
    16'b11101010_10000001 : OUT <= 1;  //234 / 129 = 1
    16'b11101010_10000010 : OUT <= 1;  //234 / 130 = 1
    16'b11101010_10000011 : OUT <= 1;  //234 / 131 = 1
    16'b11101010_10000100 : OUT <= 1;  //234 / 132 = 1
    16'b11101010_10000101 : OUT <= 1;  //234 / 133 = 1
    16'b11101010_10000110 : OUT <= 1;  //234 / 134 = 1
    16'b11101010_10000111 : OUT <= 1;  //234 / 135 = 1
    16'b11101010_10001000 : OUT <= 1;  //234 / 136 = 1
    16'b11101010_10001001 : OUT <= 1;  //234 / 137 = 1
    16'b11101010_10001010 : OUT <= 1;  //234 / 138 = 1
    16'b11101010_10001011 : OUT <= 1;  //234 / 139 = 1
    16'b11101010_10001100 : OUT <= 1;  //234 / 140 = 1
    16'b11101010_10001101 : OUT <= 1;  //234 / 141 = 1
    16'b11101010_10001110 : OUT <= 1;  //234 / 142 = 1
    16'b11101010_10001111 : OUT <= 1;  //234 / 143 = 1
    16'b11101010_10010000 : OUT <= 1;  //234 / 144 = 1
    16'b11101010_10010001 : OUT <= 1;  //234 / 145 = 1
    16'b11101010_10010010 : OUT <= 1;  //234 / 146 = 1
    16'b11101010_10010011 : OUT <= 1;  //234 / 147 = 1
    16'b11101010_10010100 : OUT <= 1;  //234 / 148 = 1
    16'b11101010_10010101 : OUT <= 1;  //234 / 149 = 1
    16'b11101010_10010110 : OUT <= 1;  //234 / 150 = 1
    16'b11101010_10010111 : OUT <= 1;  //234 / 151 = 1
    16'b11101010_10011000 : OUT <= 1;  //234 / 152 = 1
    16'b11101010_10011001 : OUT <= 1;  //234 / 153 = 1
    16'b11101010_10011010 : OUT <= 1;  //234 / 154 = 1
    16'b11101010_10011011 : OUT <= 1;  //234 / 155 = 1
    16'b11101010_10011100 : OUT <= 1;  //234 / 156 = 1
    16'b11101010_10011101 : OUT <= 1;  //234 / 157 = 1
    16'b11101010_10011110 : OUT <= 1;  //234 / 158 = 1
    16'b11101010_10011111 : OUT <= 1;  //234 / 159 = 1
    16'b11101010_10100000 : OUT <= 1;  //234 / 160 = 1
    16'b11101010_10100001 : OUT <= 1;  //234 / 161 = 1
    16'b11101010_10100010 : OUT <= 1;  //234 / 162 = 1
    16'b11101010_10100011 : OUT <= 1;  //234 / 163 = 1
    16'b11101010_10100100 : OUT <= 1;  //234 / 164 = 1
    16'b11101010_10100101 : OUT <= 1;  //234 / 165 = 1
    16'b11101010_10100110 : OUT <= 1;  //234 / 166 = 1
    16'b11101010_10100111 : OUT <= 1;  //234 / 167 = 1
    16'b11101010_10101000 : OUT <= 1;  //234 / 168 = 1
    16'b11101010_10101001 : OUT <= 1;  //234 / 169 = 1
    16'b11101010_10101010 : OUT <= 1;  //234 / 170 = 1
    16'b11101010_10101011 : OUT <= 1;  //234 / 171 = 1
    16'b11101010_10101100 : OUT <= 1;  //234 / 172 = 1
    16'b11101010_10101101 : OUT <= 1;  //234 / 173 = 1
    16'b11101010_10101110 : OUT <= 1;  //234 / 174 = 1
    16'b11101010_10101111 : OUT <= 1;  //234 / 175 = 1
    16'b11101010_10110000 : OUT <= 1;  //234 / 176 = 1
    16'b11101010_10110001 : OUT <= 1;  //234 / 177 = 1
    16'b11101010_10110010 : OUT <= 1;  //234 / 178 = 1
    16'b11101010_10110011 : OUT <= 1;  //234 / 179 = 1
    16'b11101010_10110100 : OUT <= 1;  //234 / 180 = 1
    16'b11101010_10110101 : OUT <= 1;  //234 / 181 = 1
    16'b11101010_10110110 : OUT <= 1;  //234 / 182 = 1
    16'b11101010_10110111 : OUT <= 1;  //234 / 183 = 1
    16'b11101010_10111000 : OUT <= 1;  //234 / 184 = 1
    16'b11101010_10111001 : OUT <= 1;  //234 / 185 = 1
    16'b11101010_10111010 : OUT <= 1;  //234 / 186 = 1
    16'b11101010_10111011 : OUT <= 1;  //234 / 187 = 1
    16'b11101010_10111100 : OUT <= 1;  //234 / 188 = 1
    16'b11101010_10111101 : OUT <= 1;  //234 / 189 = 1
    16'b11101010_10111110 : OUT <= 1;  //234 / 190 = 1
    16'b11101010_10111111 : OUT <= 1;  //234 / 191 = 1
    16'b11101010_11000000 : OUT <= 1;  //234 / 192 = 1
    16'b11101010_11000001 : OUT <= 1;  //234 / 193 = 1
    16'b11101010_11000010 : OUT <= 1;  //234 / 194 = 1
    16'b11101010_11000011 : OUT <= 1;  //234 / 195 = 1
    16'b11101010_11000100 : OUT <= 1;  //234 / 196 = 1
    16'b11101010_11000101 : OUT <= 1;  //234 / 197 = 1
    16'b11101010_11000110 : OUT <= 1;  //234 / 198 = 1
    16'b11101010_11000111 : OUT <= 1;  //234 / 199 = 1
    16'b11101010_11001000 : OUT <= 1;  //234 / 200 = 1
    16'b11101010_11001001 : OUT <= 1;  //234 / 201 = 1
    16'b11101010_11001010 : OUT <= 1;  //234 / 202 = 1
    16'b11101010_11001011 : OUT <= 1;  //234 / 203 = 1
    16'b11101010_11001100 : OUT <= 1;  //234 / 204 = 1
    16'b11101010_11001101 : OUT <= 1;  //234 / 205 = 1
    16'b11101010_11001110 : OUT <= 1;  //234 / 206 = 1
    16'b11101010_11001111 : OUT <= 1;  //234 / 207 = 1
    16'b11101010_11010000 : OUT <= 1;  //234 / 208 = 1
    16'b11101010_11010001 : OUT <= 1;  //234 / 209 = 1
    16'b11101010_11010010 : OUT <= 1;  //234 / 210 = 1
    16'b11101010_11010011 : OUT <= 1;  //234 / 211 = 1
    16'b11101010_11010100 : OUT <= 1;  //234 / 212 = 1
    16'b11101010_11010101 : OUT <= 1;  //234 / 213 = 1
    16'b11101010_11010110 : OUT <= 1;  //234 / 214 = 1
    16'b11101010_11010111 : OUT <= 1;  //234 / 215 = 1
    16'b11101010_11011000 : OUT <= 1;  //234 / 216 = 1
    16'b11101010_11011001 : OUT <= 1;  //234 / 217 = 1
    16'b11101010_11011010 : OUT <= 1;  //234 / 218 = 1
    16'b11101010_11011011 : OUT <= 1;  //234 / 219 = 1
    16'b11101010_11011100 : OUT <= 1;  //234 / 220 = 1
    16'b11101010_11011101 : OUT <= 1;  //234 / 221 = 1
    16'b11101010_11011110 : OUT <= 1;  //234 / 222 = 1
    16'b11101010_11011111 : OUT <= 1;  //234 / 223 = 1
    16'b11101010_11100000 : OUT <= 1;  //234 / 224 = 1
    16'b11101010_11100001 : OUT <= 1;  //234 / 225 = 1
    16'b11101010_11100010 : OUT <= 1;  //234 / 226 = 1
    16'b11101010_11100011 : OUT <= 1;  //234 / 227 = 1
    16'b11101010_11100100 : OUT <= 1;  //234 / 228 = 1
    16'b11101010_11100101 : OUT <= 1;  //234 / 229 = 1
    16'b11101010_11100110 : OUT <= 1;  //234 / 230 = 1
    16'b11101010_11100111 : OUT <= 1;  //234 / 231 = 1
    16'b11101010_11101000 : OUT <= 1;  //234 / 232 = 1
    16'b11101010_11101001 : OUT <= 1;  //234 / 233 = 1
    16'b11101010_11101010 : OUT <= 1;  //234 / 234 = 1
    16'b11101010_11101011 : OUT <= 0;  //234 / 235 = 0
    16'b11101010_11101100 : OUT <= 0;  //234 / 236 = 0
    16'b11101010_11101101 : OUT <= 0;  //234 / 237 = 0
    16'b11101010_11101110 : OUT <= 0;  //234 / 238 = 0
    16'b11101010_11101111 : OUT <= 0;  //234 / 239 = 0
    16'b11101010_11110000 : OUT <= 0;  //234 / 240 = 0
    16'b11101010_11110001 : OUT <= 0;  //234 / 241 = 0
    16'b11101010_11110010 : OUT <= 0;  //234 / 242 = 0
    16'b11101010_11110011 : OUT <= 0;  //234 / 243 = 0
    16'b11101010_11110100 : OUT <= 0;  //234 / 244 = 0
    16'b11101010_11110101 : OUT <= 0;  //234 / 245 = 0
    16'b11101010_11110110 : OUT <= 0;  //234 / 246 = 0
    16'b11101010_11110111 : OUT <= 0;  //234 / 247 = 0
    16'b11101010_11111000 : OUT <= 0;  //234 / 248 = 0
    16'b11101010_11111001 : OUT <= 0;  //234 / 249 = 0
    16'b11101010_11111010 : OUT <= 0;  //234 / 250 = 0
    16'b11101010_11111011 : OUT <= 0;  //234 / 251 = 0
    16'b11101010_11111100 : OUT <= 0;  //234 / 252 = 0
    16'b11101010_11111101 : OUT <= 0;  //234 / 253 = 0
    16'b11101010_11111110 : OUT <= 0;  //234 / 254 = 0
    16'b11101010_11111111 : OUT <= 0;  //234 / 255 = 0
    16'b11101011_00000000 : OUT <= 0;  //235 / 0 = 0
    16'b11101011_00000001 : OUT <= 235;  //235 / 1 = 235
    16'b11101011_00000010 : OUT <= 117;  //235 / 2 = 117
    16'b11101011_00000011 : OUT <= 78;  //235 / 3 = 78
    16'b11101011_00000100 : OUT <= 58;  //235 / 4 = 58
    16'b11101011_00000101 : OUT <= 47;  //235 / 5 = 47
    16'b11101011_00000110 : OUT <= 39;  //235 / 6 = 39
    16'b11101011_00000111 : OUT <= 33;  //235 / 7 = 33
    16'b11101011_00001000 : OUT <= 29;  //235 / 8 = 29
    16'b11101011_00001001 : OUT <= 26;  //235 / 9 = 26
    16'b11101011_00001010 : OUT <= 23;  //235 / 10 = 23
    16'b11101011_00001011 : OUT <= 21;  //235 / 11 = 21
    16'b11101011_00001100 : OUT <= 19;  //235 / 12 = 19
    16'b11101011_00001101 : OUT <= 18;  //235 / 13 = 18
    16'b11101011_00001110 : OUT <= 16;  //235 / 14 = 16
    16'b11101011_00001111 : OUT <= 15;  //235 / 15 = 15
    16'b11101011_00010000 : OUT <= 14;  //235 / 16 = 14
    16'b11101011_00010001 : OUT <= 13;  //235 / 17 = 13
    16'b11101011_00010010 : OUT <= 13;  //235 / 18 = 13
    16'b11101011_00010011 : OUT <= 12;  //235 / 19 = 12
    16'b11101011_00010100 : OUT <= 11;  //235 / 20 = 11
    16'b11101011_00010101 : OUT <= 11;  //235 / 21 = 11
    16'b11101011_00010110 : OUT <= 10;  //235 / 22 = 10
    16'b11101011_00010111 : OUT <= 10;  //235 / 23 = 10
    16'b11101011_00011000 : OUT <= 9;  //235 / 24 = 9
    16'b11101011_00011001 : OUT <= 9;  //235 / 25 = 9
    16'b11101011_00011010 : OUT <= 9;  //235 / 26 = 9
    16'b11101011_00011011 : OUT <= 8;  //235 / 27 = 8
    16'b11101011_00011100 : OUT <= 8;  //235 / 28 = 8
    16'b11101011_00011101 : OUT <= 8;  //235 / 29 = 8
    16'b11101011_00011110 : OUT <= 7;  //235 / 30 = 7
    16'b11101011_00011111 : OUT <= 7;  //235 / 31 = 7
    16'b11101011_00100000 : OUT <= 7;  //235 / 32 = 7
    16'b11101011_00100001 : OUT <= 7;  //235 / 33 = 7
    16'b11101011_00100010 : OUT <= 6;  //235 / 34 = 6
    16'b11101011_00100011 : OUT <= 6;  //235 / 35 = 6
    16'b11101011_00100100 : OUT <= 6;  //235 / 36 = 6
    16'b11101011_00100101 : OUT <= 6;  //235 / 37 = 6
    16'b11101011_00100110 : OUT <= 6;  //235 / 38 = 6
    16'b11101011_00100111 : OUT <= 6;  //235 / 39 = 6
    16'b11101011_00101000 : OUT <= 5;  //235 / 40 = 5
    16'b11101011_00101001 : OUT <= 5;  //235 / 41 = 5
    16'b11101011_00101010 : OUT <= 5;  //235 / 42 = 5
    16'b11101011_00101011 : OUT <= 5;  //235 / 43 = 5
    16'b11101011_00101100 : OUT <= 5;  //235 / 44 = 5
    16'b11101011_00101101 : OUT <= 5;  //235 / 45 = 5
    16'b11101011_00101110 : OUT <= 5;  //235 / 46 = 5
    16'b11101011_00101111 : OUT <= 5;  //235 / 47 = 5
    16'b11101011_00110000 : OUT <= 4;  //235 / 48 = 4
    16'b11101011_00110001 : OUT <= 4;  //235 / 49 = 4
    16'b11101011_00110010 : OUT <= 4;  //235 / 50 = 4
    16'b11101011_00110011 : OUT <= 4;  //235 / 51 = 4
    16'b11101011_00110100 : OUT <= 4;  //235 / 52 = 4
    16'b11101011_00110101 : OUT <= 4;  //235 / 53 = 4
    16'b11101011_00110110 : OUT <= 4;  //235 / 54 = 4
    16'b11101011_00110111 : OUT <= 4;  //235 / 55 = 4
    16'b11101011_00111000 : OUT <= 4;  //235 / 56 = 4
    16'b11101011_00111001 : OUT <= 4;  //235 / 57 = 4
    16'b11101011_00111010 : OUT <= 4;  //235 / 58 = 4
    16'b11101011_00111011 : OUT <= 3;  //235 / 59 = 3
    16'b11101011_00111100 : OUT <= 3;  //235 / 60 = 3
    16'b11101011_00111101 : OUT <= 3;  //235 / 61 = 3
    16'b11101011_00111110 : OUT <= 3;  //235 / 62 = 3
    16'b11101011_00111111 : OUT <= 3;  //235 / 63 = 3
    16'b11101011_01000000 : OUT <= 3;  //235 / 64 = 3
    16'b11101011_01000001 : OUT <= 3;  //235 / 65 = 3
    16'b11101011_01000010 : OUT <= 3;  //235 / 66 = 3
    16'b11101011_01000011 : OUT <= 3;  //235 / 67 = 3
    16'b11101011_01000100 : OUT <= 3;  //235 / 68 = 3
    16'b11101011_01000101 : OUT <= 3;  //235 / 69 = 3
    16'b11101011_01000110 : OUT <= 3;  //235 / 70 = 3
    16'b11101011_01000111 : OUT <= 3;  //235 / 71 = 3
    16'b11101011_01001000 : OUT <= 3;  //235 / 72 = 3
    16'b11101011_01001001 : OUT <= 3;  //235 / 73 = 3
    16'b11101011_01001010 : OUT <= 3;  //235 / 74 = 3
    16'b11101011_01001011 : OUT <= 3;  //235 / 75 = 3
    16'b11101011_01001100 : OUT <= 3;  //235 / 76 = 3
    16'b11101011_01001101 : OUT <= 3;  //235 / 77 = 3
    16'b11101011_01001110 : OUT <= 3;  //235 / 78 = 3
    16'b11101011_01001111 : OUT <= 2;  //235 / 79 = 2
    16'b11101011_01010000 : OUT <= 2;  //235 / 80 = 2
    16'b11101011_01010001 : OUT <= 2;  //235 / 81 = 2
    16'b11101011_01010010 : OUT <= 2;  //235 / 82 = 2
    16'b11101011_01010011 : OUT <= 2;  //235 / 83 = 2
    16'b11101011_01010100 : OUT <= 2;  //235 / 84 = 2
    16'b11101011_01010101 : OUT <= 2;  //235 / 85 = 2
    16'b11101011_01010110 : OUT <= 2;  //235 / 86 = 2
    16'b11101011_01010111 : OUT <= 2;  //235 / 87 = 2
    16'b11101011_01011000 : OUT <= 2;  //235 / 88 = 2
    16'b11101011_01011001 : OUT <= 2;  //235 / 89 = 2
    16'b11101011_01011010 : OUT <= 2;  //235 / 90 = 2
    16'b11101011_01011011 : OUT <= 2;  //235 / 91 = 2
    16'b11101011_01011100 : OUT <= 2;  //235 / 92 = 2
    16'b11101011_01011101 : OUT <= 2;  //235 / 93 = 2
    16'b11101011_01011110 : OUT <= 2;  //235 / 94 = 2
    16'b11101011_01011111 : OUT <= 2;  //235 / 95 = 2
    16'b11101011_01100000 : OUT <= 2;  //235 / 96 = 2
    16'b11101011_01100001 : OUT <= 2;  //235 / 97 = 2
    16'b11101011_01100010 : OUT <= 2;  //235 / 98 = 2
    16'b11101011_01100011 : OUT <= 2;  //235 / 99 = 2
    16'b11101011_01100100 : OUT <= 2;  //235 / 100 = 2
    16'b11101011_01100101 : OUT <= 2;  //235 / 101 = 2
    16'b11101011_01100110 : OUT <= 2;  //235 / 102 = 2
    16'b11101011_01100111 : OUT <= 2;  //235 / 103 = 2
    16'b11101011_01101000 : OUT <= 2;  //235 / 104 = 2
    16'b11101011_01101001 : OUT <= 2;  //235 / 105 = 2
    16'b11101011_01101010 : OUT <= 2;  //235 / 106 = 2
    16'b11101011_01101011 : OUT <= 2;  //235 / 107 = 2
    16'b11101011_01101100 : OUT <= 2;  //235 / 108 = 2
    16'b11101011_01101101 : OUT <= 2;  //235 / 109 = 2
    16'b11101011_01101110 : OUT <= 2;  //235 / 110 = 2
    16'b11101011_01101111 : OUT <= 2;  //235 / 111 = 2
    16'b11101011_01110000 : OUT <= 2;  //235 / 112 = 2
    16'b11101011_01110001 : OUT <= 2;  //235 / 113 = 2
    16'b11101011_01110010 : OUT <= 2;  //235 / 114 = 2
    16'b11101011_01110011 : OUT <= 2;  //235 / 115 = 2
    16'b11101011_01110100 : OUT <= 2;  //235 / 116 = 2
    16'b11101011_01110101 : OUT <= 2;  //235 / 117 = 2
    16'b11101011_01110110 : OUT <= 1;  //235 / 118 = 1
    16'b11101011_01110111 : OUT <= 1;  //235 / 119 = 1
    16'b11101011_01111000 : OUT <= 1;  //235 / 120 = 1
    16'b11101011_01111001 : OUT <= 1;  //235 / 121 = 1
    16'b11101011_01111010 : OUT <= 1;  //235 / 122 = 1
    16'b11101011_01111011 : OUT <= 1;  //235 / 123 = 1
    16'b11101011_01111100 : OUT <= 1;  //235 / 124 = 1
    16'b11101011_01111101 : OUT <= 1;  //235 / 125 = 1
    16'b11101011_01111110 : OUT <= 1;  //235 / 126 = 1
    16'b11101011_01111111 : OUT <= 1;  //235 / 127 = 1
    16'b11101011_10000000 : OUT <= 1;  //235 / 128 = 1
    16'b11101011_10000001 : OUT <= 1;  //235 / 129 = 1
    16'b11101011_10000010 : OUT <= 1;  //235 / 130 = 1
    16'b11101011_10000011 : OUT <= 1;  //235 / 131 = 1
    16'b11101011_10000100 : OUT <= 1;  //235 / 132 = 1
    16'b11101011_10000101 : OUT <= 1;  //235 / 133 = 1
    16'b11101011_10000110 : OUT <= 1;  //235 / 134 = 1
    16'b11101011_10000111 : OUT <= 1;  //235 / 135 = 1
    16'b11101011_10001000 : OUT <= 1;  //235 / 136 = 1
    16'b11101011_10001001 : OUT <= 1;  //235 / 137 = 1
    16'b11101011_10001010 : OUT <= 1;  //235 / 138 = 1
    16'b11101011_10001011 : OUT <= 1;  //235 / 139 = 1
    16'b11101011_10001100 : OUT <= 1;  //235 / 140 = 1
    16'b11101011_10001101 : OUT <= 1;  //235 / 141 = 1
    16'b11101011_10001110 : OUT <= 1;  //235 / 142 = 1
    16'b11101011_10001111 : OUT <= 1;  //235 / 143 = 1
    16'b11101011_10010000 : OUT <= 1;  //235 / 144 = 1
    16'b11101011_10010001 : OUT <= 1;  //235 / 145 = 1
    16'b11101011_10010010 : OUT <= 1;  //235 / 146 = 1
    16'b11101011_10010011 : OUT <= 1;  //235 / 147 = 1
    16'b11101011_10010100 : OUT <= 1;  //235 / 148 = 1
    16'b11101011_10010101 : OUT <= 1;  //235 / 149 = 1
    16'b11101011_10010110 : OUT <= 1;  //235 / 150 = 1
    16'b11101011_10010111 : OUT <= 1;  //235 / 151 = 1
    16'b11101011_10011000 : OUT <= 1;  //235 / 152 = 1
    16'b11101011_10011001 : OUT <= 1;  //235 / 153 = 1
    16'b11101011_10011010 : OUT <= 1;  //235 / 154 = 1
    16'b11101011_10011011 : OUT <= 1;  //235 / 155 = 1
    16'b11101011_10011100 : OUT <= 1;  //235 / 156 = 1
    16'b11101011_10011101 : OUT <= 1;  //235 / 157 = 1
    16'b11101011_10011110 : OUT <= 1;  //235 / 158 = 1
    16'b11101011_10011111 : OUT <= 1;  //235 / 159 = 1
    16'b11101011_10100000 : OUT <= 1;  //235 / 160 = 1
    16'b11101011_10100001 : OUT <= 1;  //235 / 161 = 1
    16'b11101011_10100010 : OUT <= 1;  //235 / 162 = 1
    16'b11101011_10100011 : OUT <= 1;  //235 / 163 = 1
    16'b11101011_10100100 : OUT <= 1;  //235 / 164 = 1
    16'b11101011_10100101 : OUT <= 1;  //235 / 165 = 1
    16'b11101011_10100110 : OUT <= 1;  //235 / 166 = 1
    16'b11101011_10100111 : OUT <= 1;  //235 / 167 = 1
    16'b11101011_10101000 : OUT <= 1;  //235 / 168 = 1
    16'b11101011_10101001 : OUT <= 1;  //235 / 169 = 1
    16'b11101011_10101010 : OUT <= 1;  //235 / 170 = 1
    16'b11101011_10101011 : OUT <= 1;  //235 / 171 = 1
    16'b11101011_10101100 : OUT <= 1;  //235 / 172 = 1
    16'b11101011_10101101 : OUT <= 1;  //235 / 173 = 1
    16'b11101011_10101110 : OUT <= 1;  //235 / 174 = 1
    16'b11101011_10101111 : OUT <= 1;  //235 / 175 = 1
    16'b11101011_10110000 : OUT <= 1;  //235 / 176 = 1
    16'b11101011_10110001 : OUT <= 1;  //235 / 177 = 1
    16'b11101011_10110010 : OUT <= 1;  //235 / 178 = 1
    16'b11101011_10110011 : OUT <= 1;  //235 / 179 = 1
    16'b11101011_10110100 : OUT <= 1;  //235 / 180 = 1
    16'b11101011_10110101 : OUT <= 1;  //235 / 181 = 1
    16'b11101011_10110110 : OUT <= 1;  //235 / 182 = 1
    16'b11101011_10110111 : OUT <= 1;  //235 / 183 = 1
    16'b11101011_10111000 : OUT <= 1;  //235 / 184 = 1
    16'b11101011_10111001 : OUT <= 1;  //235 / 185 = 1
    16'b11101011_10111010 : OUT <= 1;  //235 / 186 = 1
    16'b11101011_10111011 : OUT <= 1;  //235 / 187 = 1
    16'b11101011_10111100 : OUT <= 1;  //235 / 188 = 1
    16'b11101011_10111101 : OUT <= 1;  //235 / 189 = 1
    16'b11101011_10111110 : OUT <= 1;  //235 / 190 = 1
    16'b11101011_10111111 : OUT <= 1;  //235 / 191 = 1
    16'b11101011_11000000 : OUT <= 1;  //235 / 192 = 1
    16'b11101011_11000001 : OUT <= 1;  //235 / 193 = 1
    16'b11101011_11000010 : OUT <= 1;  //235 / 194 = 1
    16'b11101011_11000011 : OUT <= 1;  //235 / 195 = 1
    16'b11101011_11000100 : OUT <= 1;  //235 / 196 = 1
    16'b11101011_11000101 : OUT <= 1;  //235 / 197 = 1
    16'b11101011_11000110 : OUT <= 1;  //235 / 198 = 1
    16'b11101011_11000111 : OUT <= 1;  //235 / 199 = 1
    16'b11101011_11001000 : OUT <= 1;  //235 / 200 = 1
    16'b11101011_11001001 : OUT <= 1;  //235 / 201 = 1
    16'b11101011_11001010 : OUT <= 1;  //235 / 202 = 1
    16'b11101011_11001011 : OUT <= 1;  //235 / 203 = 1
    16'b11101011_11001100 : OUT <= 1;  //235 / 204 = 1
    16'b11101011_11001101 : OUT <= 1;  //235 / 205 = 1
    16'b11101011_11001110 : OUT <= 1;  //235 / 206 = 1
    16'b11101011_11001111 : OUT <= 1;  //235 / 207 = 1
    16'b11101011_11010000 : OUT <= 1;  //235 / 208 = 1
    16'b11101011_11010001 : OUT <= 1;  //235 / 209 = 1
    16'b11101011_11010010 : OUT <= 1;  //235 / 210 = 1
    16'b11101011_11010011 : OUT <= 1;  //235 / 211 = 1
    16'b11101011_11010100 : OUT <= 1;  //235 / 212 = 1
    16'b11101011_11010101 : OUT <= 1;  //235 / 213 = 1
    16'b11101011_11010110 : OUT <= 1;  //235 / 214 = 1
    16'b11101011_11010111 : OUT <= 1;  //235 / 215 = 1
    16'b11101011_11011000 : OUT <= 1;  //235 / 216 = 1
    16'b11101011_11011001 : OUT <= 1;  //235 / 217 = 1
    16'b11101011_11011010 : OUT <= 1;  //235 / 218 = 1
    16'b11101011_11011011 : OUT <= 1;  //235 / 219 = 1
    16'b11101011_11011100 : OUT <= 1;  //235 / 220 = 1
    16'b11101011_11011101 : OUT <= 1;  //235 / 221 = 1
    16'b11101011_11011110 : OUT <= 1;  //235 / 222 = 1
    16'b11101011_11011111 : OUT <= 1;  //235 / 223 = 1
    16'b11101011_11100000 : OUT <= 1;  //235 / 224 = 1
    16'b11101011_11100001 : OUT <= 1;  //235 / 225 = 1
    16'b11101011_11100010 : OUT <= 1;  //235 / 226 = 1
    16'b11101011_11100011 : OUT <= 1;  //235 / 227 = 1
    16'b11101011_11100100 : OUT <= 1;  //235 / 228 = 1
    16'b11101011_11100101 : OUT <= 1;  //235 / 229 = 1
    16'b11101011_11100110 : OUT <= 1;  //235 / 230 = 1
    16'b11101011_11100111 : OUT <= 1;  //235 / 231 = 1
    16'b11101011_11101000 : OUT <= 1;  //235 / 232 = 1
    16'b11101011_11101001 : OUT <= 1;  //235 / 233 = 1
    16'b11101011_11101010 : OUT <= 1;  //235 / 234 = 1
    16'b11101011_11101011 : OUT <= 1;  //235 / 235 = 1
    16'b11101011_11101100 : OUT <= 0;  //235 / 236 = 0
    16'b11101011_11101101 : OUT <= 0;  //235 / 237 = 0
    16'b11101011_11101110 : OUT <= 0;  //235 / 238 = 0
    16'b11101011_11101111 : OUT <= 0;  //235 / 239 = 0
    16'b11101011_11110000 : OUT <= 0;  //235 / 240 = 0
    16'b11101011_11110001 : OUT <= 0;  //235 / 241 = 0
    16'b11101011_11110010 : OUT <= 0;  //235 / 242 = 0
    16'b11101011_11110011 : OUT <= 0;  //235 / 243 = 0
    16'b11101011_11110100 : OUT <= 0;  //235 / 244 = 0
    16'b11101011_11110101 : OUT <= 0;  //235 / 245 = 0
    16'b11101011_11110110 : OUT <= 0;  //235 / 246 = 0
    16'b11101011_11110111 : OUT <= 0;  //235 / 247 = 0
    16'b11101011_11111000 : OUT <= 0;  //235 / 248 = 0
    16'b11101011_11111001 : OUT <= 0;  //235 / 249 = 0
    16'b11101011_11111010 : OUT <= 0;  //235 / 250 = 0
    16'b11101011_11111011 : OUT <= 0;  //235 / 251 = 0
    16'b11101011_11111100 : OUT <= 0;  //235 / 252 = 0
    16'b11101011_11111101 : OUT <= 0;  //235 / 253 = 0
    16'b11101011_11111110 : OUT <= 0;  //235 / 254 = 0
    16'b11101011_11111111 : OUT <= 0;  //235 / 255 = 0
    16'b11101100_00000000 : OUT <= 0;  //236 / 0 = 0
    16'b11101100_00000001 : OUT <= 236;  //236 / 1 = 236
    16'b11101100_00000010 : OUT <= 118;  //236 / 2 = 118
    16'b11101100_00000011 : OUT <= 78;  //236 / 3 = 78
    16'b11101100_00000100 : OUT <= 59;  //236 / 4 = 59
    16'b11101100_00000101 : OUT <= 47;  //236 / 5 = 47
    16'b11101100_00000110 : OUT <= 39;  //236 / 6 = 39
    16'b11101100_00000111 : OUT <= 33;  //236 / 7 = 33
    16'b11101100_00001000 : OUT <= 29;  //236 / 8 = 29
    16'b11101100_00001001 : OUT <= 26;  //236 / 9 = 26
    16'b11101100_00001010 : OUT <= 23;  //236 / 10 = 23
    16'b11101100_00001011 : OUT <= 21;  //236 / 11 = 21
    16'b11101100_00001100 : OUT <= 19;  //236 / 12 = 19
    16'b11101100_00001101 : OUT <= 18;  //236 / 13 = 18
    16'b11101100_00001110 : OUT <= 16;  //236 / 14 = 16
    16'b11101100_00001111 : OUT <= 15;  //236 / 15 = 15
    16'b11101100_00010000 : OUT <= 14;  //236 / 16 = 14
    16'b11101100_00010001 : OUT <= 13;  //236 / 17 = 13
    16'b11101100_00010010 : OUT <= 13;  //236 / 18 = 13
    16'b11101100_00010011 : OUT <= 12;  //236 / 19 = 12
    16'b11101100_00010100 : OUT <= 11;  //236 / 20 = 11
    16'b11101100_00010101 : OUT <= 11;  //236 / 21 = 11
    16'b11101100_00010110 : OUT <= 10;  //236 / 22 = 10
    16'b11101100_00010111 : OUT <= 10;  //236 / 23 = 10
    16'b11101100_00011000 : OUT <= 9;  //236 / 24 = 9
    16'b11101100_00011001 : OUT <= 9;  //236 / 25 = 9
    16'b11101100_00011010 : OUT <= 9;  //236 / 26 = 9
    16'b11101100_00011011 : OUT <= 8;  //236 / 27 = 8
    16'b11101100_00011100 : OUT <= 8;  //236 / 28 = 8
    16'b11101100_00011101 : OUT <= 8;  //236 / 29 = 8
    16'b11101100_00011110 : OUT <= 7;  //236 / 30 = 7
    16'b11101100_00011111 : OUT <= 7;  //236 / 31 = 7
    16'b11101100_00100000 : OUT <= 7;  //236 / 32 = 7
    16'b11101100_00100001 : OUT <= 7;  //236 / 33 = 7
    16'b11101100_00100010 : OUT <= 6;  //236 / 34 = 6
    16'b11101100_00100011 : OUT <= 6;  //236 / 35 = 6
    16'b11101100_00100100 : OUT <= 6;  //236 / 36 = 6
    16'b11101100_00100101 : OUT <= 6;  //236 / 37 = 6
    16'b11101100_00100110 : OUT <= 6;  //236 / 38 = 6
    16'b11101100_00100111 : OUT <= 6;  //236 / 39 = 6
    16'b11101100_00101000 : OUT <= 5;  //236 / 40 = 5
    16'b11101100_00101001 : OUT <= 5;  //236 / 41 = 5
    16'b11101100_00101010 : OUT <= 5;  //236 / 42 = 5
    16'b11101100_00101011 : OUT <= 5;  //236 / 43 = 5
    16'b11101100_00101100 : OUT <= 5;  //236 / 44 = 5
    16'b11101100_00101101 : OUT <= 5;  //236 / 45 = 5
    16'b11101100_00101110 : OUT <= 5;  //236 / 46 = 5
    16'b11101100_00101111 : OUT <= 5;  //236 / 47 = 5
    16'b11101100_00110000 : OUT <= 4;  //236 / 48 = 4
    16'b11101100_00110001 : OUT <= 4;  //236 / 49 = 4
    16'b11101100_00110010 : OUT <= 4;  //236 / 50 = 4
    16'b11101100_00110011 : OUT <= 4;  //236 / 51 = 4
    16'b11101100_00110100 : OUT <= 4;  //236 / 52 = 4
    16'b11101100_00110101 : OUT <= 4;  //236 / 53 = 4
    16'b11101100_00110110 : OUT <= 4;  //236 / 54 = 4
    16'b11101100_00110111 : OUT <= 4;  //236 / 55 = 4
    16'b11101100_00111000 : OUT <= 4;  //236 / 56 = 4
    16'b11101100_00111001 : OUT <= 4;  //236 / 57 = 4
    16'b11101100_00111010 : OUT <= 4;  //236 / 58 = 4
    16'b11101100_00111011 : OUT <= 4;  //236 / 59 = 4
    16'b11101100_00111100 : OUT <= 3;  //236 / 60 = 3
    16'b11101100_00111101 : OUT <= 3;  //236 / 61 = 3
    16'b11101100_00111110 : OUT <= 3;  //236 / 62 = 3
    16'b11101100_00111111 : OUT <= 3;  //236 / 63 = 3
    16'b11101100_01000000 : OUT <= 3;  //236 / 64 = 3
    16'b11101100_01000001 : OUT <= 3;  //236 / 65 = 3
    16'b11101100_01000010 : OUT <= 3;  //236 / 66 = 3
    16'b11101100_01000011 : OUT <= 3;  //236 / 67 = 3
    16'b11101100_01000100 : OUT <= 3;  //236 / 68 = 3
    16'b11101100_01000101 : OUT <= 3;  //236 / 69 = 3
    16'b11101100_01000110 : OUT <= 3;  //236 / 70 = 3
    16'b11101100_01000111 : OUT <= 3;  //236 / 71 = 3
    16'b11101100_01001000 : OUT <= 3;  //236 / 72 = 3
    16'b11101100_01001001 : OUT <= 3;  //236 / 73 = 3
    16'b11101100_01001010 : OUT <= 3;  //236 / 74 = 3
    16'b11101100_01001011 : OUT <= 3;  //236 / 75 = 3
    16'b11101100_01001100 : OUT <= 3;  //236 / 76 = 3
    16'b11101100_01001101 : OUT <= 3;  //236 / 77 = 3
    16'b11101100_01001110 : OUT <= 3;  //236 / 78 = 3
    16'b11101100_01001111 : OUT <= 2;  //236 / 79 = 2
    16'b11101100_01010000 : OUT <= 2;  //236 / 80 = 2
    16'b11101100_01010001 : OUT <= 2;  //236 / 81 = 2
    16'b11101100_01010010 : OUT <= 2;  //236 / 82 = 2
    16'b11101100_01010011 : OUT <= 2;  //236 / 83 = 2
    16'b11101100_01010100 : OUT <= 2;  //236 / 84 = 2
    16'b11101100_01010101 : OUT <= 2;  //236 / 85 = 2
    16'b11101100_01010110 : OUT <= 2;  //236 / 86 = 2
    16'b11101100_01010111 : OUT <= 2;  //236 / 87 = 2
    16'b11101100_01011000 : OUT <= 2;  //236 / 88 = 2
    16'b11101100_01011001 : OUT <= 2;  //236 / 89 = 2
    16'b11101100_01011010 : OUT <= 2;  //236 / 90 = 2
    16'b11101100_01011011 : OUT <= 2;  //236 / 91 = 2
    16'b11101100_01011100 : OUT <= 2;  //236 / 92 = 2
    16'b11101100_01011101 : OUT <= 2;  //236 / 93 = 2
    16'b11101100_01011110 : OUT <= 2;  //236 / 94 = 2
    16'b11101100_01011111 : OUT <= 2;  //236 / 95 = 2
    16'b11101100_01100000 : OUT <= 2;  //236 / 96 = 2
    16'b11101100_01100001 : OUT <= 2;  //236 / 97 = 2
    16'b11101100_01100010 : OUT <= 2;  //236 / 98 = 2
    16'b11101100_01100011 : OUT <= 2;  //236 / 99 = 2
    16'b11101100_01100100 : OUT <= 2;  //236 / 100 = 2
    16'b11101100_01100101 : OUT <= 2;  //236 / 101 = 2
    16'b11101100_01100110 : OUT <= 2;  //236 / 102 = 2
    16'b11101100_01100111 : OUT <= 2;  //236 / 103 = 2
    16'b11101100_01101000 : OUT <= 2;  //236 / 104 = 2
    16'b11101100_01101001 : OUT <= 2;  //236 / 105 = 2
    16'b11101100_01101010 : OUT <= 2;  //236 / 106 = 2
    16'b11101100_01101011 : OUT <= 2;  //236 / 107 = 2
    16'b11101100_01101100 : OUT <= 2;  //236 / 108 = 2
    16'b11101100_01101101 : OUT <= 2;  //236 / 109 = 2
    16'b11101100_01101110 : OUT <= 2;  //236 / 110 = 2
    16'b11101100_01101111 : OUT <= 2;  //236 / 111 = 2
    16'b11101100_01110000 : OUT <= 2;  //236 / 112 = 2
    16'b11101100_01110001 : OUT <= 2;  //236 / 113 = 2
    16'b11101100_01110010 : OUT <= 2;  //236 / 114 = 2
    16'b11101100_01110011 : OUT <= 2;  //236 / 115 = 2
    16'b11101100_01110100 : OUT <= 2;  //236 / 116 = 2
    16'b11101100_01110101 : OUT <= 2;  //236 / 117 = 2
    16'b11101100_01110110 : OUT <= 2;  //236 / 118 = 2
    16'b11101100_01110111 : OUT <= 1;  //236 / 119 = 1
    16'b11101100_01111000 : OUT <= 1;  //236 / 120 = 1
    16'b11101100_01111001 : OUT <= 1;  //236 / 121 = 1
    16'b11101100_01111010 : OUT <= 1;  //236 / 122 = 1
    16'b11101100_01111011 : OUT <= 1;  //236 / 123 = 1
    16'b11101100_01111100 : OUT <= 1;  //236 / 124 = 1
    16'b11101100_01111101 : OUT <= 1;  //236 / 125 = 1
    16'b11101100_01111110 : OUT <= 1;  //236 / 126 = 1
    16'b11101100_01111111 : OUT <= 1;  //236 / 127 = 1
    16'b11101100_10000000 : OUT <= 1;  //236 / 128 = 1
    16'b11101100_10000001 : OUT <= 1;  //236 / 129 = 1
    16'b11101100_10000010 : OUT <= 1;  //236 / 130 = 1
    16'b11101100_10000011 : OUT <= 1;  //236 / 131 = 1
    16'b11101100_10000100 : OUT <= 1;  //236 / 132 = 1
    16'b11101100_10000101 : OUT <= 1;  //236 / 133 = 1
    16'b11101100_10000110 : OUT <= 1;  //236 / 134 = 1
    16'b11101100_10000111 : OUT <= 1;  //236 / 135 = 1
    16'b11101100_10001000 : OUT <= 1;  //236 / 136 = 1
    16'b11101100_10001001 : OUT <= 1;  //236 / 137 = 1
    16'b11101100_10001010 : OUT <= 1;  //236 / 138 = 1
    16'b11101100_10001011 : OUT <= 1;  //236 / 139 = 1
    16'b11101100_10001100 : OUT <= 1;  //236 / 140 = 1
    16'b11101100_10001101 : OUT <= 1;  //236 / 141 = 1
    16'b11101100_10001110 : OUT <= 1;  //236 / 142 = 1
    16'b11101100_10001111 : OUT <= 1;  //236 / 143 = 1
    16'b11101100_10010000 : OUT <= 1;  //236 / 144 = 1
    16'b11101100_10010001 : OUT <= 1;  //236 / 145 = 1
    16'b11101100_10010010 : OUT <= 1;  //236 / 146 = 1
    16'b11101100_10010011 : OUT <= 1;  //236 / 147 = 1
    16'b11101100_10010100 : OUT <= 1;  //236 / 148 = 1
    16'b11101100_10010101 : OUT <= 1;  //236 / 149 = 1
    16'b11101100_10010110 : OUT <= 1;  //236 / 150 = 1
    16'b11101100_10010111 : OUT <= 1;  //236 / 151 = 1
    16'b11101100_10011000 : OUT <= 1;  //236 / 152 = 1
    16'b11101100_10011001 : OUT <= 1;  //236 / 153 = 1
    16'b11101100_10011010 : OUT <= 1;  //236 / 154 = 1
    16'b11101100_10011011 : OUT <= 1;  //236 / 155 = 1
    16'b11101100_10011100 : OUT <= 1;  //236 / 156 = 1
    16'b11101100_10011101 : OUT <= 1;  //236 / 157 = 1
    16'b11101100_10011110 : OUT <= 1;  //236 / 158 = 1
    16'b11101100_10011111 : OUT <= 1;  //236 / 159 = 1
    16'b11101100_10100000 : OUT <= 1;  //236 / 160 = 1
    16'b11101100_10100001 : OUT <= 1;  //236 / 161 = 1
    16'b11101100_10100010 : OUT <= 1;  //236 / 162 = 1
    16'b11101100_10100011 : OUT <= 1;  //236 / 163 = 1
    16'b11101100_10100100 : OUT <= 1;  //236 / 164 = 1
    16'b11101100_10100101 : OUT <= 1;  //236 / 165 = 1
    16'b11101100_10100110 : OUT <= 1;  //236 / 166 = 1
    16'b11101100_10100111 : OUT <= 1;  //236 / 167 = 1
    16'b11101100_10101000 : OUT <= 1;  //236 / 168 = 1
    16'b11101100_10101001 : OUT <= 1;  //236 / 169 = 1
    16'b11101100_10101010 : OUT <= 1;  //236 / 170 = 1
    16'b11101100_10101011 : OUT <= 1;  //236 / 171 = 1
    16'b11101100_10101100 : OUT <= 1;  //236 / 172 = 1
    16'b11101100_10101101 : OUT <= 1;  //236 / 173 = 1
    16'b11101100_10101110 : OUT <= 1;  //236 / 174 = 1
    16'b11101100_10101111 : OUT <= 1;  //236 / 175 = 1
    16'b11101100_10110000 : OUT <= 1;  //236 / 176 = 1
    16'b11101100_10110001 : OUT <= 1;  //236 / 177 = 1
    16'b11101100_10110010 : OUT <= 1;  //236 / 178 = 1
    16'b11101100_10110011 : OUT <= 1;  //236 / 179 = 1
    16'b11101100_10110100 : OUT <= 1;  //236 / 180 = 1
    16'b11101100_10110101 : OUT <= 1;  //236 / 181 = 1
    16'b11101100_10110110 : OUT <= 1;  //236 / 182 = 1
    16'b11101100_10110111 : OUT <= 1;  //236 / 183 = 1
    16'b11101100_10111000 : OUT <= 1;  //236 / 184 = 1
    16'b11101100_10111001 : OUT <= 1;  //236 / 185 = 1
    16'b11101100_10111010 : OUT <= 1;  //236 / 186 = 1
    16'b11101100_10111011 : OUT <= 1;  //236 / 187 = 1
    16'b11101100_10111100 : OUT <= 1;  //236 / 188 = 1
    16'b11101100_10111101 : OUT <= 1;  //236 / 189 = 1
    16'b11101100_10111110 : OUT <= 1;  //236 / 190 = 1
    16'b11101100_10111111 : OUT <= 1;  //236 / 191 = 1
    16'b11101100_11000000 : OUT <= 1;  //236 / 192 = 1
    16'b11101100_11000001 : OUT <= 1;  //236 / 193 = 1
    16'b11101100_11000010 : OUT <= 1;  //236 / 194 = 1
    16'b11101100_11000011 : OUT <= 1;  //236 / 195 = 1
    16'b11101100_11000100 : OUT <= 1;  //236 / 196 = 1
    16'b11101100_11000101 : OUT <= 1;  //236 / 197 = 1
    16'b11101100_11000110 : OUT <= 1;  //236 / 198 = 1
    16'b11101100_11000111 : OUT <= 1;  //236 / 199 = 1
    16'b11101100_11001000 : OUT <= 1;  //236 / 200 = 1
    16'b11101100_11001001 : OUT <= 1;  //236 / 201 = 1
    16'b11101100_11001010 : OUT <= 1;  //236 / 202 = 1
    16'b11101100_11001011 : OUT <= 1;  //236 / 203 = 1
    16'b11101100_11001100 : OUT <= 1;  //236 / 204 = 1
    16'b11101100_11001101 : OUT <= 1;  //236 / 205 = 1
    16'b11101100_11001110 : OUT <= 1;  //236 / 206 = 1
    16'b11101100_11001111 : OUT <= 1;  //236 / 207 = 1
    16'b11101100_11010000 : OUT <= 1;  //236 / 208 = 1
    16'b11101100_11010001 : OUT <= 1;  //236 / 209 = 1
    16'b11101100_11010010 : OUT <= 1;  //236 / 210 = 1
    16'b11101100_11010011 : OUT <= 1;  //236 / 211 = 1
    16'b11101100_11010100 : OUT <= 1;  //236 / 212 = 1
    16'b11101100_11010101 : OUT <= 1;  //236 / 213 = 1
    16'b11101100_11010110 : OUT <= 1;  //236 / 214 = 1
    16'b11101100_11010111 : OUT <= 1;  //236 / 215 = 1
    16'b11101100_11011000 : OUT <= 1;  //236 / 216 = 1
    16'b11101100_11011001 : OUT <= 1;  //236 / 217 = 1
    16'b11101100_11011010 : OUT <= 1;  //236 / 218 = 1
    16'b11101100_11011011 : OUT <= 1;  //236 / 219 = 1
    16'b11101100_11011100 : OUT <= 1;  //236 / 220 = 1
    16'b11101100_11011101 : OUT <= 1;  //236 / 221 = 1
    16'b11101100_11011110 : OUT <= 1;  //236 / 222 = 1
    16'b11101100_11011111 : OUT <= 1;  //236 / 223 = 1
    16'b11101100_11100000 : OUT <= 1;  //236 / 224 = 1
    16'b11101100_11100001 : OUT <= 1;  //236 / 225 = 1
    16'b11101100_11100010 : OUT <= 1;  //236 / 226 = 1
    16'b11101100_11100011 : OUT <= 1;  //236 / 227 = 1
    16'b11101100_11100100 : OUT <= 1;  //236 / 228 = 1
    16'b11101100_11100101 : OUT <= 1;  //236 / 229 = 1
    16'b11101100_11100110 : OUT <= 1;  //236 / 230 = 1
    16'b11101100_11100111 : OUT <= 1;  //236 / 231 = 1
    16'b11101100_11101000 : OUT <= 1;  //236 / 232 = 1
    16'b11101100_11101001 : OUT <= 1;  //236 / 233 = 1
    16'b11101100_11101010 : OUT <= 1;  //236 / 234 = 1
    16'b11101100_11101011 : OUT <= 1;  //236 / 235 = 1
    16'b11101100_11101100 : OUT <= 1;  //236 / 236 = 1
    16'b11101100_11101101 : OUT <= 0;  //236 / 237 = 0
    16'b11101100_11101110 : OUT <= 0;  //236 / 238 = 0
    16'b11101100_11101111 : OUT <= 0;  //236 / 239 = 0
    16'b11101100_11110000 : OUT <= 0;  //236 / 240 = 0
    16'b11101100_11110001 : OUT <= 0;  //236 / 241 = 0
    16'b11101100_11110010 : OUT <= 0;  //236 / 242 = 0
    16'b11101100_11110011 : OUT <= 0;  //236 / 243 = 0
    16'b11101100_11110100 : OUT <= 0;  //236 / 244 = 0
    16'b11101100_11110101 : OUT <= 0;  //236 / 245 = 0
    16'b11101100_11110110 : OUT <= 0;  //236 / 246 = 0
    16'b11101100_11110111 : OUT <= 0;  //236 / 247 = 0
    16'b11101100_11111000 : OUT <= 0;  //236 / 248 = 0
    16'b11101100_11111001 : OUT <= 0;  //236 / 249 = 0
    16'b11101100_11111010 : OUT <= 0;  //236 / 250 = 0
    16'b11101100_11111011 : OUT <= 0;  //236 / 251 = 0
    16'b11101100_11111100 : OUT <= 0;  //236 / 252 = 0
    16'b11101100_11111101 : OUT <= 0;  //236 / 253 = 0
    16'b11101100_11111110 : OUT <= 0;  //236 / 254 = 0
    16'b11101100_11111111 : OUT <= 0;  //236 / 255 = 0
    16'b11101101_00000000 : OUT <= 0;  //237 / 0 = 0
    16'b11101101_00000001 : OUT <= 237;  //237 / 1 = 237
    16'b11101101_00000010 : OUT <= 118;  //237 / 2 = 118
    16'b11101101_00000011 : OUT <= 79;  //237 / 3 = 79
    16'b11101101_00000100 : OUT <= 59;  //237 / 4 = 59
    16'b11101101_00000101 : OUT <= 47;  //237 / 5 = 47
    16'b11101101_00000110 : OUT <= 39;  //237 / 6 = 39
    16'b11101101_00000111 : OUT <= 33;  //237 / 7 = 33
    16'b11101101_00001000 : OUT <= 29;  //237 / 8 = 29
    16'b11101101_00001001 : OUT <= 26;  //237 / 9 = 26
    16'b11101101_00001010 : OUT <= 23;  //237 / 10 = 23
    16'b11101101_00001011 : OUT <= 21;  //237 / 11 = 21
    16'b11101101_00001100 : OUT <= 19;  //237 / 12 = 19
    16'b11101101_00001101 : OUT <= 18;  //237 / 13 = 18
    16'b11101101_00001110 : OUT <= 16;  //237 / 14 = 16
    16'b11101101_00001111 : OUT <= 15;  //237 / 15 = 15
    16'b11101101_00010000 : OUT <= 14;  //237 / 16 = 14
    16'b11101101_00010001 : OUT <= 13;  //237 / 17 = 13
    16'b11101101_00010010 : OUT <= 13;  //237 / 18 = 13
    16'b11101101_00010011 : OUT <= 12;  //237 / 19 = 12
    16'b11101101_00010100 : OUT <= 11;  //237 / 20 = 11
    16'b11101101_00010101 : OUT <= 11;  //237 / 21 = 11
    16'b11101101_00010110 : OUT <= 10;  //237 / 22 = 10
    16'b11101101_00010111 : OUT <= 10;  //237 / 23 = 10
    16'b11101101_00011000 : OUT <= 9;  //237 / 24 = 9
    16'b11101101_00011001 : OUT <= 9;  //237 / 25 = 9
    16'b11101101_00011010 : OUT <= 9;  //237 / 26 = 9
    16'b11101101_00011011 : OUT <= 8;  //237 / 27 = 8
    16'b11101101_00011100 : OUT <= 8;  //237 / 28 = 8
    16'b11101101_00011101 : OUT <= 8;  //237 / 29 = 8
    16'b11101101_00011110 : OUT <= 7;  //237 / 30 = 7
    16'b11101101_00011111 : OUT <= 7;  //237 / 31 = 7
    16'b11101101_00100000 : OUT <= 7;  //237 / 32 = 7
    16'b11101101_00100001 : OUT <= 7;  //237 / 33 = 7
    16'b11101101_00100010 : OUT <= 6;  //237 / 34 = 6
    16'b11101101_00100011 : OUT <= 6;  //237 / 35 = 6
    16'b11101101_00100100 : OUT <= 6;  //237 / 36 = 6
    16'b11101101_00100101 : OUT <= 6;  //237 / 37 = 6
    16'b11101101_00100110 : OUT <= 6;  //237 / 38 = 6
    16'b11101101_00100111 : OUT <= 6;  //237 / 39 = 6
    16'b11101101_00101000 : OUT <= 5;  //237 / 40 = 5
    16'b11101101_00101001 : OUT <= 5;  //237 / 41 = 5
    16'b11101101_00101010 : OUT <= 5;  //237 / 42 = 5
    16'b11101101_00101011 : OUT <= 5;  //237 / 43 = 5
    16'b11101101_00101100 : OUT <= 5;  //237 / 44 = 5
    16'b11101101_00101101 : OUT <= 5;  //237 / 45 = 5
    16'b11101101_00101110 : OUT <= 5;  //237 / 46 = 5
    16'b11101101_00101111 : OUT <= 5;  //237 / 47 = 5
    16'b11101101_00110000 : OUT <= 4;  //237 / 48 = 4
    16'b11101101_00110001 : OUT <= 4;  //237 / 49 = 4
    16'b11101101_00110010 : OUT <= 4;  //237 / 50 = 4
    16'b11101101_00110011 : OUT <= 4;  //237 / 51 = 4
    16'b11101101_00110100 : OUT <= 4;  //237 / 52 = 4
    16'b11101101_00110101 : OUT <= 4;  //237 / 53 = 4
    16'b11101101_00110110 : OUT <= 4;  //237 / 54 = 4
    16'b11101101_00110111 : OUT <= 4;  //237 / 55 = 4
    16'b11101101_00111000 : OUT <= 4;  //237 / 56 = 4
    16'b11101101_00111001 : OUT <= 4;  //237 / 57 = 4
    16'b11101101_00111010 : OUT <= 4;  //237 / 58 = 4
    16'b11101101_00111011 : OUT <= 4;  //237 / 59 = 4
    16'b11101101_00111100 : OUT <= 3;  //237 / 60 = 3
    16'b11101101_00111101 : OUT <= 3;  //237 / 61 = 3
    16'b11101101_00111110 : OUT <= 3;  //237 / 62 = 3
    16'b11101101_00111111 : OUT <= 3;  //237 / 63 = 3
    16'b11101101_01000000 : OUT <= 3;  //237 / 64 = 3
    16'b11101101_01000001 : OUT <= 3;  //237 / 65 = 3
    16'b11101101_01000010 : OUT <= 3;  //237 / 66 = 3
    16'b11101101_01000011 : OUT <= 3;  //237 / 67 = 3
    16'b11101101_01000100 : OUT <= 3;  //237 / 68 = 3
    16'b11101101_01000101 : OUT <= 3;  //237 / 69 = 3
    16'b11101101_01000110 : OUT <= 3;  //237 / 70 = 3
    16'b11101101_01000111 : OUT <= 3;  //237 / 71 = 3
    16'b11101101_01001000 : OUT <= 3;  //237 / 72 = 3
    16'b11101101_01001001 : OUT <= 3;  //237 / 73 = 3
    16'b11101101_01001010 : OUT <= 3;  //237 / 74 = 3
    16'b11101101_01001011 : OUT <= 3;  //237 / 75 = 3
    16'b11101101_01001100 : OUT <= 3;  //237 / 76 = 3
    16'b11101101_01001101 : OUT <= 3;  //237 / 77 = 3
    16'b11101101_01001110 : OUT <= 3;  //237 / 78 = 3
    16'b11101101_01001111 : OUT <= 3;  //237 / 79 = 3
    16'b11101101_01010000 : OUT <= 2;  //237 / 80 = 2
    16'b11101101_01010001 : OUT <= 2;  //237 / 81 = 2
    16'b11101101_01010010 : OUT <= 2;  //237 / 82 = 2
    16'b11101101_01010011 : OUT <= 2;  //237 / 83 = 2
    16'b11101101_01010100 : OUT <= 2;  //237 / 84 = 2
    16'b11101101_01010101 : OUT <= 2;  //237 / 85 = 2
    16'b11101101_01010110 : OUT <= 2;  //237 / 86 = 2
    16'b11101101_01010111 : OUT <= 2;  //237 / 87 = 2
    16'b11101101_01011000 : OUT <= 2;  //237 / 88 = 2
    16'b11101101_01011001 : OUT <= 2;  //237 / 89 = 2
    16'b11101101_01011010 : OUT <= 2;  //237 / 90 = 2
    16'b11101101_01011011 : OUT <= 2;  //237 / 91 = 2
    16'b11101101_01011100 : OUT <= 2;  //237 / 92 = 2
    16'b11101101_01011101 : OUT <= 2;  //237 / 93 = 2
    16'b11101101_01011110 : OUT <= 2;  //237 / 94 = 2
    16'b11101101_01011111 : OUT <= 2;  //237 / 95 = 2
    16'b11101101_01100000 : OUT <= 2;  //237 / 96 = 2
    16'b11101101_01100001 : OUT <= 2;  //237 / 97 = 2
    16'b11101101_01100010 : OUT <= 2;  //237 / 98 = 2
    16'b11101101_01100011 : OUT <= 2;  //237 / 99 = 2
    16'b11101101_01100100 : OUT <= 2;  //237 / 100 = 2
    16'b11101101_01100101 : OUT <= 2;  //237 / 101 = 2
    16'b11101101_01100110 : OUT <= 2;  //237 / 102 = 2
    16'b11101101_01100111 : OUT <= 2;  //237 / 103 = 2
    16'b11101101_01101000 : OUT <= 2;  //237 / 104 = 2
    16'b11101101_01101001 : OUT <= 2;  //237 / 105 = 2
    16'b11101101_01101010 : OUT <= 2;  //237 / 106 = 2
    16'b11101101_01101011 : OUT <= 2;  //237 / 107 = 2
    16'b11101101_01101100 : OUT <= 2;  //237 / 108 = 2
    16'b11101101_01101101 : OUT <= 2;  //237 / 109 = 2
    16'b11101101_01101110 : OUT <= 2;  //237 / 110 = 2
    16'b11101101_01101111 : OUT <= 2;  //237 / 111 = 2
    16'b11101101_01110000 : OUT <= 2;  //237 / 112 = 2
    16'b11101101_01110001 : OUT <= 2;  //237 / 113 = 2
    16'b11101101_01110010 : OUT <= 2;  //237 / 114 = 2
    16'b11101101_01110011 : OUT <= 2;  //237 / 115 = 2
    16'b11101101_01110100 : OUT <= 2;  //237 / 116 = 2
    16'b11101101_01110101 : OUT <= 2;  //237 / 117 = 2
    16'b11101101_01110110 : OUT <= 2;  //237 / 118 = 2
    16'b11101101_01110111 : OUT <= 1;  //237 / 119 = 1
    16'b11101101_01111000 : OUT <= 1;  //237 / 120 = 1
    16'b11101101_01111001 : OUT <= 1;  //237 / 121 = 1
    16'b11101101_01111010 : OUT <= 1;  //237 / 122 = 1
    16'b11101101_01111011 : OUT <= 1;  //237 / 123 = 1
    16'b11101101_01111100 : OUT <= 1;  //237 / 124 = 1
    16'b11101101_01111101 : OUT <= 1;  //237 / 125 = 1
    16'b11101101_01111110 : OUT <= 1;  //237 / 126 = 1
    16'b11101101_01111111 : OUT <= 1;  //237 / 127 = 1
    16'b11101101_10000000 : OUT <= 1;  //237 / 128 = 1
    16'b11101101_10000001 : OUT <= 1;  //237 / 129 = 1
    16'b11101101_10000010 : OUT <= 1;  //237 / 130 = 1
    16'b11101101_10000011 : OUT <= 1;  //237 / 131 = 1
    16'b11101101_10000100 : OUT <= 1;  //237 / 132 = 1
    16'b11101101_10000101 : OUT <= 1;  //237 / 133 = 1
    16'b11101101_10000110 : OUT <= 1;  //237 / 134 = 1
    16'b11101101_10000111 : OUT <= 1;  //237 / 135 = 1
    16'b11101101_10001000 : OUT <= 1;  //237 / 136 = 1
    16'b11101101_10001001 : OUT <= 1;  //237 / 137 = 1
    16'b11101101_10001010 : OUT <= 1;  //237 / 138 = 1
    16'b11101101_10001011 : OUT <= 1;  //237 / 139 = 1
    16'b11101101_10001100 : OUT <= 1;  //237 / 140 = 1
    16'b11101101_10001101 : OUT <= 1;  //237 / 141 = 1
    16'b11101101_10001110 : OUT <= 1;  //237 / 142 = 1
    16'b11101101_10001111 : OUT <= 1;  //237 / 143 = 1
    16'b11101101_10010000 : OUT <= 1;  //237 / 144 = 1
    16'b11101101_10010001 : OUT <= 1;  //237 / 145 = 1
    16'b11101101_10010010 : OUT <= 1;  //237 / 146 = 1
    16'b11101101_10010011 : OUT <= 1;  //237 / 147 = 1
    16'b11101101_10010100 : OUT <= 1;  //237 / 148 = 1
    16'b11101101_10010101 : OUT <= 1;  //237 / 149 = 1
    16'b11101101_10010110 : OUT <= 1;  //237 / 150 = 1
    16'b11101101_10010111 : OUT <= 1;  //237 / 151 = 1
    16'b11101101_10011000 : OUT <= 1;  //237 / 152 = 1
    16'b11101101_10011001 : OUT <= 1;  //237 / 153 = 1
    16'b11101101_10011010 : OUT <= 1;  //237 / 154 = 1
    16'b11101101_10011011 : OUT <= 1;  //237 / 155 = 1
    16'b11101101_10011100 : OUT <= 1;  //237 / 156 = 1
    16'b11101101_10011101 : OUT <= 1;  //237 / 157 = 1
    16'b11101101_10011110 : OUT <= 1;  //237 / 158 = 1
    16'b11101101_10011111 : OUT <= 1;  //237 / 159 = 1
    16'b11101101_10100000 : OUT <= 1;  //237 / 160 = 1
    16'b11101101_10100001 : OUT <= 1;  //237 / 161 = 1
    16'b11101101_10100010 : OUT <= 1;  //237 / 162 = 1
    16'b11101101_10100011 : OUT <= 1;  //237 / 163 = 1
    16'b11101101_10100100 : OUT <= 1;  //237 / 164 = 1
    16'b11101101_10100101 : OUT <= 1;  //237 / 165 = 1
    16'b11101101_10100110 : OUT <= 1;  //237 / 166 = 1
    16'b11101101_10100111 : OUT <= 1;  //237 / 167 = 1
    16'b11101101_10101000 : OUT <= 1;  //237 / 168 = 1
    16'b11101101_10101001 : OUT <= 1;  //237 / 169 = 1
    16'b11101101_10101010 : OUT <= 1;  //237 / 170 = 1
    16'b11101101_10101011 : OUT <= 1;  //237 / 171 = 1
    16'b11101101_10101100 : OUT <= 1;  //237 / 172 = 1
    16'b11101101_10101101 : OUT <= 1;  //237 / 173 = 1
    16'b11101101_10101110 : OUT <= 1;  //237 / 174 = 1
    16'b11101101_10101111 : OUT <= 1;  //237 / 175 = 1
    16'b11101101_10110000 : OUT <= 1;  //237 / 176 = 1
    16'b11101101_10110001 : OUT <= 1;  //237 / 177 = 1
    16'b11101101_10110010 : OUT <= 1;  //237 / 178 = 1
    16'b11101101_10110011 : OUT <= 1;  //237 / 179 = 1
    16'b11101101_10110100 : OUT <= 1;  //237 / 180 = 1
    16'b11101101_10110101 : OUT <= 1;  //237 / 181 = 1
    16'b11101101_10110110 : OUT <= 1;  //237 / 182 = 1
    16'b11101101_10110111 : OUT <= 1;  //237 / 183 = 1
    16'b11101101_10111000 : OUT <= 1;  //237 / 184 = 1
    16'b11101101_10111001 : OUT <= 1;  //237 / 185 = 1
    16'b11101101_10111010 : OUT <= 1;  //237 / 186 = 1
    16'b11101101_10111011 : OUT <= 1;  //237 / 187 = 1
    16'b11101101_10111100 : OUT <= 1;  //237 / 188 = 1
    16'b11101101_10111101 : OUT <= 1;  //237 / 189 = 1
    16'b11101101_10111110 : OUT <= 1;  //237 / 190 = 1
    16'b11101101_10111111 : OUT <= 1;  //237 / 191 = 1
    16'b11101101_11000000 : OUT <= 1;  //237 / 192 = 1
    16'b11101101_11000001 : OUT <= 1;  //237 / 193 = 1
    16'b11101101_11000010 : OUT <= 1;  //237 / 194 = 1
    16'b11101101_11000011 : OUT <= 1;  //237 / 195 = 1
    16'b11101101_11000100 : OUT <= 1;  //237 / 196 = 1
    16'b11101101_11000101 : OUT <= 1;  //237 / 197 = 1
    16'b11101101_11000110 : OUT <= 1;  //237 / 198 = 1
    16'b11101101_11000111 : OUT <= 1;  //237 / 199 = 1
    16'b11101101_11001000 : OUT <= 1;  //237 / 200 = 1
    16'b11101101_11001001 : OUT <= 1;  //237 / 201 = 1
    16'b11101101_11001010 : OUT <= 1;  //237 / 202 = 1
    16'b11101101_11001011 : OUT <= 1;  //237 / 203 = 1
    16'b11101101_11001100 : OUT <= 1;  //237 / 204 = 1
    16'b11101101_11001101 : OUT <= 1;  //237 / 205 = 1
    16'b11101101_11001110 : OUT <= 1;  //237 / 206 = 1
    16'b11101101_11001111 : OUT <= 1;  //237 / 207 = 1
    16'b11101101_11010000 : OUT <= 1;  //237 / 208 = 1
    16'b11101101_11010001 : OUT <= 1;  //237 / 209 = 1
    16'b11101101_11010010 : OUT <= 1;  //237 / 210 = 1
    16'b11101101_11010011 : OUT <= 1;  //237 / 211 = 1
    16'b11101101_11010100 : OUT <= 1;  //237 / 212 = 1
    16'b11101101_11010101 : OUT <= 1;  //237 / 213 = 1
    16'b11101101_11010110 : OUT <= 1;  //237 / 214 = 1
    16'b11101101_11010111 : OUT <= 1;  //237 / 215 = 1
    16'b11101101_11011000 : OUT <= 1;  //237 / 216 = 1
    16'b11101101_11011001 : OUT <= 1;  //237 / 217 = 1
    16'b11101101_11011010 : OUT <= 1;  //237 / 218 = 1
    16'b11101101_11011011 : OUT <= 1;  //237 / 219 = 1
    16'b11101101_11011100 : OUT <= 1;  //237 / 220 = 1
    16'b11101101_11011101 : OUT <= 1;  //237 / 221 = 1
    16'b11101101_11011110 : OUT <= 1;  //237 / 222 = 1
    16'b11101101_11011111 : OUT <= 1;  //237 / 223 = 1
    16'b11101101_11100000 : OUT <= 1;  //237 / 224 = 1
    16'b11101101_11100001 : OUT <= 1;  //237 / 225 = 1
    16'b11101101_11100010 : OUT <= 1;  //237 / 226 = 1
    16'b11101101_11100011 : OUT <= 1;  //237 / 227 = 1
    16'b11101101_11100100 : OUT <= 1;  //237 / 228 = 1
    16'b11101101_11100101 : OUT <= 1;  //237 / 229 = 1
    16'b11101101_11100110 : OUT <= 1;  //237 / 230 = 1
    16'b11101101_11100111 : OUT <= 1;  //237 / 231 = 1
    16'b11101101_11101000 : OUT <= 1;  //237 / 232 = 1
    16'b11101101_11101001 : OUT <= 1;  //237 / 233 = 1
    16'b11101101_11101010 : OUT <= 1;  //237 / 234 = 1
    16'b11101101_11101011 : OUT <= 1;  //237 / 235 = 1
    16'b11101101_11101100 : OUT <= 1;  //237 / 236 = 1
    16'b11101101_11101101 : OUT <= 1;  //237 / 237 = 1
    16'b11101101_11101110 : OUT <= 0;  //237 / 238 = 0
    16'b11101101_11101111 : OUT <= 0;  //237 / 239 = 0
    16'b11101101_11110000 : OUT <= 0;  //237 / 240 = 0
    16'b11101101_11110001 : OUT <= 0;  //237 / 241 = 0
    16'b11101101_11110010 : OUT <= 0;  //237 / 242 = 0
    16'b11101101_11110011 : OUT <= 0;  //237 / 243 = 0
    16'b11101101_11110100 : OUT <= 0;  //237 / 244 = 0
    16'b11101101_11110101 : OUT <= 0;  //237 / 245 = 0
    16'b11101101_11110110 : OUT <= 0;  //237 / 246 = 0
    16'b11101101_11110111 : OUT <= 0;  //237 / 247 = 0
    16'b11101101_11111000 : OUT <= 0;  //237 / 248 = 0
    16'b11101101_11111001 : OUT <= 0;  //237 / 249 = 0
    16'b11101101_11111010 : OUT <= 0;  //237 / 250 = 0
    16'b11101101_11111011 : OUT <= 0;  //237 / 251 = 0
    16'b11101101_11111100 : OUT <= 0;  //237 / 252 = 0
    16'b11101101_11111101 : OUT <= 0;  //237 / 253 = 0
    16'b11101101_11111110 : OUT <= 0;  //237 / 254 = 0
    16'b11101101_11111111 : OUT <= 0;  //237 / 255 = 0
    16'b11101110_00000000 : OUT <= 0;  //238 / 0 = 0
    16'b11101110_00000001 : OUT <= 238;  //238 / 1 = 238
    16'b11101110_00000010 : OUT <= 119;  //238 / 2 = 119
    16'b11101110_00000011 : OUT <= 79;  //238 / 3 = 79
    16'b11101110_00000100 : OUT <= 59;  //238 / 4 = 59
    16'b11101110_00000101 : OUT <= 47;  //238 / 5 = 47
    16'b11101110_00000110 : OUT <= 39;  //238 / 6 = 39
    16'b11101110_00000111 : OUT <= 34;  //238 / 7 = 34
    16'b11101110_00001000 : OUT <= 29;  //238 / 8 = 29
    16'b11101110_00001001 : OUT <= 26;  //238 / 9 = 26
    16'b11101110_00001010 : OUT <= 23;  //238 / 10 = 23
    16'b11101110_00001011 : OUT <= 21;  //238 / 11 = 21
    16'b11101110_00001100 : OUT <= 19;  //238 / 12 = 19
    16'b11101110_00001101 : OUT <= 18;  //238 / 13 = 18
    16'b11101110_00001110 : OUT <= 17;  //238 / 14 = 17
    16'b11101110_00001111 : OUT <= 15;  //238 / 15 = 15
    16'b11101110_00010000 : OUT <= 14;  //238 / 16 = 14
    16'b11101110_00010001 : OUT <= 14;  //238 / 17 = 14
    16'b11101110_00010010 : OUT <= 13;  //238 / 18 = 13
    16'b11101110_00010011 : OUT <= 12;  //238 / 19 = 12
    16'b11101110_00010100 : OUT <= 11;  //238 / 20 = 11
    16'b11101110_00010101 : OUT <= 11;  //238 / 21 = 11
    16'b11101110_00010110 : OUT <= 10;  //238 / 22 = 10
    16'b11101110_00010111 : OUT <= 10;  //238 / 23 = 10
    16'b11101110_00011000 : OUT <= 9;  //238 / 24 = 9
    16'b11101110_00011001 : OUT <= 9;  //238 / 25 = 9
    16'b11101110_00011010 : OUT <= 9;  //238 / 26 = 9
    16'b11101110_00011011 : OUT <= 8;  //238 / 27 = 8
    16'b11101110_00011100 : OUT <= 8;  //238 / 28 = 8
    16'b11101110_00011101 : OUT <= 8;  //238 / 29 = 8
    16'b11101110_00011110 : OUT <= 7;  //238 / 30 = 7
    16'b11101110_00011111 : OUT <= 7;  //238 / 31 = 7
    16'b11101110_00100000 : OUT <= 7;  //238 / 32 = 7
    16'b11101110_00100001 : OUT <= 7;  //238 / 33 = 7
    16'b11101110_00100010 : OUT <= 7;  //238 / 34 = 7
    16'b11101110_00100011 : OUT <= 6;  //238 / 35 = 6
    16'b11101110_00100100 : OUT <= 6;  //238 / 36 = 6
    16'b11101110_00100101 : OUT <= 6;  //238 / 37 = 6
    16'b11101110_00100110 : OUT <= 6;  //238 / 38 = 6
    16'b11101110_00100111 : OUT <= 6;  //238 / 39 = 6
    16'b11101110_00101000 : OUT <= 5;  //238 / 40 = 5
    16'b11101110_00101001 : OUT <= 5;  //238 / 41 = 5
    16'b11101110_00101010 : OUT <= 5;  //238 / 42 = 5
    16'b11101110_00101011 : OUT <= 5;  //238 / 43 = 5
    16'b11101110_00101100 : OUT <= 5;  //238 / 44 = 5
    16'b11101110_00101101 : OUT <= 5;  //238 / 45 = 5
    16'b11101110_00101110 : OUT <= 5;  //238 / 46 = 5
    16'b11101110_00101111 : OUT <= 5;  //238 / 47 = 5
    16'b11101110_00110000 : OUT <= 4;  //238 / 48 = 4
    16'b11101110_00110001 : OUT <= 4;  //238 / 49 = 4
    16'b11101110_00110010 : OUT <= 4;  //238 / 50 = 4
    16'b11101110_00110011 : OUT <= 4;  //238 / 51 = 4
    16'b11101110_00110100 : OUT <= 4;  //238 / 52 = 4
    16'b11101110_00110101 : OUT <= 4;  //238 / 53 = 4
    16'b11101110_00110110 : OUT <= 4;  //238 / 54 = 4
    16'b11101110_00110111 : OUT <= 4;  //238 / 55 = 4
    16'b11101110_00111000 : OUT <= 4;  //238 / 56 = 4
    16'b11101110_00111001 : OUT <= 4;  //238 / 57 = 4
    16'b11101110_00111010 : OUT <= 4;  //238 / 58 = 4
    16'b11101110_00111011 : OUT <= 4;  //238 / 59 = 4
    16'b11101110_00111100 : OUT <= 3;  //238 / 60 = 3
    16'b11101110_00111101 : OUT <= 3;  //238 / 61 = 3
    16'b11101110_00111110 : OUT <= 3;  //238 / 62 = 3
    16'b11101110_00111111 : OUT <= 3;  //238 / 63 = 3
    16'b11101110_01000000 : OUT <= 3;  //238 / 64 = 3
    16'b11101110_01000001 : OUT <= 3;  //238 / 65 = 3
    16'b11101110_01000010 : OUT <= 3;  //238 / 66 = 3
    16'b11101110_01000011 : OUT <= 3;  //238 / 67 = 3
    16'b11101110_01000100 : OUT <= 3;  //238 / 68 = 3
    16'b11101110_01000101 : OUT <= 3;  //238 / 69 = 3
    16'b11101110_01000110 : OUT <= 3;  //238 / 70 = 3
    16'b11101110_01000111 : OUT <= 3;  //238 / 71 = 3
    16'b11101110_01001000 : OUT <= 3;  //238 / 72 = 3
    16'b11101110_01001001 : OUT <= 3;  //238 / 73 = 3
    16'b11101110_01001010 : OUT <= 3;  //238 / 74 = 3
    16'b11101110_01001011 : OUT <= 3;  //238 / 75 = 3
    16'b11101110_01001100 : OUT <= 3;  //238 / 76 = 3
    16'b11101110_01001101 : OUT <= 3;  //238 / 77 = 3
    16'b11101110_01001110 : OUT <= 3;  //238 / 78 = 3
    16'b11101110_01001111 : OUT <= 3;  //238 / 79 = 3
    16'b11101110_01010000 : OUT <= 2;  //238 / 80 = 2
    16'b11101110_01010001 : OUT <= 2;  //238 / 81 = 2
    16'b11101110_01010010 : OUT <= 2;  //238 / 82 = 2
    16'b11101110_01010011 : OUT <= 2;  //238 / 83 = 2
    16'b11101110_01010100 : OUT <= 2;  //238 / 84 = 2
    16'b11101110_01010101 : OUT <= 2;  //238 / 85 = 2
    16'b11101110_01010110 : OUT <= 2;  //238 / 86 = 2
    16'b11101110_01010111 : OUT <= 2;  //238 / 87 = 2
    16'b11101110_01011000 : OUT <= 2;  //238 / 88 = 2
    16'b11101110_01011001 : OUT <= 2;  //238 / 89 = 2
    16'b11101110_01011010 : OUT <= 2;  //238 / 90 = 2
    16'b11101110_01011011 : OUT <= 2;  //238 / 91 = 2
    16'b11101110_01011100 : OUT <= 2;  //238 / 92 = 2
    16'b11101110_01011101 : OUT <= 2;  //238 / 93 = 2
    16'b11101110_01011110 : OUT <= 2;  //238 / 94 = 2
    16'b11101110_01011111 : OUT <= 2;  //238 / 95 = 2
    16'b11101110_01100000 : OUT <= 2;  //238 / 96 = 2
    16'b11101110_01100001 : OUT <= 2;  //238 / 97 = 2
    16'b11101110_01100010 : OUT <= 2;  //238 / 98 = 2
    16'b11101110_01100011 : OUT <= 2;  //238 / 99 = 2
    16'b11101110_01100100 : OUT <= 2;  //238 / 100 = 2
    16'b11101110_01100101 : OUT <= 2;  //238 / 101 = 2
    16'b11101110_01100110 : OUT <= 2;  //238 / 102 = 2
    16'b11101110_01100111 : OUT <= 2;  //238 / 103 = 2
    16'b11101110_01101000 : OUT <= 2;  //238 / 104 = 2
    16'b11101110_01101001 : OUT <= 2;  //238 / 105 = 2
    16'b11101110_01101010 : OUT <= 2;  //238 / 106 = 2
    16'b11101110_01101011 : OUT <= 2;  //238 / 107 = 2
    16'b11101110_01101100 : OUT <= 2;  //238 / 108 = 2
    16'b11101110_01101101 : OUT <= 2;  //238 / 109 = 2
    16'b11101110_01101110 : OUT <= 2;  //238 / 110 = 2
    16'b11101110_01101111 : OUT <= 2;  //238 / 111 = 2
    16'b11101110_01110000 : OUT <= 2;  //238 / 112 = 2
    16'b11101110_01110001 : OUT <= 2;  //238 / 113 = 2
    16'b11101110_01110010 : OUT <= 2;  //238 / 114 = 2
    16'b11101110_01110011 : OUT <= 2;  //238 / 115 = 2
    16'b11101110_01110100 : OUT <= 2;  //238 / 116 = 2
    16'b11101110_01110101 : OUT <= 2;  //238 / 117 = 2
    16'b11101110_01110110 : OUT <= 2;  //238 / 118 = 2
    16'b11101110_01110111 : OUT <= 2;  //238 / 119 = 2
    16'b11101110_01111000 : OUT <= 1;  //238 / 120 = 1
    16'b11101110_01111001 : OUT <= 1;  //238 / 121 = 1
    16'b11101110_01111010 : OUT <= 1;  //238 / 122 = 1
    16'b11101110_01111011 : OUT <= 1;  //238 / 123 = 1
    16'b11101110_01111100 : OUT <= 1;  //238 / 124 = 1
    16'b11101110_01111101 : OUT <= 1;  //238 / 125 = 1
    16'b11101110_01111110 : OUT <= 1;  //238 / 126 = 1
    16'b11101110_01111111 : OUT <= 1;  //238 / 127 = 1
    16'b11101110_10000000 : OUT <= 1;  //238 / 128 = 1
    16'b11101110_10000001 : OUT <= 1;  //238 / 129 = 1
    16'b11101110_10000010 : OUT <= 1;  //238 / 130 = 1
    16'b11101110_10000011 : OUT <= 1;  //238 / 131 = 1
    16'b11101110_10000100 : OUT <= 1;  //238 / 132 = 1
    16'b11101110_10000101 : OUT <= 1;  //238 / 133 = 1
    16'b11101110_10000110 : OUT <= 1;  //238 / 134 = 1
    16'b11101110_10000111 : OUT <= 1;  //238 / 135 = 1
    16'b11101110_10001000 : OUT <= 1;  //238 / 136 = 1
    16'b11101110_10001001 : OUT <= 1;  //238 / 137 = 1
    16'b11101110_10001010 : OUT <= 1;  //238 / 138 = 1
    16'b11101110_10001011 : OUT <= 1;  //238 / 139 = 1
    16'b11101110_10001100 : OUT <= 1;  //238 / 140 = 1
    16'b11101110_10001101 : OUT <= 1;  //238 / 141 = 1
    16'b11101110_10001110 : OUT <= 1;  //238 / 142 = 1
    16'b11101110_10001111 : OUT <= 1;  //238 / 143 = 1
    16'b11101110_10010000 : OUT <= 1;  //238 / 144 = 1
    16'b11101110_10010001 : OUT <= 1;  //238 / 145 = 1
    16'b11101110_10010010 : OUT <= 1;  //238 / 146 = 1
    16'b11101110_10010011 : OUT <= 1;  //238 / 147 = 1
    16'b11101110_10010100 : OUT <= 1;  //238 / 148 = 1
    16'b11101110_10010101 : OUT <= 1;  //238 / 149 = 1
    16'b11101110_10010110 : OUT <= 1;  //238 / 150 = 1
    16'b11101110_10010111 : OUT <= 1;  //238 / 151 = 1
    16'b11101110_10011000 : OUT <= 1;  //238 / 152 = 1
    16'b11101110_10011001 : OUT <= 1;  //238 / 153 = 1
    16'b11101110_10011010 : OUT <= 1;  //238 / 154 = 1
    16'b11101110_10011011 : OUT <= 1;  //238 / 155 = 1
    16'b11101110_10011100 : OUT <= 1;  //238 / 156 = 1
    16'b11101110_10011101 : OUT <= 1;  //238 / 157 = 1
    16'b11101110_10011110 : OUT <= 1;  //238 / 158 = 1
    16'b11101110_10011111 : OUT <= 1;  //238 / 159 = 1
    16'b11101110_10100000 : OUT <= 1;  //238 / 160 = 1
    16'b11101110_10100001 : OUT <= 1;  //238 / 161 = 1
    16'b11101110_10100010 : OUT <= 1;  //238 / 162 = 1
    16'b11101110_10100011 : OUT <= 1;  //238 / 163 = 1
    16'b11101110_10100100 : OUT <= 1;  //238 / 164 = 1
    16'b11101110_10100101 : OUT <= 1;  //238 / 165 = 1
    16'b11101110_10100110 : OUT <= 1;  //238 / 166 = 1
    16'b11101110_10100111 : OUT <= 1;  //238 / 167 = 1
    16'b11101110_10101000 : OUT <= 1;  //238 / 168 = 1
    16'b11101110_10101001 : OUT <= 1;  //238 / 169 = 1
    16'b11101110_10101010 : OUT <= 1;  //238 / 170 = 1
    16'b11101110_10101011 : OUT <= 1;  //238 / 171 = 1
    16'b11101110_10101100 : OUT <= 1;  //238 / 172 = 1
    16'b11101110_10101101 : OUT <= 1;  //238 / 173 = 1
    16'b11101110_10101110 : OUT <= 1;  //238 / 174 = 1
    16'b11101110_10101111 : OUT <= 1;  //238 / 175 = 1
    16'b11101110_10110000 : OUT <= 1;  //238 / 176 = 1
    16'b11101110_10110001 : OUT <= 1;  //238 / 177 = 1
    16'b11101110_10110010 : OUT <= 1;  //238 / 178 = 1
    16'b11101110_10110011 : OUT <= 1;  //238 / 179 = 1
    16'b11101110_10110100 : OUT <= 1;  //238 / 180 = 1
    16'b11101110_10110101 : OUT <= 1;  //238 / 181 = 1
    16'b11101110_10110110 : OUT <= 1;  //238 / 182 = 1
    16'b11101110_10110111 : OUT <= 1;  //238 / 183 = 1
    16'b11101110_10111000 : OUT <= 1;  //238 / 184 = 1
    16'b11101110_10111001 : OUT <= 1;  //238 / 185 = 1
    16'b11101110_10111010 : OUT <= 1;  //238 / 186 = 1
    16'b11101110_10111011 : OUT <= 1;  //238 / 187 = 1
    16'b11101110_10111100 : OUT <= 1;  //238 / 188 = 1
    16'b11101110_10111101 : OUT <= 1;  //238 / 189 = 1
    16'b11101110_10111110 : OUT <= 1;  //238 / 190 = 1
    16'b11101110_10111111 : OUT <= 1;  //238 / 191 = 1
    16'b11101110_11000000 : OUT <= 1;  //238 / 192 = 1
    16'b11101110_11000001 : OUT <= 1;  //238 / 193 = 1
    16'b11101110_11000010 : OUT <= 1;  //238 / 194 = 1
    16'b11101110_11000011 : OUT <= 1;  //238 / 195 = 1
    16'b11101110_11000100 : OUT <= 1;  //238 / 196 = 1
    16'b11101110_11000101 : OUT <= 1;  //238 / 197 = 1
    16'b11101110_11000110 : OUT <= 1;  //238 / 198 = 1
    16'b11101110_11000111 : OUT <= 1;  //238 / 199 = 1
    16'b11101110_11001000 : OUT <= 1;  //238 / 200 = 1
    16'b11101110_11001001 : OUT <= 1;  //238 / 201 = 1
    16'b11101110_11001010 : OUT <= 1;  //238 / 202 = 1
    16'b11101110_11001011 : OUT <= 1;  //238 / 203 = 1
    16'b11101110_11001100 : OUT <= 1;  //238 / 204 = 1
    16'b11101110_11001101 : OUT <= 1;  //238 / 205 = 1
    16'b11101110_11001110 : OUT <= 1;  //238 / 206 = 1
    16'b11101110_11001111 : OUT <= 1;  //238 / 207 = 1
    16'b11101110_11010000 : OUT <= 1;  //238 / 208 = 1
    16'b11101110_11010001 : OUT <= 1;  //238 / 209 = 1
    16'b11101110_11010010 : OUT <= 1;  //238 / 210 = 1
    16'b11101110_11010011 : OUT <= 1;  //238 / 211 = 1
    16'b11101110_11010100 : OUT <= 1;  //238 / 212 = 1
    16'b11101110_11010101 : OUT <= 1;  //238 / 213 = 1
    16'b11101110_11010110 : OUT <= 1;  //238 / 214 = 1
    16'b11101110_11010111 : OUT <= 1;  //238 / 215 = 1
    16'b11101110_11011000 : OUT <= 1;  //238 / 216 = 1
    16'b11101110_11011001 : OUT <= 1;  //238 / 217 = 1
    16'b11101110_11011010 : OUT <= 1;  //238 / 218 = 1
    16'b11101110_11011011 : OUT <= 1;  //238 / 219 = 1
    16'b11101110_11011100 : OUT <= 1;  //238 / 220 = 1
    16'b11101110_11011101 : OUT <= 1;  //238 / 221 = 1
    16'b11101110_11011110 : OUT <= 1;  //238 / 222 = 1
    16'b11101110_11011111 : OUT <= 1;  //238 / 223 = 1
    16'b11101110_11100000 : OUT <= 1;  //238 / 224 = 1
    16'b11101110_11100001 : OUT <= 1;  //238 / 225 = 1
    16'b11101110_11100010 : OUT <= 1;  //238 / 226 = 1
    16'b11101110_11100011 : OUT <= 1;  //238 / 227 = 1
    16'b11101110_11100100 : OUT <= 1;  //238 / 228 = 1
    16'b11101110_11100101 : OUT <= 1;  //238 / 229 = 1
    16'b11101110_11100110 : OUT <= 1;  //238 / 230 = 1
    16'b11101110_11100111 : OUT <= 1;  //238 / 231 = 1
    16'b11101110_11101000 : OUT <= 1;  //238 / 232 = 1
    16'b11101110_11101001 : OUT <= 1;  //238 / 233 = 1
    16'b11101110_11101010 : OUT <= 1;  //238 / 234 = 1
    16'b11101110_11101011 : OUT <= 1;  //238 / 235 = 1
    16'b11101110_11101100 : OUT <= 1;  //238 / 236 = 1
    16'b11101110_11101101 : OUT <= 1;  //238 / 237 = 1
    16'b11101110_11101110 : OUT <= 1;  //238 / 238 = 1
    16'b11101110_11101111 : OUT <= 0;  //238 / 239 = 0
    16'b11101110_11110000 : OUT <= 0;  //238 / 240 = 0
    16'b11101110_11110001 : OUT <= 0;  //238 / 241 = 0
    16'b11101110_11110010 : OUT <= 0;  //238 / 242 = 0
    16'b11101110_11110011 : OUT <= 0;  //238 / 243 = 0
    16'b11101110_11110100 : OUT <= 0;  //238 / 244 = 0
    16'b11101110_11110101 : OUT <= 0;  //238 / 245 = 0
    16'b11101110_11110110 : OUT <= 0;  //238 / 246 = 0
    16'b11101110_11110111 : OUT <= 0;  //238 / 247 = 0
    16'b11101110_11111000 : OUT <= 0;  //238 / 248 = 0
    16'b11101110_11111001 : OUT <= 0;  //238 / 249 = 0
    16'b11101110_11111010 : OUT <= 0;  //238 / 250 = 0
    16'b11101110_11111011 : OUT <= 0;  //238 / 251 = 0
    16'b11101110_11111100 : OUT <= 0;  //238 / 252 = 0
    16'b11101110_11111101 : OUT <= 0;  //238 / 253 = 0
    16'b11101110_11111110 : OUT <= 0;  //238 / 254 = 0
    16'b11101110_11111111 : OUT <= 0;  //238 / 255 = 0
    16'b11101111_00000000 : OUT <= 0;  //239 / 0 = 0
    16'b11101111_00000001 : OUT <= 239;  //239 / 1 = 239
    16'b11101111_00000010 : OUT <= 119;  //239 / 2 = 119
    16'b11101111_00000011 : OUT <= 79;  //239 / 3 = 79
    16'b11101111_00000100 : OUT <= 59;  //239 / 4 = 59
    16'b11101111_00000101 : OUT <= 47;  //239 / 5 = 47
    16'b11101111_00000110 : OUT <= 39;  //239 / 6 = 39
    16'b11101111_00000111 : OUT <= 34;  //239 / 7 = 34
    16'b11101111_00001000 : OUT <= 29;  //239 / 8 = 29
    16'b11101111_00001001 : OUT <= 26;  //239 / 9 = 26
    16'b11101111_00001010 : OUT <= 23;  //239 / 10 = 23
    16'b11101111_00001011 : OUT <= 21;  //239 / 11 = 21
    16'b11101111_00001100 : OUT <= 19;  //239 / 12 = 19
    16'b11101111_00001101 : OUT <= 18;  //239 / 13 = 18
    16'b11101111_00001110 : OUT <= 17;  //239 / 14 = 17
    16'b11101111_00001111 : OUT <= 15;  //239 / 15 = 15
    16'b11101111_00010000 : OUT <= 14;  //239 / 16 = 14
    16'b11101111_00010001 : OUT <= 14;  //239 / 17 = 14
    16'b11101111_00010010 : OUT <= 13;  //239 / 18 = 13
    16'b11101111_00010011 : OUT <= 12;  //239 / 19 = 12
    16'b11101111_00010100 : OUT <= 11;  //239 / 20 = 11
    16'b11101111_00010101 : OUT <= 11;  //239 / 21 = 11
    16'b11101111_00010110 : OUT <= 10;  //239 / 22 = 10
    16'b11101111_00010111 : OUT <= 10;  //239 / 23 = 10
    16'b11101111_00011000 : OUT <= 9;  //239 / 24 = 9
    16'b11101111_00011001 : OUT <= 9;  //239 / 25 = 9
    16'b11101111_00011010 : OUT <= 9;  //239 / 26 = 9
    16'b11101111_00011011 : OUT <= 8;  //239 / 27 = 8
    16'b11101111_00011100 : OUT <= 8;  //239 / 28 = 8
    16'b11101111_00011101 : OUT <= 8;  //239 / 29 = 8
    16'b11101111_00011110 : OUT <= 7;  //239 / 30 = 7
    16'b11101111_00011111 : OUT <= 7;  //239 / 31 = 7
    16'b11101111_00100000 : OUT <= 7;  //239 / 32 = 7
    16'b11101111_00100001 : OUT <= 7;  //239 / 33 = 7
    16'b11101111_00100010 : OUT <= 7;  //239 / 34 = 7
    16'b11101111_00100011 : OUT <= 6;  //239 / 35 = 6
    16'b11101111_00100100 : OUT <= 6;  //239 / 36 = 6
    16'b11101111_00100101 : OUT <= 6;  //239 / 37 = 6
    16'b11101111_00100110 : OUT <= 6;  //239 / 38 = 6
    16'b11101111_00100111 : OUT <= 6;  //239 / 39 = 6
    16'b11101111_00101000 : OUT <= 5;  //239 / 40 = 5
    16'b11101111_00101001 : OUT <= 5;  //239 / 41 = 5
    16'b11101111_00101010 : OUT <= 5;  //239 / 42 = 5
    16'b11101111_00101011 : OUT <= 5;  //239 / 43 = 5
    16'b11101111_00101100 : OUT <= 5;  //239 / 44 = 5
    16'b11101111_00101101 : OUT <= 5;  //239 / 45 = 5
    16'b11101111_00101110 : OUT <= 5;  //239 / 46 = 5
    16'b11101111_00101111 : OUT <= 5;  //239 / 47 = 5
    16'b11101111_00110000 : OUT <= 4;  //239 / 48 = 4
    16'b11101111_00110001 : OUT <= 4;  //239 / 49 = 4
    16'b11101111_00110010 : OUT <= 4;  //239 / 50 = 4
    16'b11101111_00110011 : OUT <= 4;  //239 / 51 = 4
    16'b11101111_00110100 : OUT <= 4;  //239 / 52 = 4
    16'b11101111_00110101 : OUT <= 4;  //239 / 53 = 4
    16'b11101111_00110110 : OUT <= 4;  //239 / 54 = 4
    16'b11101111_00110111 : OUT <= 4;  //239 / 55 = 4
    16'b11101111_00111000 : OUT <= 4;  //239 / 56 = 4
    16'b11101111_00111001 : OUT <= 4;  //239 / 57 = 4
    16'b11101111_00111010 : OUT <= 4;  //239 / 58 = 4
    16'b11101111_00111011 : OUT <= 4;  //239 / 59 = 4
    16'b11101111_00111100 : OUT <= 3;  //239 / 60 = 3
    16'b11101111_00111101 : OUT <= 3;  //239 / 61 = 3
    16'b11101111_00111110 : OUT <= 3;  //239 / 62 = 3
    16'b11101111_00111111 : OUT <= 3;  //239 / 63 = 3
    16'b11101111_01000000 : OUT <= 3;  //239 / 64 = 3
    16'b11101111_01000001 : OUT <= 3;  //239 / 65 = 3
    16'b11101111_01000010 : OUT <= 3;  //239 / 66 = 3
    16'b11101111_01000011 : OUT <= 3;  //239 / 67 = 3
    16'b11101111_01000100 : OUT <= 3;  //239 / 68 = 3
    16'b11101111_01000101 : OUT <= 3;  //239 / 69 = 3
    16'b11101111_01000110 : OUT <= 3;  //239 / 70 = 3
    16'b11101111_01000111 : OUT <= 3;  //239 / 71 = 3
    16'b11101111_01001000 : OUT <= 3;  //239 / 72 = 3
    16'b11101111_01001001 : OUT <= 3;  //239 / 73 = 3
    16'b11101111_01001010 : OUT <= 3;  //239 / 74 = 3
    16'b11101111_01001011 : OUT <= 3;  //239 / 75 = 3
    16'b11101111_01001100 : OUT <= 3;  //239 / 76 = 3
    16'b11101111_01001101 : OUT <= 3;  //239 / 77 = 3
    16'b11101111_01001110 : OUT <= 3;  //239 / 78 = 3
    16'b11101111_01001111 : OUT <= 3;  //239 / 79 = 3
    16'b11101111_01010000 : OUT <= 2;  //239 / 80 = 2
    16'b11101111_01010001 : OUT <= 2;  //239 / 81 = 2
    16'b11101111_01010010 : OUT <= 2;  //239 / 82 = 2
    16'b11101111_01010011 : OUT <= 2;  //239 / 83 = 2
    16'b11101111_01010100 : OUT <= 2;  //239 / 84 = 2
    16'b11101111_01010101 : OUT <= 2;  //239 / 85 = 2
    16'b11101111_01010110 : OUT <= 2;  //239 / 86 = 2
    16'b11101111_01010111 : OUT <= 2;  //239 / 87 = 2
    16'b11101111_01011000 : OUT <= 2;  //239 / 88 = 2
    16'b11101111_01011001 : OUT <= 2;  //239 / 89 = 2
    16'b11101111_01011010 : OUT <= 2;  //239 / 90 = 2
    16'b11101111_01011011 : OUT <= 2;  //239 / 91 = 2
    16'b11101111_01011100 : OUT <= 2;  //239 / 92 = 2
    16'b11101111_01011101 : OUT <= 2;  //239 / 93 = 2
    16'b11101111_01011110 : OUT <= 2;  //239 / 94 = 2
    16'b11101111_01011111 : OUT <= 2;  //239 / 95 = 2
    16'b11101111_01100000 : OUT <= 2;  //239 / 96 = 2
    16'b11101111_01100001 : OUT <= 2;  //239 / 97 = 2
    16'b11101111_01100010 : OUT <= 2;  //239 / 98 = 2
    16'b11101111_01100011 : OUT <= 2;  //239 / 99 = 2
    16'b11101111_01100100 : OUT <= 2;  //239 / 100 = 2
    16'b11101111_01100101 : OUT <= 2;  //239 / 101 = 2
    16'b11101111_01100110 : OUT <= 2;  //239 / 102 = 2
    16'b11101111_01100111 : OUT <= 2;  //239 / 103 = 2
    16'b11101111_01101000 : OUT <= 2;  //239 / 104 = 2
    16'b11101111_01101001 : OUT <= 2;  //239 / 105 = 2
    16'b11101111_01101010 : OUT <= 2;  //239 / 106 = 2
    16'b11101111_01101011 : OUT <= 2;  //239 / 107 = 2
    16'b11101111_01101100 : OUT <= 2;  //239 / 108 = 2
    16'b11101111_01101101 : OUT <= 2;  //239 / 109 = 2
    16'b11101111_01101110 : OUT <= 2;  //239 / 110 = 2
    16'b11101111_01101111 : OUT <= 2;  //239 / 111 = 2
    16'b11101111_01110000 : OUT <= 2;  //239 / 112 = 2
    16'b11101111_01110001 : OUT <= 2;  //239 / 113 = 2
    16'b11101111_01110010 : OUT <= 2;  //239 / 114 = 2
    16'b11101111_01110011 : OUT <= 2;  //239 / 115 = 2
    16'b11101111_01110100 : OUT <= 2;  //239 / 116 = 2
    16'b11101111_01110101 : OUT <= 2;  //239 / 117 = 2
    16'b11101111_01110110 : OUT <= 2;  //239 / 118 = 2
    16'b11101111_01110111 : OUT <= 2;  //239 / 119 = 2
    16'b11101111_01111000 : OUT <= 1;  //239 / 120 = 1
    16'b11101111_01111001 : OUT <= 1;  //239 / 121 = 1
    16'b11101111_01111010 : OUT <= 1;  //239 / 122 = 1
    16'b11101111_01111011 : OUT <= 1;  //239 / 123 = 1
    16'b11101111_01111100 : OUT <= 1;  //239 / 124 = 1
    16'b11101111_01111101 : OUT <= 1;  //239 / 125 = 1
    16'b11101111_01111110 : OUT <= 1;  //239 / 126 = 1
    16'b11101111_01111111 : OUT <= 1;  //239 / 127 = 1
    16'b11101111_10000000 : OUT <= 1;  //239 / 128 = 1
    16'b11101111_10000001 : OUT <= 1;  //239 / 129 = 1
    16'b11101111_10000010 : OUT <= 1;  //239 / 130 = 1
    16'b11101111_10000011 : OUT <= 1;  //239 / 131 = 1
    16'b11101111_10000100 : OUT <= 1;  //239 / 132 = 1
    16'b11101111_10000101 : OUT <= 1;  //239 / 133 = 1
    16'b11101111_10000110 : OUT <= 1;  //239 / 134 = 1
    16'b11101111_10000111 : OUT <= 1;  //239 / 135 = 1
    16'b11101111_10001000 : OUT <= 1;  //239 / 136 = 1
    16'b11101111_10001001 : OUT <= 1;  //239 / 137 = 1
    16'b11101111_10001010 : OUT <= 1;  //239 / 138 = 1
    16'b11101111_10001011 : OUT <= 1;  //239 / 139 = 1
    16'b11101111_10001100 : OUT <= 1;  //239 / 140 = 1
    16'b11101111_10001101 : OUT <= 1;  //239 / 141 = 1
    16'b11101111_10001110 : OUT <= 1;  //239 / 142 = 1
    16'b11101111_10001111 : OUT <= 1;  //239 / 143 = 1
    16'b11101111_10010000 : OUT <= 1;  //239 / 144 = 1
    16'b11101111_10010001 : OUT <= 1;  //239 / 145 = 1
    16'b11101111_10010010 : OUT <= 1;  //239 / 146 = 1
    16'b11101111_10010011 : OUT <= 1;  //239 / 147 = 1
    16'b11101111_10010100 : OUT <= 1;  //239 / 148 = 1
    16'b11101111_10010101 : OUT <= 1;  //239 / 149 = 1
    16'b11101111_10010110 : OUT <= 1;  //239 / 150 = 1
    16'b11101111_10010111 : OUT <= 1;  //239 / 151 = 1
    16'b11101111_10011000 : OUT <= 1;  //239 / 152 = 1
    16'b11101111_10011001 : OUT <= 1;  //239 / 153 = 1
    16'b11101111_10011010 : OUT <= 1;  //239 / 154 = 1
    16'b11101111_10011011 : OUT <= 1;  //239 / 155 = 1
    16'b11101111_10011100 : OUT <= 1;  //239 / 156 = 1
    16'b11101111_10011101 : OUT <= 1;  //239 / 157 = 1
    16'b11101111_10011110 : OUT <= 1;  //239 / 158 = 1
    16'b11101111_10011111 : OUT <= 1;  //239 / 159 = 1
    16'b11101111_10100000 : OUT <= 1;  //239 / 160 = 1
    16'b11101111_10100001 : OUT <= 1;  //239 / 161 = 1
    16'b11101111_10100010 : OUT <= 1;  //239 / 162 = 1
    16'b11101111_10100011 : OUT <= 1;  //239 / 163 = 1
    16'b11101111_10100100 : OUT <= 1;  //239 / 164 = 1
    16'b11101111_10100101 : OUT <= 1;  //239 / 165 = 1
    16'b11101111_10100110 : OUT <= 1;  //239 / 166 = 1
    16'b11101111_10100111 : OUT <= 1;  //239 / 167 = 1
    16'b11101111_10101000 : OUT <= 1;  //239 / 168 = 1
    16'b11101111_10101001 : OUT <= 1;  //239 / 169 = 1
    16'b11101111_10101010 : OUT <= 1;  //239 / 170 = 1
    16'b11101111_10101011 : OUT <= 1;  //239 / 171 = 1
    16'b11101111_10101100 : OUT <= 1;  //239 / 172 = 1
    16'b11101111_10101101 : OUT <= 1;  //239 / 173 = 1
    16'b11101111_10101110 : OUT <= 1;  //239 / 174 = 1
    16'b11101111_10101111 : OUT <= 1;  //239 / 175 = 1
    16'b11101111_10110000 : OUT <= 1;  //239 / 176 = 1
    16'b11101111_10110001 : OUT <= 1;  //239 / 177 = 1
    16'b11101111_10110010 : OUT <= 1;  //239 / 178 = 1
    16'b11101111_10110011 : OUT <= 1;  //239 / 179 = 1
    16'b11101111_10110100 : OUT <= 1;  //239 / 180 = 1
    16'b11101111_10110101 : OUT <= 1;  //239 / 181 = 1
    16'b11101111_10110110 : OUT <= 1;  //239 / 182 = 1
    16'b11101111_10110111 : OUT <= 1;  //239 / 183 = 1
    16'b11101111_10111000 : OUT <= 1;  //239 / 184 = 1
    16'b11101111_10111001 : OUT <= 1;  //239 / 185 = 1
    16'b11101111_10111010 : OUT <= 1;  //239 / 186 = 1
    16'b11101111_10111011 : OUT <= 1;  //239 / 187 = 1
    16'b11101111_10111100 : OUT <= 1;  //239 / 188 = 1
    16'b11101111_10111101 : OUT <= 1;  //239 / 189 = 1
    16'b11101111_10111110 : OUT <= 1;  //239 / 190 = 1
    16'b11101111_10111111 : OUT <= 1;  //239 / 191 = 1
    16'b11101111_11000000 : OUT <= 1;  //239 / 192 = 1
    16'b11101111_11000001 : OUT <= 1;  //239 / 193 = 1
    16'b11101111_11000010 : OUT <= 1;  //239 / 194 = 1
    16'b11101111_11000011 : OUT <= 1;  //239 / 195 = 1
    16'b11101111_11000100 : OUT <= 1;  //239 / 196 = 1
    16'b11101111_11000101 : OUT <= 1;  //239 / 197 = 1
    16'b11101111_11000110 : OUT <= 1;  //239 / 198 = 1
    16'b11101111_11000111 : OUT <= 1;  //239 / 199 = 1
    16'b11101111_11001000 : OUT <= 1;  //239 / 200 = 1
    16'b11101111_11001001 : OUT <= 1;  //239 / 201 = 1
    16'b11101111_11001010 : OUT <= 1;  //239 / 202 = 1
    16'b11101111_11001011 : OUT <= 1;  //239 / 203 = 1
    16'b11101111_11001100 : OUT <= 1;  //239 / 204 = 1
    16'b11101111_11001101 : OUT <= 1;  //239 / 205 = 1
    16'b11101111_11001110 : OUT <= 1;  //239 / 206 = 1
    16'b11101111_11001111 : OUT <= 1;  //239 / 207 = 1
    16'b11101111_11010000 : OUT <= 1;  //239 / 208 = 1
    16'b11101111_11010001 : OUT <= 1;  //239 / 209 = 1
    16'b11101111_11010010 : OUT <= 1;  //239 / 210 = 1
    16'b11101111_11010011 : OUT <= 1;  //239 / 211 = 1
    16'b11101111_11010100 : OUT <= 1;  //239 / 212 = 1
    16'b11101111_11010101 : OUT <= 1;  //239 / 213 = 1
    16'b11101111_11010110 : OUT <= 1;  //239 / 214 = 1
    16'b11101111_11010111 : OUT <= 1;  //239 / 215 = 1
    16'b11101111_11011000 : OUT <= 1;  //239 / 216 = 1
    16'b11101111_11011001 : OUT <= 1;  //239 / 217 = 1
    16'b11101111_11011010 : OUT <= 1;  //239 / 218 = 1
    16'b11101111_11011011 : OUT <= 1;  //239 / 219 = 1
    16'b11101111_11011100 : OUT <= 1;  //239 / 220 = 1
    16'b11101111_11011101 : OUT <= 1;  //239 / 221 = 1
    16'b11101111_11011110 : OUT <= 1;  //239 / 222 = 1
    16'b11101111_11011111 : OUT <= 1;  //239 / 223 = 1
    16'b11101111_11100000 : OUT <= 1;  //239 / 224 = 1
    16'b11101111_11100001 : OUT <= 1;  //239 / 225 = 1
    16'b11101111_11100010 : OUT <= 1;  //239 / 226 = 1
    16'b11101111_11100011 : OUT <= 1;  //239 / 227 = 1
    16'b11101111_11100100 : OUT <= 1;  //239 / 228 = 1
    16'b11101111_11100101 : OUT <= 1;  //239 / 229 = 1
    16'b11101111_11100110 : OUT <= 1;  //239 / 230 = 1
    16'b11101111_11100111 : OUT <= 1;  //239 / 231 = 1
    16'b11101111_11101000 : OUT <= 1;  //239 / 232 = 1
    16'b11101111_11101001 : OUT <= 1;  //239 / 233 = 1
    16'b11101111_11101010 : OUT <= 1;  //239 / 234 = 1
    16'b11101111_11101011 : OUT <= 1;  //239 / 235 = 1
    16'b11101111_11101100 : OUT <= 1;  //239 / 236 = 1
    16'b11101111_11101101 : OUT <= 1;  //239 / 237 = 1
    16'b11101111_11101110 : OUT <= 1;  //239 / 238 = 1
    16'b11101111_11101111 : OUT <= 1;  //239 / 239 = 1
    16'b11101111_11110000 : OUT <= 0;  //239 / 240 = 0
    16'b11101111_11110001 : OUT <= 0;  //239 / 241 = 0
    16'b11101111_11110010 : OUT <= 0;  //239 / 242 = 0
    16'b11101111_11110011 : OUT <= 0;  //239 / 243 = 0
    16'b11101111_11110100 : OUT <= 0;  //239 / 244 = 0
    16'b11101111_11110101 : OUT <= 0;  //239 / 245 = 0
    16'b11101111_11110110 : OUT <= 0;  //239 / 246 = 0
    16'b11101111_11110111 : OUT <= 0;  //239 / 247 = 0
    16'b11101111_11111000 : OUT <= 0;  //239 / 248 = 0
    16'b11101111_11111001 : OUT <= 0;  //239 / 249 = 0
    16'b11101111_11111010 : OUT <= 0;  //239 / 250 = 0
    16'b11101111_11111011 : OUT <= 0;  //239 / 251 = 0
    16'b11101111_11111100 : OUT <= 0;  //239 / 252 = 0
    16'b11101111_11111101 : OUT <= 0;  //239 / 253 = 0
    16'b11101111_11111110 : OUT <= 0;  //239 / 254 = 0
    16'b11101111_11111111 : OUT <= 0;  //239 / 255 = 0
    16'b11110000_00000000 : OUT <= 0;  //240 / 0 = 0
    16'b11110000_00000001 : OUT <= 240;  //240 / 1 = 240
    16'b11110000_00000010 : OUT <= 120;  //240 / 2 = 120
    16'b11110000_00000011 : OUT <= 80;  //240 / 3 = 80
    16'b11110000_00000100 : OUT <= 60;  //240 / 4 = 60
    16'b11110000_00000101 : OUT <= 48;  //240 / 5 = 48
    16'b11110000_00000110 : OUT <= 40;  //240 / 6 = 40
    16'b11110000_00000111 : OUT <= 34;  //240 / 7 = 34
    16'b11110000_00001000 : OUT <= 30;  //240 / 8 = 30
    16'b11110000_00001001 : OUT <= 26;  //240 / 9 = 26
    16'b11110000_00001010 : OUT <= 24;  //240 / 10 = 24
    16'b11110000_00001011 : OUT <= 21;  //240 / 11 = 21
    16'b11110000_00001100 : OUT <= 20;  //240 / 12 = 20
    16'b11110000_00001101 : OUT <= 18;  //240 / 13 = 18
    16'b11110000_00001110 : OUT <= 17;  //240 / 14 = 17
    16'b11110000_00001111 : OUT <= 16;  //240 / 15 = 16
    16'b11110000_00010000 : OUT <= 15;  //240 / 16 = 15
    16'b11110000_00010001 : OUT <= 14;  //240 / 17 = 14
    16'b11110000_00010010 : OUT <= 13;  //240 / 18 = 13
    16'b11110000_00010011 : OUT <= 12;  //240 / 19 = 12
    16'b11110000_00010100 : OUT <= 12;  //240 / 20 = 12
    16'b11110000_00010101 : OUT <= 11;  //240 / 21 = 11
    16'b11110000_00010110 : OUT <= 10;  //240 / 22 = 10
    16'b11110000_00010111 : OUT <= 10;  //240 / 23 = 10
    16'b11110000_00011000 : OUT <= 10;  //240 / 24 = 10
    16'b11110000_00011001 : OUT <= 9;  //240 / 25 = 9
    16'b11110000_00011010 : OUT <= 9;  //240 / 26 = 9
    16'b11110000_00011011 : OUT <= 8;  //240 / 27 = 8
    16'b11110000_00011100 : OUT <= 8;  //240 / 28 = 8
    16'b11110000_00011101 : OUT <= 8;  //240 / 29 = 8
    16'b11110000_00011110 : OUT <= 8;  //240 / 30 = 8
    16'b11110000_00011111 : OUT <= 7;  //240 / 31 = 7
    16'b11110000_00100000 : OUT <= 7;  //240 / 32 = 7
    16'b11110000_00100001 : OUT <= 7;  //240 / 33 = 7
    16'b11110000_00100010 : OUT <= 7;  //240 / 34 = 7
    16'b11110000_00100011 : OUT <= 6;  //240 / 35 = 6
    16'b11110000_00100100 : OUT <= 6;  //240 / 36 = 6
    16'b11110000_00100101 : OUT <= 6;  //240 / 37 = 6
    16'b11110000_00100110 : OUT <= 6;  //240 / 38 = 6
    16'b11110000_00100111 : OUT <= 6;  //240 / 39 = 6
    16'b11110000_00101000 : OUT <= 6;  //240 / 40 = 6
    16'b11110000_00101001 : OUT <= 5;  //240 / 41 = 5
    16'b11110000_00101010 : OUT <= 5;  //240 / 42 = 5
    16'b11110000_00101011 : OUT <= 5;  //240 / 43 = 5
    16'b11110000_00101100 : OUT <= 5;  //240 / 44 = 5
    16'b11110000_00101101 : OUT <= 5;  //240 / 45 = 5
    16'b11110000_00101110 : OUT <= 5;  //240 / 46 = 5
    16'b11110000_00101111 : OUT <= 5;  //240 / 47 = 5
    16'b11110000_00110000 : OUT <= 5;  //240 / 48 = 5
    16'b11110000_00110001 : OUT <= 4;  //240 / 49 = 4
    16'b11110000_00110010 : OUT <= 4;  //240 / 50 = 4
    16'b11110000_00110011 : OUT <= 4;  //240 / 51 = 4
    16'b11110000_00110100 : OUT <= 4;  //240 / 52 = 4
    16'b11110000_00110101 : OUT <= 4;  //240 / 53 = 4
    16'b11110000_00110110 : OUT <= 4;  //240 / 54 = 4
    16'b11110000_00110111 : OUT <= 4;  //240 / 55 = 4
    16'b11110000_00111000 : OUT <= 4;  //240 / 56 = 4
    16'b11110000_00111001 : OUT <= 4;  //240 / 57 = 4
    16'b11110000_00111010 : OUT <= 4;  //240 / 58 = 4
    16'b11110000_00111011 : OUT <= 4;  //240 / 59 = 4
    16'b11110000_00111100 : OUT <= 4;  //240 / 60 = 4
    16'b11110000_00111101 : OUT <= 3;  //240 / 61 = 3
    16'b11110000_00111110 : OUT <= 3;  //240 / 62 = 3
    16'b11110000_00111111 : OUT <= 3;  //240 / 63 = 3
    16'b11110000_01000000 : OUT <= 3;  //240 / 64 = 3
    16'b11110000_01000001 : OUT <= 3;  //240 / 65 = 3
    16'b11110000_01000010 : OUT <= 3;  //240 / 66 = 3
    16'b11110000_01000011 : OUT <= 3;  //240 / 67 = 3
    16'b11110000_01000100 : OUT <= 3;  //240 / 68 = 3
    16'b11110000_01000101 : OUT <= 3;  //240 / 69 = 3
    16'b11110000_01000110 : OUT <= 3;  //240 / 70 = 3
    16'b11110000_01000111 : OUT <= 3;  //240 / 71 = 3
    16'b11110000_01001000 : OUT <= 3;  //240 / 72 = 3
    16'b11110000_01001001 : OUT <= 3;  //240 / 73 = 3
    16'b11110000_01001010 : OUT <= 3;  //240 / 74 = 3
    16'b11110000_01001011 : OUT <= 3;  //240 / 75 = 3
    16'b11110000_01001100 : OUT <= 3;  //240 / 76 = 3
    16'b11110000_01001101 : OUT <= 3;  //240 / 77 = 3
    16'b11110000_01001110 : OUT <= 3;  //240 / 78 = 3
    16'b11110000_01001111 : OUT <= 3;  //240 / 79 = 3
    16'b11110000_01010000 : OUT <= 3;  //240 / 80 = 3
    16'b11110000_01010001 : OUT <= 2;  //240 / 81 = 2
    16'b11110000_01010010 : OUT <= 2;  //240 / 82 = 2
    16'b11110000_01010011 : OUT <= 2;  //240 / 83 = 2
    16'b11110000_01010100 : OUT <= 2;  //240 / 84 = 2
    16'b11110000_01010101 : OUT <= 2;  //240 / 85 = 2
    16'b11110000_01010110 : OUT <= 2;  //240 / 86 = 2
    16'b11110000_01010111 : OUT <= 2;  //240 / 87 = 2
    16'b11110000_01011000 : OUT <= 2;  //240 / 88 = 2
    16'b11110000_01011001 : OUT <= 2;  //240 / 89 = 2
    16'b11110000_01011010 : OUT <= 2;  //240 / 90 = 2
    16'b11110000_01011011 : OUT <= 2;  //240 / 91 = 2
    16'b11110000_01011100 : OUT <= 2;  //240 / 92 = 2
    16'b11110000_01011101 : OUT <= 2;  //240 / 93 = 2
    16'b11110000_01011110 : OUT <= 2;  //240 / 94 = 2
    16'b11110000_01011111 : OUT <= 2;  //240 / 95 = 2
    16'b11110000_01100000 : OUT <= 2;  //240 / 96 = 2
    16'b11110000_01100001 : OUT <= 2;  //240 / 97 = 2
    16'b11110000_01100010 : OUT <= 2;  //240 / 98 = 2
    16'b11110000_01100011 : OUT <= 2;  //240 / 99 = 2
    16'b11110000_01100100 : OUT <= 2;  //240 / 100 = 2
    16'b11110000_01100101 : OUT <= 2;  //240 / 101 = 2
    16'b11110000_01100110 : OUT <= 2;  //240 / 102 = 2
    16'b11110000_01100111 : OUT <= 2;  //240 / 103 = 2
    16'b11110000_01101000 : OUT <= 2;  //240 / 104 = 2
    16'b11110000_01101001 : OUT <= 2;  //240 / 105 = 2
    16'b11110000_01101010 : OUT <= 2;  //240 / 106 = 2
    16'b11110000_01101011 : OUT <= 2;  //240 / 107 = 2
    16'b11110000_01101100 : OUT <= 2;  //240 / 108 = 2
    16'b11110000_01101101 : OUT <= 2;  //240 / 109 = 2
    16'b11110000_01101110 : OUT <= 2;  //240 / 110 = 2
    16'b11110000_01101111 : OUT <= 2;  //240 / 111 = 2
    16'b11110000_01110000 : OUT <= 2;  //240 / 112 = 2
    16'b11110000_01110001 : OUT <= 2;  //240 / 113 = 2
    16'b11110000_01110010 : OUT <= 2;  //240 / 114 = 2
    16'b11110000_01110011 : OUT <= 2;  //240 / 115 = 2
    16'b11110000_01110100 : OUT <= 2;  //240 / 116 = 2
    16'b11110000_01110101 : OUT <= 2;  //240 / 117 = 2
    16'b11110000_01110110 : OUT <= 2;  //240 / 118 = 2
    16'b11110000_01110111 : OUT <= 2;  //240 / 119 = 2
    16'b11110000_01111000 : OUT <= 2;  //240 / 120 = 2
    16'b11110000_01111001 : OUT <= 1;  //240 / 121 = 1
    16'b11110000_01111010 : OUT <= 1;  //240 / 122 = 1
    16'b11110000_01111011 : OUT <= 1;  //240 / 123 = 1
    16'b11110000_01111100 : OUT <= 1;  //240 / 124 = 1
    16'b11110000_01111101 : OUT <= 1;  //240 / 125 = 1
    16'b11110000_01111110 : OUT <= 1;  //240 / 126 = 1
    16'b11110000_01111111 : OUT <= 1;  //240 / 127 = 1
    16'b11110000_10000000 : OUT <= 1;  //240 / 128 = 1
    16'b11110000_10000001 : OUT <= 1;  //240 / 129 = 1
    16'b11110000_10000010 : OUT <= 1;  //240 / 130 = 1
    16'b11110000_10000011 : OUT <= 1;  //240 / 131 = 1
    16'b11110000_10000100 : OUT <= 1;  //240 / 132 = 1
    16'b11110000_10000101 : OUT <= 1;  //240 / 133 = 1
    16'b11110000_10000110 : OUT <= 1;  //240 / 134 = 1
    16'b11110000_10000111 : OUT <= 1;  //240 / 135 = 1
    16'b11110000_10001000 : OUT <= 1;  //240 / 136 = 1
    16'b11110000_10001001 : OUT <= 1;  //240 / 137 = 1
    16'b11110000_10001010 : OUT <= 1;  //240 / 138 = 1
    16'b11110000_10001011 : OUT <= 1;  //240 / 139 = 1
    16'b11110000_10001100 : OUT <= 1;  //240 / 140 = 1
    16'b11110000_10001101 : OUT <= 1;  //240 / 141 = 1
    16'b11110000_10001110 : OUT <= 1;  //240 / 142 = 1
    16'b11110000_10001111 : OUT <= 1;  //240 / 143 = 1
    16'b11110000_10010000 : OUT <= 1;  //240 / 144 = 1
    16'b11110000_10010001 : OUT <= 1;  //240 / 145 = 1
    16'b11110000_10010010 : OUT <= 1;  //240 / 146 = 1
    16'b11110000_10010011 : OUT <= 1;  //240 / 147 = 1
    16'b11110000_10010100 : OUT <= 1;  //240 / 148 = 1
    16'b11110000_10010101 : OUT <= 1;  //240 / 149 = 1
    16'b11110000_10010110 : OUT <= 1;  //240 / 150 = 1
    16'b11110000_10010111 : OUT <= 1;  //240 / 151 = 1
    16'b11110000_10011000 : OUT <= 1;  //240 / 152 = 1
    16'b11110000_10011001 : OUT <= 1;  //240 / 153 = 1
    16'b11110000_10011010 : OUT <= 1;  //240 / 154 = 1
    16'b11110000_10011011 : OUT <= 1;  //240 / 155 = 1
    16'b11110000_10011100 : OUT <= 1;  //240 / 156 = 1
    16'b11110000_10011101 : OUT <= 1;  //240 / 157 = 1
    16'b11110000_10011110 : OUT <= 1;  //240 / 158 = 1
    16'b11110000_10011111 : OUT <= 1;  //240 / 159 = 1
    16'b11110000_10100000 : OUT <= 1;  //240 / 160 = 1
    16'b11110000_10100001 : OUT <= 1;  //240 / 161 = 1
    16'b11110000_10100010 : OUT <= 1;  //240 / 162 = 1
    16'b11110000_10100011 : OUT <= 1;  //240 / 163 = 1
    16'b11110000_10100100 : OUT <= 1;  //240 / 164 = 1
    16'b11110000_10100101 : OUT <= 1;  //240 / 165 = 1
    16'b11110000_10100110 : OUT <= 1;  //240 / 166 = 1
    16'b11110000_10100111 : OUT <= 1;  //240 / 167 = 1
    16'b11110000_10101000 : OUT <= 1;  //240 / 168 = 1
    16'b11110000_10101001 : OUT <= 1;  //240 / 169 = 1
    16'b11110000_10101010 : OUT <= 1;  //240 / 170 = 1
    16'b11110000_10101011 : OUT <= 1;  //240 / 171 = 1
    16'b11110000_10101100 : OUT <= 1;  //240 / 172 = 1
    16'b11110000_10101101 : OUT <= 1;  //240 / 173 = 1
    16'b11110000_10101110 : OUT <= 1;  //240 / 174 = 1
    16'b11110000_10101111 : OUT <= 1;  //240 / 175 = 1
    16'b11110000_10110000 : OUT <= 1;  //240 / 176 = 1
    16'b11110000_10110001 : OUT <= 1;  //240 / 177 = 1
    16'b11110000_10110010 : OUT <= 1;  //240 / 178 = 1
    16'b11110000_10110011 : OUT <= 1;  //240 / 179 = 1
    16'b11110000_10110100 : OUT <= 1;  //240 / 180 = 1
    16'b11110000_10110101 : OUT <= 1;  //240 / 181 = 1
    16'b11110000_10110110 : OUT <= 1;  //240 / 182 = 1
    16'b11110000_10110111 : OUT <= 1;  //240 / 183 = 1
    16'b11110000_10111000 : OUT <= 1;  //240 / 184 = 1
    16'b11110000_10111001 : OUT <= 1;  //240 / 185 = 1
    16'b11110000_10111010 : OUT <= 1;  //240 / 186 = 1
    16'b11110000_10111011 : OUT <= 1;  //240 / 187 = 1
    16'b11110000_10111100 : OUT <= 1;  //240 / 188 = 1
    16'b11110000_10111101 : OUT <= 1;  //240 / 189 = 1
    16'b11110000_10111110 : OUT <= 1;  //240 / 190 = 1
    16'b11110000_10111111 : OUT <= 1;  //240 / 191 = 1
    16'b11110000_11000000 : OUT <= 1;  //240 / 192 = 1
    16'b11110000_11000001 : OUT <= 1;  //240 / 193 = 1
    16'b11110000_11000010 : OUT <= 1;  //240 / 194 = 1
    16'b11110000_11000011 : OUT <= 1;  //240 / 195 = 1
    16'b11110000_11000100 : OUT <= 1;  //240 / 196 = 1
    16'b11110000_11000101 : OUT <= 1;  //240 / 197 = 1
    16'b11110000_11000110 : OUT <= 1;  //240 / 198 = 1
    16'b11110000_11000111 : OUT <= 1;  //240 / 199 = 1
    16'b11110000_11001000 : OUT <= 1;  //240 / 200 = 1
    16'b11110000_11001001 : OUT <= 1;  //240 / 201 = 1
    16'b11110000_11001010 : OUT <= 1;  //240 / 202 = 1
    16'b11110000_11001011 : OUT <= 1;  //240 / 203 = 1
    16'b11110000_11001100 : OUT <= 1;  //240 / 204 = 1
    16'b11110000_11001101 : OUT <= 1;  //240 / 205 = 1
    16'b11110000_11001110 : OUT <= 1;  //240 / 206 = 1
    16'b11110000_11001111 : OUT <= 1;  //240 / 207 = 1
    16'b11110000_11010000 : OUT <= 1;  //240 / 208 = 1
    16'b11110000_11010001 : OUT <= 1;  //240 / 209 = 1
    16'b11110000_11010010 : OUT <= 1;  //240 / 210 = 1
    16'b11110000_11010011 : OUT <= 1;  //240 / 211 = 1
    16'b11110000_11010100 : OUT <= 1;  //240 / 212 = 1
    16'b11110000_11010101 : OUT <= 1;  //240 / 213 = 1
    16'b11110000_11010110 : OUT <= 1;  //240 / 214 = 1
    16'b11110000_11010111 : OUT <= 1;  //240 / 215 = 1
    16'b11110000_11011000 : OUT <= 1;  //240 / 216 = 1
    16'b11110000_11011001 : OUT <= 1;  //240 / 217 = 1
    16'b11110000_11011010 : OUT <= 1;  //240 / 218 = 1
    16'b11110000_11011011 : OUT <= 1;  //240 / 219 = 1
    16'b11110000_11011100 : OUT <= 1;  //240 / 220 = 1
    16'b11110000_11011101 : OUT <= 1;  //240 / 221 = 1
    16'b11110000_11011110 : OUT <= 1;  //240 / 222 = 1
    16'b11110000_11011111 : OUT <= 1;  //240 / 223 = 1
    16'b11110000_11100000 : OUT <= 1;  //240 / 224 = 1
    16'b11110000_11100001 : OUT <= 1;  //240 / 225 = 1
    16'b11110000_11100010 : OUT <= 1;  //240 / 226 = 1
    16'b11110000_11100011 : OUT <= 1;  //240 / 227 = 1
    16'b11110000_11100100 : OUT <= 1;  //240 / 228 = 1
    16'b11110000_11100101 : OUT <= 1;  //240 / 229 = 1
    16'b11110000_11100110 : OUT <= 1;  //240 / 230 = 1
    16'b11110000_11100111 : OUT <= 1;  //240 / 231 = 1
    16'b11110000_11101000 : OUT <= 1;  //240 / 232 = 1
    16'b11110000_11101001 : OUT <= 1;  //240 / 233 = 1
    16'b11110000_11101010 : OUT <= 1;  //240 / 234 = 1
    16'b11110000_11101011 : OUT <= 1;  //240 / 235 = 1
    16'b11110000_11101100 : OUT <= 1;  //240 / 236 = 1
    16'b11110000_11101101 : OUT <= 1;  //240 / 237 = 1
    16'b11110000_11101110 : OUT <= 1;  //240 / 238 = 1
    16'b11110000_11101111 : OUT <= 1;  //240 / 239 = 1
    16'b11110000_11110000 : OUT <= 1;  //240 / 240 = 1
    16'b11110000_11110001 : OUT <= 0;  //240 / 241 = 0
    16'b11110000_11110010 : OUT <= 0;  //240 / 242 = 0
    16'b11110000_11110011 : OUT <= 0;  //240 / 243 = 0
    16'b11110000_11110100 : OUT <= 0;  //240 / 244 = 0
    16'b11110000_11110101 : OUT <= 0;  //240 / 245 = 0
    16'b11110000_11110110 : OUT <= 0;  //240 / 246 = 0
    16'b11110000_11110111 : OUT <= 0;  //240 / 247 = 0
    16'b11110000_11111000 : OUT <= 0;  //240 / 248 = 0
    16'b11110000_11111001 : OUT <= 0;  //240 / 249 = 0
    16'b11110000_11111010 : OUT <= 0;  //240 / 250 = 0
    16'b11110000_11111011 : OUT <= 0;  //240 / 251 = 0
    16'b11110000_11111100 : OUT <= 0;  //240 / 252 = 0
    16'b11110000_11111101 : OUT <= 0;  //240 / 253 = 0
    16'b11110000_11111110 : OUT <= 0;  //240 / 254 = 0
    16'b11110000_11111111 : OUT <= 0;  //240 / 255 = 0
    16'b11110001_00000000 : OUT <= 0;  //241 / 0 = 0
    16'b11110001_00000001 : OUT <= 241;  //241 / 1 = 241
    16'b11110001_00000010 : OUT <= 120;  //241 / 2 = 120
    16'b11110001_00000011 : OUT <= 80;  //241 / 3 = 80
    16'b11110001_00000100 : OUT <= 60;  //241 / 4 = 60
    16'b11110001_00000101 : OUT <= 48;  //241 / 5 = 48
    16'b11110001_00000110 : OUT <= 40;  //241 / 6 = 40
    16'b11110001_00000111 : OUT <= 34;  //241 / 7 = 34
    16'b11110001_00001000 : OUT <= 30;  //241 / 8 = 30
    16'b11110001_00001001 : OUT <= 26;  //241 / 9 = 26
    16'b11110001_00001010 : OUT <= 24;  //241 / 10 = 24
    16'b11110001_00001011 : OUT <= 21;  //241 / 11 = 21
    16'b11110001_00001100 : OUT <= 20;  //241 / 12 = 20
    16'b11110001_00001101 : OUT <= 18;  //241 / 13 = 18
    16'b11110001_00001110 : OUT <= 17;  //241 / 14 = 17
    16'b11110001_00001111 : OUT <= 16;  //241 / 15 = 16
    16'b11110001_00010000 : OUT <= 15;  //241 / 16 = 15
    16'b11110001_00010001 : OUT <= 14;  //241 / 17 = 14
    16'b11110001_00010010 : OUT <= 13;  //241 / 18 = 13
    16'b11110001_00010011 : OUT <= 12;  //241 / 19 = 12
    16'b11110001_00010100 : OUT <= 12;  //241 / 20 = 12
    16'b11110001_00010101 : OUT <= 11;  //241 / 21 = 11
    16'b11110001_00010110 : OUT <= 10;  //241 / 22 = 10
    16'b11110001_00010111 : OUT <= 10;  //241 / 23 = 10
    16'b11110001_00011000 : OUT <= 10;  //241 / 24 = 10
    16'b11110001_00011001 : OUT <= 9;  //241 / 25 = 9
    16'b11110001_00011010 : OUT <= 9;  //241 / 26 = 9
    16'b11110001_00011011 : OUT <= 8;  //241 / 27 = 8
    16'b11110001_00011100 : OUT <= 8;  //241 / 28 = 8
    16'b11110001_00011101 : OUT <= 8;  //241 / 29 = 8
    16'b11110001_00011110 : OUT <= 8;  //241 / 30 = 8
    16'b11110001_00011111 : OUT <= 7;  //241 / 31 = 7
    16'b11110001_00100000 : OUT <= 7;  //241 / 32 = 7
    16'b11110001_00100001 : OUT <= 7;  //241 / 33 = 7
    16'b11110001_00100010 : OUT <= 7;  //241 / 34 = 7
    16'b11110001_00100011 : OUT <= 6;  //241 / 35 = 6
    16'b11110001_00100100 : OUT <= 6;  //241 / 36 = 6
    16'b11110001_00100101 : OUT <= 6;  //241 / 37 = 6
    16'b11110001_00100110 : OUT <= 6;  //241 / 38 = 6
    16'b11110001_00100111 : OUT <= 6;  //241 / 39 = 6
    16'b11110001_00101000 : OUT <= 6;  //241 / 40 = 6
    16'b11110001_00101001 : OUT <= 5;  //241 / 41 = 5
    16'b11110001_00101010 : OUT <= 5;  //241 / 42 = 5
    16'b11110001_00101011 : OUT <= 5;  //241 / 43 = 5
    16'b11110001_00101100 : OUT <= 5;  //241 / 44 = 5
    16'b11110001_00101101 : OUT <= 5;  //241 / 45 = 5
    16'b11110001_00101110 : OUT <= 5;  //241 / 46 = 5
    16'b11110001_00101111 : OUT <= 5;  //241 / 47 = 5
    16'b11110001_00110000 : OUT <= 5;  //241 / 48 = 5
    16'b11110001_00110001 : OUT <= 4;  //241 / 49 = 4
    16'b11110001_00110010 : OUT <= 4;  //241 / 50 = 4
    16'b11110001_00110011 : OUT <= 4;  //241 / 51 = 4
    16'b11110001_00110100 : OUT <= 4;  //241 / 52 = 4
    16'b11110001_00110101 : OUT <= 4;  //241 / 53 = 4
    16'b11110001_00110110 : OUT <= 4;  //241 / 54 = 4
    16'b11110001_00110111 : OUT <= 4;  //241 / 55 = 4
    16'b11110001_00111000 : OUT <= 4;  //241 / 56 = 4
    16'b11110001_00111001 : OUT <= 4;  //241 / 57 = 4
    16'b11110001_00111010 : OUT <= 4;  //241 / 58 = 4
    16'b11110001_00111011 : OUT <= 4;  //241 / 59 = 4
    16'b11110001_00111100 : OUT <= 4;  //241 / 60 = 4
    16'b11110001_00111101 : OUT <= 3;  //241 / 61 = 3
    16'b11110001_00111110 : OUT <= 3;  //241 / 62 = 3
    16'b11110001_00111111 : OUT <= 3;  //241 / 63 = 3
    16'b11110001_01000000 : OUT <= 3;  //241 / 64 = 3
    16'b11110001_01000001 : OUT <= 3;  //241 / 65 = 3
    16'b11110001_01000010 : OUT <= 3;  //241 / 66 = 3
    16'b11110001_01000011 : OUT <= 3;  //241 / 67 = 3
    16'b11110001_01000100 : OUT <= 3;  //241 / 68 = 3
    16'b11110001_01000101 : OUT <= 3;  //241 / 69 = 3
    16'b11110001_01000110 : OUT <= 3;  //241 / 70 = 3
    16'b11110001_01000111 : OUT <= 3;  //241 / 71 = 3
    16'b11110001_01001000 : OUT <= 3;  //241 / 72 = 3
    16'b11110001_01001001 : OUT <= 3;  //241 / 73 = 3
    16'b11110001_01001010 : OUT <= 3;  //241 / 74 = 3
    16'b11110001_01001011 : OUT <= 3;  //241 / 75 = 3
    16'b11110001_01001100 : OUT <= 3;  //241 / 76 = 3
    16'b11110001_01001101 : OUT <= 3;  //241 / 77 = 3
    16'b11110001_01001110 : OUT <= 3;  //241 / 78 = 3
    16'b11110001_01001111 : OUT <= 3;  //241 / 79 = 3
    16'b11110001_01010000 : OUT <= 3;  //241 / 80 = 3
    16'b11110001_01010001 : OUT <= 2;  //241 / 81 = 2
    16'b11110001_01010010 : OUT <= 2;  //241 / 82 = 2
    16'b11110001_01010011 : OUT <= 2;  //241 / 83 = 2
    16'b11110001_01010100 : OUT <= 2;  //241 / 84 = 2
    16'b11110001_01010101 : OUT <= 2;  //241 / 85 = 2
    16'b11110001_01010110 : OUT <= 2;  //241 / 86 = 2
    16'b11110001_01010111 : OUT <= 2;  //241 / 87 = 2
    16'b11110001_01011000 : OUT <= 2;  //241 / 88 = 2
    16'b11110001_01011001 : OUT <= 2;  //241 / 89 = 2
    16'b11110001_01011010 : OUT <= 2;  //241 / 90 = 2
    16'b11110001_01011011 : OUT <= 2;  //241 / 91 = 2
    16'b11110001_01011100 : OUT <= 2;  //241 / 92 = 2
    16'b11110001_01011101 : OUT <= 2;  //241 / 93 = 2
    16'b11110001_01011110 : OUT <= 2;  //241 / 94 = 2
    16'b11110001_01011111 : OUT <= 2;  //241 / 95 = 2
    16'b11110001_01100000 : OUT <= 2;  //241 / 96 = 2
    16'b11110001_01100001 : OUT <= 2;  //241 / 97 = 2
    16'b11110001_01100010 : OUT <= 2;  //241 / 98 = 2
    16'b11110001_01100011 : OUT <= 2;  //241 / 99 = 2
    16'b11110001_01100100 : OUT <= 2;  //241 / 100 = 2
    16'b11110001_01100101 : OUT <= 2;  //241 / 101 = 2
    16'b11110001_01100110 : OUT <= 2;  //241 / 102 = 2
    16'b11110001_01100111 : OUT <= 2;  //241 / 103 = 2
    16'b11110001_01101000 : OUT <= 2;  //241 / 104 = 2
    16'b11110001_01101001 : OUT <= 2;  //241 / 105 = 2
    16'b11110001_01101010 : OUT <= 2;  //241 / 106 = 2
    16'b11110001_01101011 : OUT <= 2;  //241 / 107 = 2
    16'b11110001_01101100 : OUT <= 2;  //241 / 108 = 2
    16'b11110001_01101101 : OUT <= 2;  //241 / 109 = 2
    16'b11110001_01101110 : OUT <= 2;  //241 / 110 = 2
    16'b11110001_01101111 : OUT <= 2;  //241 / 111 = 2
    16'b11110001_01110000 : OUT <= 2;  //241 / 112 = 2
    16'b11110001_01110001 : OUT <= 2;  //241 / 113 = 2
    16'b11110001_01110010 : OUT <= 2;  //241 / 114 = 2
    16'b11110001_01110011 : OUT <= 2;  //241 / 115 = 2
    16'b11110001_01110100 : OUT <= 2;  //241 / 116 = 2
    16'b11110001_01110101 : OUT <= 2;  //241 / 117 = 2
    16'b11110001_01110110 : OUT <= 2;  //241 / 118 = 2
    16'b11110001_01110111 : OUT <= 2;  //241 / 119 = 2
    16'b11110001_01111000 : OUT <= 2;  //241 / 120 = 2
    16'b11110001_01111001 : OUT <= 1;  //241 / 121 = 1
    16'b11110001_01111010 : OUT <= 1;  //241 / 122 = 1
    16'b11110001_01111011 : OUT <= 1;  //241 / 123 = 1
    16'b11110001_01111100 : OUT <= 1;  //241 / 124 = 1
    16'b11110001_01111101 : OUT <= 1;  //241 / 125 = 1
    16'b11110001_01111110 : OUT <= 1;  //241 / 126 = 1
    16'b11110001_01111111 : OUT <= 1;  //241 / 127 = 1
    16'b11110001_10000000 : OUT <= 1;  //241 / 128 = 1
    16'b11110001_10000001 : OUT <= 1;  //241 / 129 = 1
    16'b11110001_10000010 : OUT <= 1;  //241 / 130 = 1
    16'b11110001_10000011 : OUT <= 1;  //241 / 131 = 1
    16'b11110001_10000100 : OUT <= 1;  //241 / 132 = 1
    16'b11110001_10000101 : OUT <= 1;  //241 / 133 = 1
    16'b11110001_10000110 : OUT <= 1;  //241 / 134 = 1
    16'b11110001_10000111 : OUT <= 1;  //241 / 135 = 1
    16'b11110001_10001000 : OUT <= 1;  //241 / 136 = 1
    16'b11110001_10001001 : OUT <= 1;  //241 / 137 = 1
    16'b11110001_10001010 : OUT <= 1;  //241 / 138 = 1
    16'b11110001_10001011 : OUT <= 1;  //241 / 139 = 1
    16'b11110001_10001100 : OUT <= 1;  //241 / 140 = 1
    16'b11110001_10001101 : OUT <= 1;  //241 / 141 = 1
    16'b11110001_10001110 : OUT <= 1;  //241 / 142 = 1
    16'b11110001_10001111 : OUT <= 1;  //241 / 143 = 1
    16'b11110001_10010000 : OUT <= 1;  //241 / 144 = 1
    16'b11110001_10010001 : OUT <= 1;  //241 / 145 = 1
    16'b11110001_10010010 : OUT <= 1;  //241 / 146 = 1
    16'b11110001_10010011 : OUT <= 1;  //241 / 147 = 1
    16'b11110001_10010100 : OUT <= 1;  //241 / 148 = 1
    16'b11110001_10010101 : OUT <= 1;  //241 / 149 = 1
    16'b11110001_10010110 : OUT <= 1;  //241 / 150 = 1
    16'b11110001_10010111 : OUT <= 1;  //241 / 151 = 1
    16'b11110001_10011000 : OUT <= 1;  //241 / 152 = 1
    16'b11110001_10011001 : OUT <= 1;  //241 / 153 = 1
    16'b11110001_10011010 : OUT <= 1;  //241 / 154 = 1
    16'b11110001_10011011 : OUT <= 1;  //241 / 155 = 1
    16'b11110001_10011100 : OUT <= 1;  //241 / 156 = 1
    16'b11110001_10011101 : OUT <= 1;  //241 / 157 = 1
    16'b11110001_10011110 : OUT <= 1;  //241 / 158 = 1
    16'b11110001_10011111 : OUT <= 1;  //241 / 159 = 1
    16'b11110001_10100000 : OUT <= 1;  //241 / 160 = 1
    16'b11110001_10100001 : OUT <= 1;  //241 / 161 = 1
    16'b11110001_10100010 : OUT <= 1;  //241 / 162 = 1
    16'b11110001_10100011 : OUT <= 1;  //241 / 163 = 1
    16'b11110001_10100100 : OUT <= 1;  //241 / 164 = 1
    16'b11110001_10100101 : OUT <= 1;  //241 / 165 = 1
    16'b11110001_10100110 : OUT <= 1;  //241 / 166 = 1
    16'b11110001_10100111 : OUT <= 1;  //241 / 167 = 1
    16'b11110001_10101000 : OUT <= 1;  //241 / 168 = 1
    16'b11110001_10101001 : OUT <= 1;  //241 / 169 = 1
    16'b11110001_10101010 : OUT <= 1;  //241 / 170 = 1
    16'b11110001_10101011 : OUT <= 1;  //241 / 171 = 1
    16'b11110001_10101100 : OUT <= 1;  //241 / 172 = 1
    16'b11110001_10101101 : OUT <= 1;  //241 / 173 = 1
    16'b11110001_10101110 : OUT <= 1;  //241 / 174 = 1
    16'b11110001_10101111 : OUT <= 1;  //241 / 175 = 1
    16'b11110001_10110000 : OUT <= 1;  //241 / 176 = 1
    16'b11110001_10110001 : OUT <= 1;  //241 / 177 = 1
    16'b11110001_10110010 : OUT <= 1;  //241 / 178 = 1
    16'b11110001_10110011 : OUT <= 1;  //241 / 179 = 1
    16'b11110001_10110100 : OUT <= 1;  //241 / 180 = 1
    16'b11110001_10110101 : OUT <= 1;  //241 / 181 = 1
    16'b11110001_10110110 : OUT <= 1;  //241 / 182 = 1
    16'b11110001_10110111 : OUT <= 1;  //241 / 183 = 1
    16'b11110001_10111000 : OUT <= 1;  //241 / 184 = 1
    16'b11110001_10111001 : OUT <= 1;  //241 / 185 = 1
    16'b11110001_10111010 : OUT <= 1;  //241 / 186 = 1
    16'b11110001_10111011 : OUT <= 1;  //241 / 187 = 1
    16'b11110001_10111100 : OUT <= 1;  //241 / 188 = 1
    16'b11110001_10111101 : OUT <= 1;  //241 / 189 = 1
    16'b11110001_10111110 : OUT <= 1;  //241 / 190 = 1
    16'b11110001_10111111 : OUT <= 1;  //241 / 191 = 1
    16'b11110001_11000000 : OUT <= 1;  //241 / 192 = 1
    16'b11110001_11000001 : OUT <= 1;  //241 / 193 = 1
    16'b11110001_11000010 : OUT <= 1;  //241 / 194 = 1
    16'b11110001_11000011 : OUT <= 1;  //241 / 195 = 1
    16'b11110001_11000100 : OUT <= 1;  //241 / 196 = 1
    16'b11110001_11000101 : OUT <= 1;  //241 / 197 = 1
    16'b11110001_11000110 : OUT <= 1;  //241 / 198 = 1
    16'b11110001_11000111 : OUT <= 1;  //241 / 199 = 1
    16'b11110001_11001000 : OUT <= 1;  //241 / 200 = 1
    16'b11110001_11001001 : OUT <= 1;  //241 / 201 = 1
    16'b11110001_11001010 : OUT <= 1;  //241 / 202 = 1
    16'b11110001_11001011 : OUT <= 1;  //241 / 203 = 1
    16'b11110001_11001100 : OUT <= 1;  //241 / 204 = 1
    16'b11110001_11001101 : OUT <= 1;  //241 / 205 = 1
    16'b11110001_11001110 : OUT <= 1;  //241 / 206 = 1
    16'b11110001_11001111 : OUT <= 1;  //241 / 207 = 1
    16'b11110001_11010000 : OUT <= 1;  //241 / 208 = 1
    16'b11110001_11010001 : OUT <= 1;  //241 / 209 = 1
    16'b11110001_11010010 : OUT <= 1;  //241 / 210 = 1
    16'b11110001_11010011 : OUT <= 1;  //241 / 211 = 1
    16'b11110001_11010100 : OUT <= 1;  //241 / 212 = 1
    16'b11110001_11010101 : OUT <= 1;  //241 / 213 = 1
    16'b11110001_11010110 : OUT <= 1;  //241 / 214 = 1
    16'b11110001_11010111 : OUT <= 1;  //241 / 215 = 1
    16'b11110001_11011000 : OUT <= 1;  //241 / 216 = 1
    16'b11110001_11011001 : OUT <= 1;  //241 / 217 = 1
    16'b11110001_11011010 : OUT <= 1;  //241 / 218 = 1
    16'b11110001_11011011 : OUT <= 1;  //241 / 219 = 1
    16'b11110001_11011100 : OUT <= 1;  //241 / 220 = 1
    16'b11110001_11011101 : OUT <= 1;  //241 / 221 = 1
    16'b11110001_11011110 : OUT <= 1;  //241 / 222 = 1
    16'b11110001_11011111 : OUT <= 1;  //241 / 223 = 1
    16'b11110001_11100000 : OUT <= 1;  //241 / 224 = 1
    16'b11110001_11100001 : OUT <= 1;  //241 / 225 = 1
    16'b11110001_11100010 : OUT <= 1;  //241 / 226 = 1
    16'b11110001_11100011 : OUT <= 1;  //241 / 227 = 1
    16'b11110001_11100100 : OUT <= 1;  //241 / 228 = 1
    16'b11110001_11100101 : OUT <= 1;  //241 / 229 = 1
    16'b11110001_11100110 : OUT <= 1;  //241 / 230 = 1
    16'b11110001_11100111 : OUT <= 1;  //241 / 231 = 1
    16'b11110001_11101000 : OUT <= 1;  //241 / 232 = 1
    16'b11110001_11101001 : OUT <= 1;  //241 / 233 = 1
    16'b11110001_11101010 : OUT <= 1;  //241 / 234 = 1
    16'b11110001_11101011 : OUT <= 1;  //241 / 235 = 1
    16'b11110001_11101100 : OUT <= 1;  //241 / 236 = 1
    16'b11110001_11101101 : OUT <= 1;  //241 / 237 = 1
    16'b11110001_11101110 : OUT <= 1;  //241 / 238 = 1
    16'b11110001_11101111 : OUT <= 1;  //241 / 239 = 1
    16'b11110001_11110000 : OUT <= 1;  //241 / 240 = 1
    16'b11110001_11110001 : OUT <= 1;  //241 / 241 = 1
    16'b11110001_11110010 : OUT <= 0;  //241 / 242 = 0
    16'b11110001_11110011 : OUT <= 0;  //241 / 243 = 0
    16'b11110001_11110100 : OUT <= 0;  //241 / 244 = 0
    16'b11110001_11110101 : OUT <= 0;  //241 / 245 = 0
    16'b11110001_11110110 : OUT <= 0;  //241 / 246 = 0
    16'b11110001_11110111 : OUT <= 0;  //241 / 247 = 0
    16'b11110001_11111000 : OUT <= 0;  //241 / 248 = 0
    16'b11110001_11111001 : OUT <= 0;  //241 / 249 = 0
    16'b11110001_11111010 : OUT <= 0;  //241 / 250 = 0
    16'b11110001_11111011 : OUT <= 0;  //241 / 251 = 0
    16'b11110001_11111100 : OUT <= 0;  //241 / 252 = 0
    16'b11110001_11111101 : OUT <= 0;  //241 / 253 = 0
    16'b11110001_11111110 : OUT <= 0;  //241 / 254 = 0
    16'b11110001_11111111 : OUT <= 0;  //241 / 255 = 0
    16'b11110010_00000000 : OUT <= 0;  //242 / 0 = 0
    16'b11110010_00000001 : OUT <= 242;  //242 / 1 = 242
    16'b11110010_00000010 : OUT <= 121;  //242 / 2 = 121
    16'b11110010_00000011 : OUT <= 80;  //242 / 3 = 80
    16'b11110010_00000100 : OUT <= 60;  //242 / 4 = 60
    16'b11110010_00000101 : OUT <= 48;  //242 / 5 = 48
    16'b11110010_00000110 : OUT <= 40;  //242 / 6 = 40
    16'b11110010_00000111 : OUT <= 34;  //242 / 7 = 34
    16'b11110010_00001000 : OUT <= 30;  //242 / 8 = 30
    16'b11110010_00001001 : OUT <= 26;  //242 / 9 = 26
    16'b11110010_00001010 : OUT <= 24;  //242 / 10 = 24
    16'b11110010_00001011 : OUT <= 22;  //242 / 11 = 22
    16'b11110010_00001100 : OUT <= 20;  //242 / 12 = 20
    16'b11110010_00001101 : OUT <= 18;  //242 / 13 = 18
    16'b11110010_00001110 : OUT <= 17;  //242 / 14 = 17
    16'b11110010_00001111 : OUT <= 16;  //242 / 15 = 16
    16'b11110010_00010000 : OUT <= 15;  //242 / 16 = 15
    16'b11110010_00010001 : OUT <= 14;  //242 / 17 = 14
    16'b11110010_00010010 : OUT <= 13;  //242 / 18 = 13
    16'b11110010_00010011 : OUT <= 12;  //242 / 19 = 12
    16'b11110010_00010100 : OUT <= 12;  //242 / 20 = 12
    16'b11110010_00010101 : OUT <= 11;  //242 / 21 = 11
    16'b11110010_00010110 : OUT <= 11;  //242 / 22 = 11
    16'b11110010_00010111 : OUT <= 10;  //242 / 23 = 10
    16'b11110010_00011000 : OUT <= 10;  //242 / 24 = 10
    16'b11110010_00011001 : OUT <= 9;  //242 / 25 = 9
    16'b11110010_00011010 : OUT <= 9;  //242 / 26 = 9
    16'b11110010_00011011 : OUT <= 8;  //242 / 27 = 8
    16'b11110010_00011100 : OUT <= 8;  //242 / 28 = 8
    16'b11110010_00011101 : OUT <= 8;  //242 / 29 = 8
    16'b11110010_00011110 : OUT <= 8;  //242 / 30 = 8
    16'b11110010_00011111 : OUT <= 7;  //242 / 31 = 7
    16'b11110010_00100000 : OUT <= 7;  //242 / 32 = 7
    16'b11110010_00100001 : OUT <= 7;  //242 / 33 = 7
    16'b11110010_00100010 : OUT <= 7;  //242 / 34 = 7
    16'b11110010_00100011 : OUT <= 6;  //242 / 35 = 6
    16'b11110010_00100100 : OUT <= 6;  //242 / 36 = 6
    16'b11110010_00100101 : OUT <= 6;  //242 / 37 = 6
    16'b11110010_00100110 : OUT <= 6;  //242 / 38 = 6
    16'b11110010_00100111 : OUT <= 6;  //242 / 39 = 6
    16'b11110010_00101000 : OUT <= 6;  //242 / 40 = 6
    16'b11110010_00101001 : OUT <= 5;  //242 / 41 = 5
    16'b11110010_00101010 : OUT <= 5;  //242 / 42 = 5
    16'b11110010_00101011 : OUT <= 5;  //242 / 43 = 5
    16'b11110010_00101100 : OUT <= 5;  //242 / 44 = 5
    16'b11110010_00101101 : OUT <= 5;  //242 / 45 = 5
    16'b11110010_00101110 : OUT <= 5;  //242 / 46 = 5
    16'b11110010_00101111 : OUT <= 5;  //242 / 47 = 5
    16'b11110010_00110000 : OUT <= 5;  //242 / 48 = 5
    16'b11110010_00110001 : OUT <= 4;  //242 / 49 = 4
    16'b11110010_00110010 : OUT <= 4;  //242 / 50 = 4
    16'b11110010_00110011 : OUT <= 4;  //242 / 51 = 4
    16'b11110010_00110100 : OUT <= 4;  //242 / 52 = 4
    16'b11110010_00110101 : OUT <= 4;  //242 / 53 = 4
    16'b11110010_00110110 : OUT <= 4;  //242 / 54 = 4
    16'b11110010_00110111 : OUT <= 4;  //242 / 55 = 4
    16'b11110010_00111000 : OUT <= 4;  //242 / 56 = 4
    16'b11110010_00111001 : OUT <= 4;  //242 / 57 = 4
    16'b11110010_00111010 : OUT <= 4;  //242 / 58 = 4
    16'b11110010_00111011 : OUT <= 4;  //242 / 59 = 4
    16'b11110010_00111100 : OUT <= 4;  //242 / 60 = 4
    16'b11110010_00111101 : OUT <= 3;  //242 / 61 = 3
    16'b11110010_00111110 : OUT <= 3;  //242 / 62 = 3
    16'b11110010_00111111 : OUT <= 3;  //242 / 63 = 3
    16'b11110010_01000000 : OUT <= 3;  //242 / 64 = 3
    16'b11110010_01000001 : OUT <= 3;  //242 / 65 = 3
    16'b11110010_01000010 : OUT <= 3;  //242 / 66 = 3
    16'b11110010_01000011 : OUT <= 3;  //242 / 67 = 3
    16'b11110010_01000100 : OUT <= 3;  //242 / 68 = 3
    16'b11110010_01000101 : OUT <= 3;  //242 / 69 = 3
    16'b11110010_01000110 : OUT <= 3;  //242 / 70 = 3
    16'b11110010_01000111 : OUT <= 3;  //242 / 71 = 3
    16'b11110010_01001000 : OUT <= 3;  //242 / 72 = 3
    16'b11110010_01001001 : OUT <= 3;  //242 / 73 = 3
    16'b11110010_01001010 : OUT <= 3;  //242 / 74 = 3
    16'b11110010_01001011 : OUT <= 3;  //242 / 75 = 3
    16'b11110010_01001100 : OUT <= 3;  //242 / 76 = 3
    16'b11110010_01001101 : OUT <= 3;  //242 / 77 = 3
    16'b11110010_01001110 : OUT <= 3;  //242 / 78 = 3
    16'b11110010_01001111 : OUT <= 3;  //242 / 79 = 3
    16'b11110010_01010000 : OUT <= 3;  //242 / 80 = 3
    16'b11110010_01010001 : OUT <= 2;  //242 / 81 = 2
    16'b11110010_01010010 : OUT <= 2;  //242 / 82 = 2
    16'b11110010_01010011 : OUT <= 2;  //242 / 83 = 2
    16'b11110010_01010100 : OUT <= 2;  //242 / 84 = 2
    16'b11110010_01010101 : OUT <= 2;  //242 / 85 = 2
    16'b11110010_01010110 : OUT <= 2;  //242 / 86 = 2
    16'b11110010_01010111 : OUT <= 2;  //242 / 87 = 2
    16'b11110010_01011000 : OUT <= 2;  //242 / 88 = 2
    16'b11110010_01011001 : OUT <= 2;  //242 / 89 = 2
    16'b11110010_01011010 : OUT <= 2;  //242 / 90 = 2
    16'b11110010_01011011 : OUT <= 2;  //242 / 91 = 2
    16'b11110010_01011100 : OUT <= 2;  //242 / 92 = 2
    16'b11110010_01011101 : OUT <= 2;  //242 / 93 = 2
    16'b11110010_01011110 : OUT <= 2;  //242 / 94 = 2
    16'b11110010_01011111 : OUT <= 2;  //242 / 95 = 2
    16'b11110010_01100000 : OUT <= 2;  //242 / 96 = 2
    16'b11110010_01100001 : OUT <= 2;  //242 / 97 = 2
    16'b11110010_01100010 : OUT <= 2;  //242 / 98 = 2
    16'b11110010_01100011 : OUT <= 2;  //242 / 99 = 2
    16'b11110010_01100100 : OUT <= 2;  //242 / 100 = 2
    16'b11110010_01100101 : OUT <= 2;  //242 / 101 = 2
    16'b11110010_01100110 : OUT <= 2;  //242 / 102 = 2
    16'b11110010_01100111 : OUT <= 2;  //242 / 103 = 2
    16'b11110010_01101000 : OUT <= 2;  //242 / 104 = 2
    16'b11110010_01101001 : OUT <= 2;  //242 / 105 = 2
    16'b11110010_01101010 : OUT <= 2;  //242 / 106 = 2
    16'b11110010_01101011 : OUT <= 2;  //242 / 107 = 2
    16'b11110010_01101100 : OUT <= 2;  //242 / 108 = 2
    16'b11110010_01101101 : OUT <= 2;  //242 / 109 = 2
    16'b11110010_01101110 : OUT <= 2;  //242 / 110 = 2
    16'b11110010_01101111 : OUT <= 2;  //242 / 111 = 2
    16'b11110010_01110000 : OUT <= 2;  //242 / 112 = 2
    16'b11110010_01110001 : OUT <= 2;  //242 / 113 = 2
    16'b11110010_01110010 : OUT <= 2;  //242 / 114 = 2
    16'b11110010_01110011 : OUT <= 2;  //242 / 115 = 2
    16'b11110010_01110100 : OUT <= 2;  //242 / 116 = 2
    16'b11110010_01110101 : OUT <= 2;  //242 / 117 = 2
    16'b11110010_01110110 : OUT <= 2;  //242 / 118 = 2
    16'b11110010_01110111 : OUT <= 2;  //242 / 119 = 2
    16'b11110010_01111000 : OUT <= 2;  //242 / 120 = 2
    16'b11110010_01111001 : OUT <= 2;  //242 / 121 = 2
    16'b11110010_01111010 : OUT <= 1;  //242 / 122 = 1
    16'b11110010_01111011 : OUT <= 1;  //242 / 123 = 1
    16'b11110010_01111100 : OUT <= 1;  //242 / 124 = 1
    16'b11110010_01111101 : OUT <= 1;  //242 / 125 = 1
    16'b11110010_01111110 : OUT <= 1;  //242 / 126 = 1
    16'b11110010_01111111 : OUT <= 1;  //242 / 127 = 1
    16'b11110010_10000000 : OUT <= 1;  //242 / 128 = 1
    16'b11110010_10000001 : OUT <= 1;  //242 / 129 = 1
    16'b11110010_10000010 : OUT <= 1;  //242 / 130 = 1
    16'b11110010_10000011 : OUT <= 1;  //242 / 131 = 1
    16'b11110010_10000100 : OUT <= 1;  //242 / 132 = 1
    16'b11110010_10000101 : OUT <= 1;  //242 / 133 = 1
    16'b11110010_10000110 : OUT <= 1;  //242 / 134 = 1
    16'b11110010_10000111 : OUT <= 1;  //242 / 135 = 1
    16'b11110010_10001000 : OUT <= 1;  //242 / 136 = 1
    16'b11110010_10001001 : OUT <= 1;  //242 / 137 = 1
    16'b11110010_10001010 : OUT <= 1;  //242 / 138 = 1
    16'b11110010_10001011 : OUT <= 1;  //242 / 139 = 1
    16'b11110010_10001100 : OUT <= 1;  //242 / 140 = 1
    16'b11110010_10001101 : OUT <= 1;  //242 / 141 = 1
    16'b11110010_10001110 : OUT <= 1;  //242 / 142 = 1
    16'b11110010_10001111 : OUT <= 1;  //242 / 143 = 1
    16'b11110010_10010000 : OUT <= 1;  //242 / 144 = 1
    16'b11110010_10010001 : OUT <= 1;  //242 / 145 = 1
    16'b11110010_10010010 : OUT <= 1;  //242 / 146 = 1
    16'b11110010_10010011 : OUT <= 1;  //242 / 147 = 1
    16'b11110010_10010100 : OUT <= 1;  //242 / 148 = 1
    16'b11110010_10010101 : OUT <= 1;  //242 / 149 = 1
    16'b11110010_10010110 : OUT <= 1;  //242 / 150 = 1
    16'b11110010_10010111 : OUT <= 1;  //242 / 151 = 1
    16'b11110010_10011000 : OUT <= 1;  //242 / 152 = 1
    16'b11110010_10011001 : OUT <= 1;  //242 / 153 = 1
    16'b11110010_10011010 : OUT <= 1;  //242 / 154 = 1
    16'b11110010_10011011 : OUT <= 1;  //242 / 155 = 1
    16'b11110010_10011100 : OUT <= 1;  //242 / 156 = 1
    16'b11110010_10011101 : OUT <= 1;  //242 / 157 = 1
    16'b11110010_10011110 : OUT <= 1;  //242 / 158 = 1
    16'b11110010_10011111 : OUT <= 1;  //242 / 159 = 1
    16'b11110010_10100000 : OUT <= 1;  //242 / 160 = 1
    16'b11110010_10100001 : OUT <= 1;  //242 / 161 = 1
    16'b11110010_10100010 : OUT <= 1;  //242 / 162 = 1
    16'b11110010_10100011 : OUT <= 1;  //242 / 163 = 1
    16'b11110010_10100100 : OUT <= 1;  //242 / 164 = 1
    16'b11110010_10100101 : OUT <= 1;  //242 / 165 = 1
    16'b11110010_10100110 : OUT <= 1;  //242 / 166 = 1
    16'b11110010_10100111 : OUT <= 1;  //242 / 167 = 1
    16'b11110010_10101000 : OUT <= 1;  //242 / 168 = 1
    16'b11110010_10101001 : OUT <= 1;  //242 / 169 = 1
    16'b11110010_10101010 : OUT <= 1;  //242 / 170 = 1
    16'b11110010_10101011 : OUT <= 1;  //242 / 171 = 1
    16'b11110010_10101100 : OUT <= 1;  //242 / 172 = 1
    16'b11110010_10101101 : OUT <= 1;  //242 / 173 = 1
    16'b11110010_10101110 : OUT <= 1;  //242 / 174 = 1
    16'b11110010_10101111 : OUT <= 1;  //242 / 175 = 1
    16'b11110010_10110000 : OUT <= 1;  //242 / 176 = 1
    16'b11110010_10110001 : OUT <= 1;  //242 / 177 = 1
    16'b11110010_10110010 : OUT <= 1;  //242 / 178 = 1
    16'b11110010_10110011 : OUT <= 1;  //242 / 179 = 1
    16'b11110010_10110100 : OUT <= 1;  //242 / 180 = 1
    16'b11110010_10110101 : OUT <= 1;  //242 / 181 = 1
    16'b11110010_10110110 : OUT <= 1;  //242 / 182 = 1
    16'b11110010_10110111 : OUT <= 1;  //242 / 183 = 1
    16'b11110010_10111000 : OUT <= 1;  //242 / 184 = 1
    16'b11110010_10111001 : OUT <= 1;  //242 / 185 = 1
    16'b11110010_10111010 : OUT <= 1;  //242 / 186 = 1
    16'b11110010_10111011 : OUT <= 1;  //242 / 187 = 1
    16'b11110010_10111100 : OUT <= 1;  //242 / 188 = 1
    16'b11110010_10111101 : OUT <= 1;  //242 / 189 = 1
    16'b11110010_10111110 : OUT <= 1;  //242 / 190 = 1
    16'b11110010_10111111 : OUT <= 1;  //242 / 191 = 1
    16'b11110010_11000000 : OUT <= 1;  //242 / 192 = 1
    16'b11110010_11000001 : OUT <= 1;  //242 / 193 = 1
    16'b11110010_11000010 : OUT <= 1;  //242 / 194 = 1
    16'b11110010_11000011 : OUT <= 1;  //242 / 195 = 1
    16'b11110010_11000100 : OUT <= 1;  //242 / 196 = 1
    16'b11110010_11000101 : OUT <= 1;  //242 / 197 = 1
    16'b11110010_11000110 : OUT <= 1;  //242 / 198 = 1
    16'b11110010_11000111 : OUT <= 1;  //242 / 199 = 1
    16'b11110010_11001000 : OUT <= 1;  //242 / 200 = 1
    16'b11110010_11001001 : OUT <= 1;  //242 / 201 = 1
    16'b11110010_11001010 : OUT <= 1;  //242 / 202 = 1
    16'b11110010_11001011 : OUT <= 1;  //242 / 203 = 1
    16'b11110010_11001100 : OUT <= 1;  //242 / 204 = 1
    16'b11110010_11001101 : OUT <= 1;  //242 / 205 = 1
    16'b11110010_11001110 : OUT <= 1;  //242 / 206 = 1
    16'b11110010_11001111 : OUT <= 1;  //242 / 207 = 1
    16'b11110010_11010000 : OUT <= 1;  //242 / 208 = 1
    16'b11110010_11010001 : OUT <= 1;  //242 / 209 = 1
    16'b11110010_11010010 : OUT <= 1;  //242 / 210 = 1
    16'b11110010_11010011 : OUT <= 1;  //242 / 211 = 1
    16'b11110010_11010100 : OUT <= 1;  //242 / 212 = 1
    16'b11110010_11010101 : OUT <= 1;  //242 / 213 = 1
    16'b11110010_11010110 : OUT <= 1;  //242 / 214 = 1
    16'b11110010_11010111 : OUT <= 1;  //242 / 215 = 1
    16'b11110010_11011000 : OUT <= 1;  //242 / 216 = 1
    16'b11110010_11011001 : OUT <= 1;  //242 / 217 = 1
    16'b11110010_11011010 : OUT <= 1;  //242 / 218 = 1
    16'b11110010_11011011 : OUT <= 1;  //242 / 219 = 1
    16'b11110010_11011100 : OUT <= 1;  //242 / 220 = 1
    16'b11110010_11011101 : OUT <= 1;  //242 / 221 = 1
    16'b11110010_11011110 : OUT <= 1;  //242 / 222 = 1
    16'b11110010_11011111 : OUT <= 1;  //242 / 223 = 1
    16'b11110010_11100000 : OUT <= 1;  //242 / 224 = 1
    16'b11110010_11100001 : OUT <= 1;  //242 / 225 = 1
    16'b11110010_11100010 : OUT <= 1;  //242 / 226 = 1
    16'b11110010_11100011 : OUT <= 1;  //242 / 227 = 1
    16'b11110010_11100100 : OUT <= 1;  //242 / 228 = 1
    16'b11110010_11100101 : OUT <= 1;  //242 / 229 = 1
    16'b11110010_11100110 : OUT <= 1;  //242 / 230 = 1
    16'b11110010_11100111 : OUT <= 1;  //242 / 231 = 1
    16'b11110010_11101000 : OUT <= 1;  //242 / 232 = 1
    16'b11110010_11101001 : OUT <= 1;  //242 / 233 = 1
    16'b11110010_11101010 : OUT <= 1;  //242 / 234 = 1
    16'b11110010_11101011 : OUT <= 1;  //242 / 235 = 1
    16'b11110010_11101100 : OUT <= 1;  //242 / 236 = 1
    16'b11110010_11101101 : OUT <= 1;  //242 / 237 = 1
    16'b11110010_11101110 : OUT <= 1;  //242 / 238 = 1
    16'b11110010_11101111 : OUT <= 1;  //242 / 239 = 1
    16'b11110010_11110000 : OUT <= 1;  //242 / 240 = 1
    16'b11110010_11110001 : OUT <= 1;  //242 / 241 = 1
    16'b11110010_11110010 : OUT <= 1;  //242 / 242 = 1
    16'b11110010_11110011 : OUT <= 0;  //242 / 243 = 0
    16'b11110010_11110100 : OUT <= 0;  //242 / 244 = 0
    16'b11110010_11110101 : OUT <= 0;  //242 / 245 = 0
    16'b11110010_11110110 : OUT <= 0;  //242 / 246 = 0
    16'b11110010_11110111 : OUT <= 0;  //242 / 247 = 0
    16'b11110010_11111000 : OUT <= 0;  //242 / 248 = 0
    16'b11110010_11111001 : OUT <= 0;  //242 / 249 = 0
    16'b11110010_11111010 : OUT <= 0;  //242 / 250 = 0
    16'b11110010_11111011 : OUT <= 0;  //242 / 251 = 0
    16'b11110010_11111100 : OUT <= 0;  //242 / 252 = 0
    16'b11110010_11111101 : OUT <= 0;  //242 / 253 = 0
    16'b11110010_11111110 : OUT <= 0;  //242 / 254 = 0
    16'b11110010_11111111 : OUT <= 0;  //242 / 255 = 0
    16'b11110011_00000000 : OUT <= 0;  //243 / 0 = 0
    16'b11110011_00000001 : OUT <= 243;  //243 / 1 = 243
    16'b11110011_00000010 : OUT <= 121;  //243 / 2 = 121
    16'b11110011_00000011 : OUT <= 81;  //243 / 3 = 81
    16'b11110011_00000100 : OUT <= 60;  //243 / 4 = 60
    16'b11110011_00000101 : OUT <= 48;  //243 / 5 = 48
    16'b11110011_00000110 : OUT <= 40;  //243 / 6 = 40
    16'b11110011_00000111 : OUT <= 34;  //243 / 7 = 34
    16'b11110011_00001000 : OUT <= 30;  //243 / 8 = 30
    16'b11110011_00001001 : OUT <= 27;  //243 / 9 = 27
    16'b11110011_00001010 : OUT <= 24;  //243 / 10 = 24
    16'b11110011_00001011 : OUT <= 22;  //243 / 11 = 22
    16'b11110011_00001100 : OUT <= 20;  //243 / 12 = 20
    16'b11110011_00001101 : OUT <= 18;  //243 / 13 = 18
    16'b11110011_00001110 : OUT <= 17;  //243 / 14 = 17
    16'b11110011_00001111 : OUT <= 16;  //243 / 15 = 16
    16'b11110011_00010000 : OUT <= 15;  //243 / 16 = 15
    16'b11110011_00010001 : OUT <= 14;  //243 / 17 = 14
    16'b11110011_00010010 : OUT <= 13;  //243 / 18 = 13
    16'b11110011_00010011 : OUT <= 12;  //243 / 19 = 12
    16'b11110011_00010100 : OUT <= 12;  //243 / 20 = 12
    16'b11110011_00010101 : OUT <= 11;  //243 / 21 = 11
    16'b11110011_00010110 : OUT <= 11;  //243 / 22 = 11
    16'b11110011_00010111 : OUT <= 10;  //243 / 23 = 10
    16'b11110011_00011000 : OUT <= 10;  //243 / 24 = 10
    16'b11110011_00011001 : OUT <= 9;  //243 / 25 = 9
    16'b11110011_00011010 : OUT <= 9;  //243 / 26 = 9
    16'b11110011_00011011 : OUT <= 9;  //243 / 27 = 9
    16'b11110011_00011100 : OUT <= 8;  //243 / 28 = 8
    16'b11110011_00011101 : OUT <= 8;  //243 / 29 = 8
    16'b11110011_00011110 : OUT <= 8;  //243 / 30 = 8
    16'b11110011_00011111 : OUT <= 7;  //243 / 31 = 7
    16'b11110011_00100000 : OUT <= 7;  //243 / 32 = 7
    16'b11110011_00100001 : OUT <= 7;  //243 / 33 = 7
    16'b11110011_00100010 : OUT <= 7;  //243 / 34 = 7
    16'b11110011_00100011 : OUT <= 6;  //243 / 35 = 6
    16'b11110011_00100100 : OUT <= 6;  //243 / 36 = 6
    16'b11110011_00100101 : OUT <= 6;  //243 / 37 = 6
    16'b11110011_00100110 : OUT <= 6;  //243 / 38 = 6
    16'b11110011_00100111 : OUT <= 6;  //243 / 39 = 6
    16'b11110011_00101000 : OUT <= 6;  //243 / 40 = 6
    16'b11110011_00101001 : OUT <= 5;  //243 / 41 = 5
    16'b11110011_00101010 : OUT <= 5;  //243 / 42 = 5
    16'b11110011_00101011 : OUT <= 5;  //243 / 43 = 5
    16'b11110011_00101100 : OUT <= 5;  //243 / 44 = 5
    16'b11110011_00101101 : OUT <= 5;  //243 / 45 = 5
    16'b11110011_00101110 : OUT <= 5;  //243 / 46 = 5
    16'b11110011_00101111 : OUT <= 5;  //243 / 47 = 5
    16'b11110011_00110000 : OUT <= 5;  //243 / 48 = 5
    16'b11110011_00110001 : OUT <= 4;  //243 / 49 = 4
    16'b11110011_00110010 : OUT <= 4;  //243 / 50 = 4
    16'b11110011_00110011 : OUT <= 4;  //243 / 51 = 4
    16'b11110011_00110100 : OUT <= 4;  //243 / 52 = 4
    16'b11110011_00110101 : OUT <= 4;  //243 / 53 = 4
    16'b11110011_00110110 : OUT <= 4;  //243 / 54 = 4
    16'b11110011_00110111 : OUT <= 4;  //243 / 55 = 4
    16'b11110011_00111000 : OUT <= 4;  //243 / 56 = 4
    16'b11110011_00111001 : OUT <= 4;  //243 / 57 = 4
    16'b11110011_00111010 : OUT <= 4;  //243 / 58 = 4
    16'b11110011_00111011 : OUT <= 4;  //243 / 59 = 4
    16'b11110011_00111100 : OUT <= 4;  //243 / 60 = 4
    16'b11110011_00111101 : OUT <= 3;  //243 / 61 = 3
    16'b11110011_00111110 : OUT <= 3;  //243 / 62 = 3
    16'b11110011_00111111 : OUT <= 3;  //243 / 63 = 3
    16'b11110011_01000000 : OUT <= 3;  //243 / 64 = 3
    16'b11110011_01000001 : OUT <= 3;  //243 / 65 = 3
    16'b11110011_01000010 : OUT <= 3;  //243 / 66 = 3
    16'b11110011_01000011 : OUT <= 3;  //243 / 67 = 3
    16'b11110011_01000100 : OUT <= 3;  //243 / 68 = 3
    16'b11110011_01000101 : OUT <= 3;  //243 / 69 = 3
    16'b11110011_01000110 : OUT <= 3;  //243 / 70 = 3
    16'b11110011_01000111 : OUT <= 3;  //243 / 71 = 3
    16'b11110011_01001000 : OUT <= 3;  //243 / 72 = 3
    16'b11110011_01001001 : OUT <= 3;  //243 / 73 = 3
    16'b11110011_01001010 : OUT <= 3;  //243 / 74 = 3
    16'b11110011_01001011 : OUT <= 3;  //243 / 75 = 3
    16'b11110011_01001100 : OUT <= 3;  //243 / 76 = 3
    16'b11110011_01001101 : OUT <= 3;  //243 / 77 = 3
    16'b11110011_01001110 : OUT <= 3;  //243 / 78 = 3
    16'b11110011_01001111 : OUT <= 3;  //243 / 79 = 3
    16'b11110011_01010000 : OUT <= 3;  //243 / 80 = 3
    16'b11110011_01010001 : OUT <= 3;  //243 / 81 = 3
    16'b11110011_01010010 : OUT <= 2;  //243 / 82 = 2
    16'b11110011_01010011 : OUT <= 2;  //243 / 83 = 2
    16'b11110011_01010100 : OUT <= 2;  //243 / 84 = 2
    16'b11110011_01010101 : OUT <= 2;  //243 / 85 = 2
    16'b11110011_01010110 : OUT <= 2;  //243 / 86 = 2
    16'b11110011_01010111 : OUT <= 2;  //243 / 87 = 2
    16'b11110011_01011000 : OUT <= 2;  //243 / 88 = 2
    16'b11110011_01011001 : OUT <= 2;  //243 / 89 = 2
    16'b11110011_01011010 : OUT <= 2;  //243 / 90 = 2
    16'b11110011_01011011 : OUT <= 2;  //243 / 91 = 2
    16'b11110011_01011100 : OUT <= 2;  //243 / 92 = 2
    16'b11110011_01011101 : OUT <= 2;  //243 / 93 = 2
    16'b11110011_01011110 : OUT <= 2;  //243 / 94 = 2
    16'b11110011_01011111 : OUT <= 2;  //243 / 95 = 2
    16'b11110011_01100000 : OUT <= 2;  //243 / 96 = 2
    16'b11110011_01100001 : OUT <= 2;  //243 / 97 = 2
    16'b11110011_01100010 : OUT <= 2;  //243 / 98 = 2
    16'b11110011_01100011 : OUT <= 2;  //243 / 99 = 2
    16'b11110011_01100100 : OUT <= 2;  //243 / 100 = 2
    16'b11110011_01100101 : OUT <= 2;  //243 / 101 = 2
    16'b11110011_01100110 : OUT <= 2;  //243 / 102 = 2
    16'b11110011_01100111 : OUT <= 2;  //243 / 103 = 2
    16'b11110011_01101000 : OUT <= 2;  //243 / 104 = 2
    16'b11110011_01101001 : OUT <= 2;  //243 / 105 = 2
    16'b11110011_01101010 : OUT <= 2;  //243 / 106 = 2
    16'b11110011_01101011 : OUT <= 2;  //243 / 107 = 2
    16'b11110011_01101100 : OUT <= 2;  //243 / 108 = 2
    16'b11110011_01101101 : OUT <= 2;  //243 / 109 = 2
    16'b11110011_01101110 : OUT <= 2;  //243 / 110 = 2
    16'b11110011_01101111 : OUT <= 2;  //243 / 111 = 2
    16'b11110011_01110000 : OUT <= 2;  //243 / 112 = 2
    16'b11110011_01110001 : OUT <= 2;  //243 / 113 = 2
    16'b11110011_01110010 : OUT <= 2;  //243 / 114 = 2
    16'b11110011_01110011 : OUT <= 2;  //243 / 115 = 2
    16'b11110011_01110100 : OUT <= 2;  //243 / 116 = 2
    16'b11110011_01110101 : OUT <= 2;  //243 / 117 = 2
    16'b11110011_01110110 : OUT <= 2;  //243 / 118 = 2
    16'b11110011_01110111 : OUT <= 2;  //243 / 119 = 2
    16'b11110011_01111000 : OUT <= 2;  //243 / 120 = 2
    16'b11110011_01111001 : OUT <= 2;  //243 / 121 = 2
    16'b11110011_01111010 : OUT <= 1;  //243 / 122 = 1
    16'b11110011_01111011 : OUT <= 1;  //243 / 123 = 1
    16'b11110011_01111100 : OUT <= 1;  //243 / 124 = 1
    16'b11110011_01111101 : OUT <= 1;  //243 / 125 = 1
    16'b11110011_01111110 : OUT <= 1;  //243 / 126 = 1
    16'b11110011_01111111 : OUT <= 1;  //243 / 127 = 1
    16'b11110011_10000000 : OUT <= 1;  //243 / 128 = 1
    16'b11110011_10000001 : OUT <= 1;  //243 / 129 = 1
    16'b11110011_10000010 : OUT <= 1;  //243 / 130 = 1
    16'b11110011_10000011 : OUT <= 1;  //243 / 131 = 1
    16'b11110011_10000100 : OUT <= 1;  //243 / 132 = 1
    16'b11110011_10000101 : OUT <= 1;  //243 / 133 = 1
    16'b11110011_10000110 : OUT <= 1;  //243 / 134 = 1
    16'b11110011_10000111 : OUT <= 1;  //243 / 135 = 1
    16'b11110011_10001000 : OUT <= 1;  //243 / 136 = 1
    16'b11110011_10001001 : OUT <= 1;  //243 / 137 = 1
    16'b11110011_10001010 : OUT <= 1;  //243 / 138 = 1
    16'b11110011_10001011 : OUT <= 1;  //243 / 139 = 1
    16'b11110011_10001100 : OUT <= 1;  //243 / 140 = 1
    16'b11110011_10001101 : OUT <= 1;  //243 / 141 = 1
    16'b11110011_10001110 : OUT <= 1;  //243 / 142 = 1
    16'b11110011_10001111 : OUT <= 1;  //243 / 143 = 1
    16'b11110011_10010000 : OUT <= 1;  //243 / 144 = 1
    16'b11110011_10010001 : OUT <= 1;  //243 / 145 = 1
    16'b11110011_10010010 : OUT <= 1;  //243 / 146 = 1
    16'b11110011_10010011 : OUT <= 1;  //243 / 147 = 1
    16'b11110011_10010100 : OUT <= 1;  //243 / 148 = 1
    16'b11110011_10010101 : OUT <= 1;  //243 / 149 = 1
    16'b11110011_10010110 : OUT <= 1;  //243 / 150 = 1
    16'b11110011_10010111 : OUT <= 1;  //243 / 151 = 1
    16'b11110011_10011000 : OUT <= 1;  //243 / 152 = 1
    16'b11110011_10011001 : OUT <= 1;  //243 / 153 = 1
    16'b11110011_10011010 : OUT <= 1;  //243 / 154 = 1
    16'b11110011_10011011 : OUT <= 1;  //243 / 155 = 1
    16'b11110011_10011100 : OUT <= 1;  //243 / 156 = 1
    16'b11110011_10011101 : OUT <= 1;  //243 / 157 = 1
    16'b11110011_10011110 : OUT <= 1;  //243 / 158 = 1
    16'b11110011_10011111 : OUT <= 1;  //243 / 159 = 1
    16'b11110011_10100000 : OUT <= 1;  //243 / 160 = 1
    16'b11110011_10100001 : OUT <= 1;  //243 / 161 = 1
    16'b11110011_10100010 : OUT <= 1;  //243 / 162 = 1
    16'b11110011_10100011 : OUT <= 1;  //243 / 163 = 1
    16'b11110011_10100100 : OUT <= 1;  //243 / 164 = 1
    16'b11110011_10100101 : OUT <= 1;  //243 / 165 = 1
    16'b11110011_10100110 : OUT <= 1;  //243 / 166 = 1
    16'b11110011_10100111 : OUT <= 1;  //243 / 167 = 1
    16'b11110011_10101000 : OUT <= 1;  //243 / 168 = 1
    16'b11110011_10101001 : OUT <= 1;  //243 / 169 = 1
    16'b11110011_10101010 : OUT <= 1;  //243 / 170 = 1
    16'b11110011_10101011 : OUT <= 1;  //243 / 171 = 1
    16'b11110011_10101100 : OUT <= 1;  //243 / 172 = 1
    16'b11110011_10101101 : OUT <= 1;  //243 / 173 = 1
    16'b11110011_10101110 : OUT <= 1;  //243 / 174 = 1
    16'b11110011_10101111 : OUT <= 1;  //243 / 175 = 1
    16'b11110011_10110000 : OUT <= 1;  //243 / 176 = 1
    16'b11110011_10110001 : OUT <= 1;  //243 / 177 = 1
    16'b11110011_10110010 : OUT <= 1;  //243 / 178 = 1
    16'b11110011_10110011 : OUT <= 1;  //243 / 179 = 1
    16'b11110011_10110100 : OUT <= 1;  //243 / 180 = 1
    16'b11110011_10110101 : OUT <= 1;  //243 / 181 = 1
    16'b11110011_10110110 : OUT <= 1;  //243 / 182 = 1
    16'b11110011_10110111 : OUT <= 1;  //243 / 183 = 1
    16'b11110011_10111000 : OUT <= 1;  //243 / 184 = 1
    16'b11110011_10111001 : OUT <= 1;  //243 / 185 = 1
    16'b11110011_10111010 : OUT <= 1;  //243 / 186 = 1
    16'b11110011_10111011 : OUT <= 1;  //243 / 187 = 1
    16'b11110011_10111100 : OUT <= 1;  //243 / 188 = 1
    16'b11110011_10111101 : OUT <= 1;  //243 / 189 = 1
    16'b11110011_10111110 : OUT <= 1;  //243 / 190 = 1
    16'b11110011_10111111 : OUT <= 1;  //243 / 191 = 1
    16'b11110011_11000000 : OUT <= 1;  //243 / 192 = 1
    16'b11110011_11000001 : OUT <= 1;  //243 / 193 = 1
    16'b11110011_11000010 : OUT <= 1;  //243 / 194 = 1
    16'b11110011_11000011 : OUT <= 1;  //243 / 195 = 1
    16'b11110011_11000100 : OUT <= 1;  //243 / 196 = 1
    16'b11110011_11000101 : OUT <= 1;  //243 / 197 = 1
    16'b11110011_11000110 : OUT <= 1;  //243 / 198 = 1
    16'b11110011_11000111 : OUT <= 1;  //243 / 199 = 1
    16'b11110011_11001000 : OUT <= 1;  //243 / 200 = 1
    16'b11110011_11001001 : OUT <= 1;  //243 / 201 = 1
    16'b11110011_11001010 : OUT <= 1;  //243 / 202 = 1
    16'b11110011_11001011 : OUT <= 1;  //243 / 203 = 1
    16'b11110011_11001100 : OUT <= 1;  //243 / 204 = 1
    16'b11110011_11001101 : OUT <= 1;  //243 / 205 = 1
    16'b11110011_11001110 : OUT <= 1;  //243 / 206 = 1
    16'b11110011_11001111 : OUT <= 1;  //243 / 207 = 1
    16'b11110011_11010000 : OUT <= 1;  //243 / 208 = 1
    16'b11110011_11010001 : OUT <= 1;  //243 / 209 = 1
    16'b11110011_11010010 : OUT <= 1;  //243 / 210 = 1
    16'b11110011_11010011 : OUT <= 1;  //243 / 211 = 1
    16'b11110011_11010100 : OUT <= 1;  //243 / 212 = 1
    16'b11110011_11010101 : OUT <= 1;  //243 / 213 = 1
    16'b11110011_11010110 : OUT <= 1;  //243 / 214 = 1
    16'b11110011_11010111 : OUT <= 1;  //243 / 215 = 1
    16'b11110011_11011000 : OUT <= 1;  //243 / 216 = 1
    16'b11110011_11011001 : OUT <= 1;  //243 / 217 = 1
    16'b11110011_11011010 : OUT <= 1;  //243 / 218 = 1
    16'b11110011_11011011 : OUT <= 1;  //243 / 219 = 1
    16'b11110011_11011100 : OUT <= 1;  //243 / 220 = 1
    16'b11110011_11011101 : OUT <= 1;  //243 / 221 = 1
    16'b11110011_11011110 : OUT <= 1;  //243 / 222 = 1
    16'b11110011_11011111 : OUT <= 1;  //243 / 223 = 1
    16'b11110011_11100000 : OUT <= 1;  //243 / 224 = 1
    16'b11110011_11100001 : OUT <= 1;  //243 / 225 = 1
    16'b11110011_11100010 : OUT <= 1;  //243 / 226 = 1
    16'b11110011_11100011 : OUT <= 1;  //243 / 227 = 1
    16'b11110011_11100100 : OUT <= 1;  //243 / 228 = 1
    16'b11110011_11100101 : OUT <= 1;  //243 / 229 = 1
    16'b11110011_11100110 : OUT <= 1;  //243 / 230 = 1
    16'b11110011_11100111 : OUT <= 1;  //243 / 231 = 1
    16'b11110011_11101000 : OUT <= 1;  //243 / 232 = 1
    16'b11110011_11101001 : OUT <= 1;  //243 / 233 = 1
    16'b11110011_11101010 : OUT <= 1;  //243 / 234 = 1
    16'b11110011_11101011 : OUT <= 1;  //243 / 235 = 1
    16'b11110011_11101100 : OUT <= 1;  //243 / 236 = 1
    16'b11110011_11101101 : OUT <= 1;  //243 / 237 = 1
    16'b11110011_11101110 : OUT <= 1;  //243 / 238 = 1
    16'b11110011_11101111 : OUT <= 1;  //243 / 239 = 1
    16'b11110011_11110000 : OUT <= 1;  //243 / 240 = 1
    16'b11110011_11110001 : OUT <= 1;  //243 / 241 = 1
    16'b11110011_11110010 : OUT <= 1;  //243 / 242 = 1
    16'b11110011_11110011 : OUT <= 1;  //243 / 243 = 1
    16'b11110011_11110100 : OUT <= 0;  //243 / 244 = 0
    16'b11110011_11110101 : OUT <= 0;  //243 / 245 = 0
    16'b11110011_11110110 : OUT <= 0;  //243 / 246 = 0
    16'b11110011_11110111 : OUT <= 0;  //243 / 247 = 0
    16'b11110011_11111000 : OUT <= 0;  //243 / 248 = 0
    16'b11110011_11111001 : OUT <= 0;  //243 / 249 = 0
    16'b11110011_11111010 : OUT <= 0;  //243 / 250 = 0
    16'b11110011_11111011 : OUT <= 0;  //243 / 251 = 0
    16'b11110011_11111100 : OUT <= 0;  //243 / 252 = 0
    16'b11110011_11111101 : OUT <= 0;  //243 / 253 = 0
    16'b11110011_11111110 : OUT <= 0;  //243 / 254 = 0
    16'b11110011_11111111 : OUT <= 0;  //243 / 255 = 0
    16'b11110100_00000000 : OUT <= 0;  //244 / 0 = 0
    16'b11110100_00000001 : OUT <= 244;  //244 / 1 = 244
    16'b11110100_00000010 : OUT <= 122;  //244 / 2 = 122
    16'b11110100_00000011 : OUT <= 81;  //244 / 3 = 81
    16'b11110100_00000100 : OUT <= 61;  //244 / 4 = 61
    16'b11110100_00000101 : OUT <= 48;  //244 / 5 = 48
    16'b11110100_00000110 : OUT <= 40;  //244 / 6 = 40
    16'b11110100_00000111 : OUT <= 34;  //244 / 7 = 34
    16'b11110100_00001000 : OUT <= 30;  //244 / 8 = 30
    16'b11110100_00001001 : OUT <= 27;  //244 / 9 = 27
    16'b11110100_00001010 : OUT <= 24;  //244 / 10 = 24
    16'b11110100_00001011 : OUT <= 22;  //244 / 11 = 22
    16'b11110100_00001100 : OUT <= 20;  //244 / 12 = 20
    16'b11110100_00001101 : OUT <= 18;  //244 / 13 = 18
    16'b11110100_00001110 : OUT <= 17;  //244 / 14 = 17
    16'b11110100_00001111 : OUT <= 16;  //244 / 15 = 16
    16'b11110100_00010000 : OUT <= 15;  //244 / 16 = 15
    16'b11110100_00010001 : OUT <= 14;  //244 / 17 = 14
    16'b11110100_00010010 : OUT <= 13;  //244 / 18 = 13
    16'b11110100_00010011 : OUT <= 12;  //244 / 19 = 12
    16'b11110100_00010100 : OUT <= 12;  //244 / 20 = 12
    16'b11110100_00010101 : OUT <= 11;  //244 / 21 = 11
    16'b11110100_00010110 : OUT <= 11;  //244 / 22 = 11
    16'b11110100_00010111 : OUT <= 10;  //244 / 23 = 10
    16'b11110100_00011000 : OUT <= 10;  //244 / 24 = 10
    16'b11110100_00011001 : OUT <= 9;  //244 / 25 = 9
    16'b11110100_00011010 : OUT <= 9;  //244 / 26 = 9
    16'b11110100_00011011 : OUT <= 9;  //244 / 27 = 9
    16'b11110100_00011100 : OUT <= 8;  //244 / 28 = 8
    16'b11110100_00011101 : OUT <= 8;  //244 / 29 = 8
    16'b11110100_00011110 : OUT <= 8;  //244 / 30 = 8
    16'b11110100_00011111 : OUT <= 7;  //244 / 31 = 7
    16'b11110100_00100000 : OUT <= 7;  //244 / 32 = 7
    16'b11110100_00100001 : OUT <= 7;  //244 / 33 = 7
    16'b11110100_00100010 : OUT <= 7;  //244 / 34 = 7
    16'b11110100_00100011 : OUT <= 6;  //244 / 35 = 6
    16'b11110100_00100100 : OUT <= 6;  //244 / 36 = 6
    16'b11110100_00100101 : OUT <= 6;  //244 / 37 = 6
    16'b11110100_00100110 : OUT <= 6;  //244 / 38 = 6
    16'b11110100_00100111 : OUT <= 6;  //244 / 39 = 6
    16'b11110100_00101000 : OUT <= 6;  //244 / 40 = 6
    16'b11110100_00101001 : OUT <= 5;  //244 / 41 = 5
    16'b11110100_00101010 : OUT <= 5;  //244 / 42 = 5
    16'b11110100_00101011 : OUT <= 5;  //244 / 43 = 5
    16'b11110100_00101100 : OUT <= 5;  //244 / 44 = 5
    16'b11110100_00101101 : OUT <= 5;  //244 / 45 = 5
    16'b11110100_00101110 : OUT <= 5;  //244 / 46 = 5
    16'b11110100_00101111 : OUT <= 5;  //244 / 47 = 5
    16'b11110100_00110000 : OUT <= 5;  //244 / 48 = 5
    16'b11110100_00110001 : OUT <= 4;  //244 / 49 = 4
    16'b11110100_00110010 : OUT <= 4;  //244 / 50 = 4
    16'b11110100_00110011 : OUT <= 4;  //244 / 51 = 4
    16'b11110100_00110100 : OUT <= 4;  //244 / 52 = 4
    16'b11110100_00110101 : OUT <= 4;  //244 / 53 = 4
    16'b11110100_00110110 : OUT <= 4;  //244 / 54 = 4
    16'b11110100_00110111 : OUT <= 4;  //244 / 55 = 4
    16'b11110100_00111000 : OUT <= 4;  //244 / 56 = 4
    16'b11110100_00111001 : OUT <= 4;  //244 / 57 = 4
    16'b11110100_00111010 : OUT <= 4;  //244 / 58 = 4
    16'b11110100_00111011 : OUT <= 4;  //244 / 59 = 4
    16'b11110100_00111100 : OUT <= 4;  //244 / 60 = 4
    16'b11110100_00111101 : OUT <= 4;  //244 / 61 = 4
    16'b11110100_00111110 : OUT <= 3;  //244 / 62 = 3
    16'b11110100_00111111 : OUT <= 3;  //244 / 63 = 3
    16'b11110100_01000000 : OUT <= 3;  //244 / 64 = 3
    16'b11110100_01000001 : OUT <= 3;  //244 / 65 = 3
    16'b11110100_01000010 : OUT <= 3;  //244 / 66 = 3
    16'b11110100_01000011 : OUT <= 3;  //244 / 67 = 3
    16'b11110100_01000100 : OUT <= 3;  //244 / 68 = 3
    16'b11110100_01000101 : OUT <= 3;  //244 / 69 = 3
    16'b11110100_01000110 : OUT <= 3;  //244 / 70 = 3
    16'b11110100_01000111 : OUT <= 3;  //244 / 71 = 3
    16'b11110100_01001000 : OUT <= 3;  //244 / 72 = 3
    16'b11110100_01001001 : OUT <= 3;  //244 / 73 = 3
    16'b11110100_01001010 : OUT <= 3;  //244 / 74 = 3
    16'b11110100_01001011 : OUT <= 3;  //244 / 75 = 3
    16'b11110100_01001100 : OUT <= 3;  //244 / 76 = 3
    16'b11110100_01001101 : OUT <= 3;  //244 / 77 = 3
    16'b11110100_01001110 : OUT <= 3;  //244 / 78 = 3
    16'b11110100_01001111 : OUT <= 3;  //244 / 79 = 3
    16'b11110100_01010000 : OUT <= 3;  //244 / 80 = 3
    16'b11110100_01010001 : OUT <= 3;  //244 / 81 = 3
    16'b11110100_01010010 : OUT <= 2;  //244 / 82 = 2
    16'b11110100_01010011 : OUT <= 2;  //244 / 83 = 2
    16'b11110100_01010100 : OUT <= 2;  //244 / 84 = 2
    16'b11110100_01010101 : OUT <= 2;  //244 / 85 = 2
    16'b11110100_01010110 : OUT <= 2;  //244 / 86 = 2
    16'b11110100_01010111 : OUT <= 2;  //244 / 87 = 2
    16'b11110100_01011000 : OUT <= 2;  //244 / 88 = 2
    16'b11110100_01011001 : OUT <= 2;  //244 / 89 = 2
    16'b11110100_01011010 : OUT <= 2;  //244 / 90 = 2
    16'b11110100_01011011 : OUT <= 2;  //244 / 91 = 2
    16'b11110100_01011100 : OUT <= 2;  //244 / 92 = 2
    16'b11110100_01011101 : OUT <= 2;  //244 / 93 = 2
    16'b11110100_01011110 : OUT <= 2;  //244 / 94 = 2
    16'b11110100_01011111 : OUT <= 2;  //244 / 95 = 2
    16'b11110100_01100000 : OUT <= 2;  //244 / 96 = 2
    16'b11110100_01100001 : OUT <= 2;  //244 / 97 = 2
    16'b11110100_01100010 : OUT <= 2;  //244 / 98 = 2
    16'b11110100_01100011 : OUT <= 2;  //244 / 99 = 2
    16'b11110100_01100100 : OUT <= 2;  //244 / 100 = 2
    16'b11110100_01100101 : OUT <= 2;  //244 / 101 = 2
    16'b11110100_01100110 : OUT <= 2;  //244 / 102 = 2
    16'b11110100_01100111 : OUT <= 2;  //244 / 103 = 2
    16'b11110100_01101000 : OUT <= 2;  //244 / 104 = 2
    16'b11110100_01101001 : OUT <= 2;  //244 / 105 = 2
    16'b11110100_01101010 : OUT <= 2;  //244 / 106 = 2
    16'b11110100_01101011 : OUT <= 2;  //244 / 107 = 2
    16'b11110100_01101100 : OUT <= 2;  //244 / 108 = 2
    16'b11110100_01101101 : OUT <= 2;  //244 / 109 = 2
    16'b11110100_01101110 : OUT <= 2;  //244 / 110 = 2
    16'b11110100_01101111 : OUT <= 2;  //244 / 111 = 2
    16'b11110100_01110000 : OUT <= 2;  //244 / 112 = 2
    16'b11110100_01110001 : OUT <= 2;  //244 / 113 = 2
    16'b11110100_01110010 : OUT <= 2;  //244 / 114 = 2
    16'b11110100_01110011 : OUT <= 2;  //244 / 115 = 2
    16'b11110100_01110100 : OUT <= 2;  //244 / 116 = 2
    16'b11110100_01110101 : OUT <= 2;  //244 / 117 = 2
    16'b11110100_01110110 : OUT <= 2;  //244 / 118 = 2
    16'b11110100_01110111 : OUT <= 2;  //244 / 119 = 2
    16'b11110100_01111000 : OUT <= 2;  //244 / 120 = 2
    16'b11110100_01111001 : OUT <= 2;  //244 / 121 = 2
    16'b11110100_01111010 : OUT <= 2;  //244 / 122 = 2
    16'b11110100_01111011 : OUT <= 1;  //244 / 123 = 1
    16'b11110100_01111100 : OUT <= 1;  //244 / 124 = 1
    16'b11110100_01111101 : OUT <= 1;  //244 / 125 = 1
    16'b11110100_01111110 : OUT <= 1;  //244 / 126 = 1
    16'b11110100_01111111 : OUT <= 1;  //244 / 127 = 1
    16'b11110100_10000000 : OUT <= 1;  //244 / 128 = 1
    16'b11110100_10000001 : OUT <= 1;  //244 / 129 = 1
    16'b11110100_10000010 : OUT <= 1;  //244 / 130 = 1
    16'b11110100_10000011 : OUT <= 1;  //244 / 131 = 1
    16'b11110100_10000100 : OUT <= 1;  //244 / 132 = 1
    16'b11110100_10000101 : OUT <= 1;  //244 / 133 = 1
    16'b11110100_10000110 : OUT <= 1;  //244 / 134 = 1
    16'b11110100_10000111 : OUT <= 1;  //244 / 135 = 1
    16'b11110100_10001000 : OUT <= 1;  //244 / 136 = 1
    16'b11110100_10001001 : OUT <= 1;  //244 / 137 = 1
    16'b11110100_10001010 : OUT <= 1;  //244 / 138 = 1
    16'b11110100_10001011 : OUT <= 1;  //244 / 139 = 1
    16'b11110100_10001100 : OUT <= 1;  //244 / 140 = 1
    16'b11110100_10001101 : OUT <= 1;  //244 / 141 = 1
    16'b11110100_10001110 : OUT <= 1;  //244 / 142 = 1
    16'b11110100_10001111 : OUT <= 1;  //244 / 143 = 1
    16'b11110100_10010000 : OUT <= 1;  //244 / 144 = 1
    16'b11110100_10010001 : OUT <= 1;  //244 / 145 = 1
    16'b11110100_10010010 : OUT <= 1;  //244 / 146 = 1
    16'b11110100_10010011 : OUT <= 1;  //244 / 147 = 1
    16'b11110100_10010100 : OUT <= 1;  //244 / 148 = 1
    16'b11110100_10010101 : OUT <= 1;  //244 / 149 = 1
    16'b11110100_10010110 : OUT <= 1;  //244 / 150 = 1
    16'b11110100_10010111 : OUT <= 1;  //244 / 151 = 1
    16'b11110100_10011000 : OUT <= 1;  //244 / 152 = 1
    16'b11110100_10011001 : OUT <= 1;  //244 / 153 = 1
    16'b11110100_10011010 : OUT <= 1;  //244 / 154 = 1
    16'b11110100_10011011 : OUT <= 1;  //244 / 155 = 1
    16'b11110100_10011100 : OUT <= 1;  //244 / 156 = 1
    16'b11110100_10011101 : OUT <= 1;  //244 / 157 = 1
    16'b11110100_10011110 : OUT <= 1;  //244 / 158 = 1
    16'b11110100_10011111 : OUT <= 1;  //244 / 159 = 1
    16'b11110100_10100000 : OUT <= 1;  //244 / 160 = 1
    16'b11110100_10100001 : OUT <= 1;  //244 / 161 = 1
    16'b11110100_10100010 : OUT <= 1;  //244 / 162 = 1
    16'b11110100_10100011 : OUT <= 1;  //244 / 163 = 1
    16'b11110100_10100100 : OUT <= 1;  //244 / 164 = 1
    16'b11110100_10100101 : OUT <= 1;  //244 / 165 = 1
    16'b11110100_10100110 : OUT <= 1;  //244 / 166 = 1
    16'b11110100_10100111 : OUT <= 1;  //244 / 167 = 1
    16'b11110100_10101000 : OUT <= 1;  //244 / 168 = 1
    16'b11110100_10101001 : OUT <= 1;  //244 / 169 = 1
    16'b11110100_10101010 : OUT <= 1;  //244 / 170 = 1
    16'b11110100_10101011 : OUT <= 1;  //244 / 171 = 1
    16'b11110100_10101100 : OUT <= 1;  //244 / 172 = 1
    16'b11110100_10101101 : OUT <= 1;  //244 / 173 = 1
    16'b11110100_10101110 : OUT <= 1;  //244 / 174 = 1
    16'b11110100_10101111 : OUT <= 1;  //244 / 175 = 1
    16'b11110100_10110000 : OUT <= 1;  //244 / 176 = 1
    16'b11110100_10110001 : OUT <= 1;  //244 / 177 = 1
    16'b11110100_10110010 : OUT <= 1;  //244 / 178 = 1
    16'b11110100_10110011 : OUT <= 1;  //244 / 179 = 1
    16'b11110100_10110100 : OUT <= 1;  //244 / 180 = 1
    16'b11110100_10110101 : OUT <= 1;  //244 / 181 = 1
    16'b11110100_10110110 : OUT <= 1;  //244 / 182 = 1
    16'b11110100_10110111 : OUT <= 1;  //244 / 183 = 1
    16'b11110100_10111000 : OUT <= 1;  //244 / 184 = 1
    16'b11110100_10111001 : OUT <= 1;  //244 / 185 = 1
    16'b11110100_10111010 : OUT <= 1;  //244 / 186 = 1
    16'b11110100_10111011 : OUT <= 1;  //244 / 187 = 1
    16'b11110100_10111100 : OUT <= 1;  //244 / 188 = 1
    16'b11110100_10111101 : OUT <= 1;  //244 / 189 = 1
    16'b11110100_10111110 : OUT <= 1;  //244 / 190 = 1
    16'b11110100_10111111 : OUT <= 1;  //244 / 191 = 1
    16'b11110100_11000000 : OUT <= 1;  //244 / 192 = 1
    16'b11110100_11000001 : OUT <= 1;  //244 / 193 = 1
    16'b11110100_11000010 : OUT <= 1;  //244 / 194 = 1
    16'b11110100_11000011 : OUT <= 1;  //244 / 195 = 1
    16'b11110100_11000100 : OUT <= 1;  //244 / 196 = 1
    16'b11110100_11000101 : OUT <= 1;  //244 / 197 = 1
    16'b11110100_11000110 : OUT <= 1;  //244 / 198 = 1
    16'b11110100_11000111 : OUT <= 1;  //244 / 199 = 1
    16'b11110100_11001000 : OUT <= 1;  //244 / 200 = 1
    16'b11110100_11001001 : OUT <= 1;  //244 / 201 = 1
    16'b11110100_11001010 : OUT <= 1;  //244 / 202 = 1
    16'b11110100_11001011 : OUT <= 1;  //244 / 203 = 1
    16'b11110100_11001100 : OUT <= 1;  //244 / 204 = 1
    16'b11110100_11001101 : OUT <= 1;  //244 / 205 = 1
    16'b11110100_11001110 : OUT <= 1;  //244 / 206 = 1
    16'b11110100_11001111 : OUT <= 1;  //244 / 207 = 1
    16'b11110100_11010000 : OUT <= 1;  //244 / 208 = 1
    16'b11110100_11010001 : OUT <= 1;  //244 / 209 = 1
    16'b11110100_11010010 : OUT <= 1;  //244 / 210 = 1
    16'b11110100_11010011 : OUT <= 1;  //244 / 211 = 1
    16'b11110100_11010100 : OUT <= 1;  //244 / 212 = 1
    16'b11110100_11010101 : OUT <= 1;  //244 / 213 = 1
    16'b11110100_11010110 : OUT <= 1;  //244 / 214 = 1
    16'b11110100_11010111 : OUT <= 1;  //244 / 215 = 1
    16'b11110100_11011000 : OUT <= 1;  //244 / 216 = 1
    16'b11110100_11011001 : OUT <= 1;  //244 / 217 = 1
    16'b11110100_11011010 : OUT <= 1;  //244 / 218 = 1
    16'b11110100_11011011 : OUT <= 1;  //244 / 219 = 1
    16'b11110100_11011100 : OUT <= 1;  //244 / 220 = 1
    16'b11110100_11011101 : OUT <= 1;  //244 / 221 = 1
    16'b11110100_11011110 : OUT <= 1;  //244 / 222 = 1
    16'b11110100_11011111 : OUT <= 1;  //244 / 223 = 1
    16'b11110100_11100000 : OUT <= 1;  //244 / 224 = 1
    16'b11110100_11100001 : OUT <= 1;  //244 / 225 = 1
    16'b11110100_11100010 : OUT <= 1;  //244 / 226 = 1
    16'b11110100_11100011 : OUT <= 1;  //244 / 227 = 1
    16'b11110100_11100100 : OUT <= 1;  //244 / 228 = 1
    16'b11110100_11100101 : OUT <= 1;  //244 / 229 = 1
    16'b11110100_11100110 : OUT <= 1;  //244 / 230 = 1
    16'b11110100_11100111 : OUT <= 1;  //244 / 231 = 1
    16'b11110100_11101000 : OUT <= 1;  //244 / 232 = 1
    16'b11110100_11101001 : OUT <= 1;  //244 / 233 = 1
    16'b11110100_11101010 : OUT <= 1;  //244 / 234 = 1
    16'b11110100_11101011 : OUT <= 1;  //244 / 235 = 1
    16'b11110100_11101100 : OUT <= 1;  //244 / 236 = 1
    16'b11110100_11101101 : OUT <= 1;  //244 / 237 = 1
    16'b11110100_11101110 : OUT <= 1;  //244 / 238 = 1
    16'b11110100_11101111 : OUT <= 1;  //244 / 239 = 1
    16'b11110100_11110000 : OUT <= 1;  //244 / 240 = 1
    16'b11110100_11110001 : OUT <= 1;  //244 / 241 = 1
    16'b11110100_11110010 : OUT <= 1;  //244 / 242 = 1
    16'b11110100_11110011 : OUT <= 1;  //244 / 243 = 1
    16'b11110100_11110100 : OUT <= 1;  //244 / 244 = 1
    16'b11110100_11110101 : OUT <= 0;  //244 / 245 = 0
    16'b11110100_11110110 : OUT <= 0;  //244 / 246 = 0
    16'b11110100_11110111 : OUT <= 0;  //244 / 247 = 0
    16'b11110100_11111000 : OUT <= 0;  //244 / 248 = 0
    16'b11110100_11111001 : OUT <= 0;  //244 / 249 = 0
    16'b11110100_11111010 : OUT <= 0;  //244 / 250 = 0
    16'b11110100_11111011 : OUT <= 0;  //244 / 251 = 0
    16'b11110100_11111100 : OUT <= 0;  //244 / 252 = 0
    16'b11110100_11111101 : OUT <= 0;  //244 / 253 = 0
    16'b11110100_11111110 : OUT <= 0;  //244 / 254 = 0
    16'b11110100_11111111 : OUT <= 0;  //244 / 255 = 0
    16'b11110101_00000000 : OUT <= 0;  //245 / 0 = 0
    16'b11110101_00000001 : OUT <= 245;  //245 / 1 = 245
    16'b11110101_00000010 : OUT <= 122;  //245 / 2 = 122
    16'b11110101_00000011 : OUT <= 81;  //245 / 3 = 81
    16'b11110101_00000100 : OUT <= 61;  //245 / 4 = 61
    16'b11110101_00000101 : OUT <= 49;  //245 / 5 = 49
    16'b11110101_00000110 : OUT <= 40;  //245 / 6 = 40
    16'b11110101_00000111 : OUT <= 35;  //245 / 7 = 35
    16'b11110101_00001000 : OUT <= 30;  //245 / 8 = 30
    16'b11110101_00001001 : OUT <= 27;  //245 / 9 = 27
    16'b11110101_00001010 : OUT <= 24;  //245 / 10 = 24
    16'b11110101_00001011 : OUT <= 22;  //245 / 11 = 22
    16'b11110101_00001100 : OUT <= 20;  //245 / 12 = 20
    16'b11110101_00001101 : OUT <= 18;  //245 / 13 = 18
    16'b11110101_00001110 : OUT <= 17;  //245 / 14 = 17
    16'b11110101_00001111 : OUT <= 16;  //245 / 15 = 16
    16'b11110101_00010000 : OUT <= 15;  //245 / 16 = 15
    16'b11110101_00010001 : OUT <= 14;  //245 / 17 = 14
    16'b11110101_00010010 : OUT <= 13;  //245 / 18 = 13
    16'b11110101_00010011 : OUT <= 12;  //245 / 19 = 12
    16'b11110101_00010100 : OUT <= 12;  //245 / 20 = 12
    16'b11110101_00010101 : OUT <= 11;  //245 / 21 = 11
    16'b11110101_00010110 : OUT <= 11;  //245 / 22 = 11
    16'b11110101_00010111 : OUT <= 10;  //245 / 23 = 10
    16'b11110101_00011000 : OUT <= 10;  //245 / 24 = 10
    16'b11110101_00011001 : OUT <= 9;  //245 / 25 = 9
    16'b11110101_00011010 : OUT <= 9;  //245 / 26 = 9
    16'b11110101_00011011 : OUT <= 9;  //245 / 27 = 9
    16'b11110101_00011100 : OUT <= 8;  //245 / 28 = 8
    16'b11110101_00011101 : OUT <= 8;  //245 / 29 = 8
    16'b11110101_00011110 : OUT <= 8;  //245 / 30 = 8
    16'b11110101_00011111 : OUT <= 7;  //245 / 31 = 7
    16'b11110101_00100000 : OUT <= 7;  //245 / 32 = 7
    16'b11110101_00100001 : OUT <= 7;  //245 / 33 = 7
    16'b11110101_00100010 : OUT <= 7;  //245 / 34 = 7
    16'b11110101_00100011 : OUT <= 7;  //245 / 35 = 7
    16'b11110101_00100100 : OUT <= 6;  //245 / 36 = 6
    16'b11110101_00100101 : OUT <= 6;  //245 / 37 = 6
    16'b11110101_00100110 : OUT <= 6;  //245 / 38 = 6
    16'b11110101_00100111 : OUT <= 6;  //245 / 39 = 6
    16'b11110101_00101000 : OUT <= 6;  //245 / 40 = 6
    16'b11110101_00101001 : OUT <= 5;  //245 / 41 = 5
    16'b11110101_00101010 : OUT <= 5;  //245 / 42 = 5
    16'b11110101_00101011 : OUT <= 5;  //245 / 43 = 5
    16'b11110101_00101100 : OUT <= 5;  //245 / 44 = 5
    16'b11110101_00101101 : OUT <= 5;  //245 / 45 = 5
    16'b11110101_00101110 : OUT <= 5;  //245 / 46 = 5
    16'b11110101_00101111 : OUT <= 5;  //245 / 47 = 5
    16'b11110101_00110000 : OUT <= 5;  //245 / 48 = 5
    16'b11110101_00110001 : OUT <= 5;  //245 / 49 = 5
    16'b11110101_00110010 : OUT <= 4;  //245 / 50 = 4
    16'b11110101_00110011 : OUT <= 4;  //245 / 51 = 4
    16'b11110101_00110100 : OUT <= 4;  //245 / 52 = 4
    16'b11110101_00110101 : OUT <= 4;  //245 / 53 = 4
    16'b11110101_00110110 : OUT <= 4;  //245 / 54 = 4
    16'b11110101_00110111 : OUT <= 4;  //245 / 55 = 4
    16'b11110101_00111000 : OUT <= 4;  //245 / 56 = 4
    16'b11110101_00111001 : OUT <= 4;  //245 / 57 = 4
    16'b11110101_00111010 : OUT <= 4;  //245 / 58 = 4
    16'b11110101_00111011 : OUT <= 4;  //245 / 59 = 4
    16'b11110101_00111100 : OUT <= 4;  //245 / 60 = 4
    16'b11110101_00111101 : OUT <= 4;  //245 / 61 = 4
    16'b11110101_00111110 : OUT <= 3;  //245 / 62 = 3
    16'b11110101_00111111 : OUT <= 3;  //245 / 63 = 3
    16'b11110101_01000000 : OUT <= 3;  //245 / 64 = 3
    16'b11110101_01000001 : OUT <= 3;  //245 / 65 = 3
    16'b11110101_01000010 : OUT <= 3;  //245 / 66 = 3
    16'b11110101_01000011 : OUT <= 3;  //245 / 67 = 3
    16'b11110101_01000100 : OUT <= 3;  //245 / 68 = 3
    16'b11110101_01000101 : OUT <= 3;  //245 / 69 = 3
    16'b11110101_01000110 : OUT <= 3;  //245 / 70 = 3
    16'b11110101_01000111 : OUT <= 3;  //245 / 71 = 3
    16'b11110101_01001000 : OUT <= 3;  //245 / 72 = 3
    16'b11110101_01001001 : OUT <= 3;  //245 / 73 = 3
    16'b11110101_01001010 : OUT <= 3;  //245 / 74 = 3
    16'b11110101_01001011 : OUT <= 3;  //245 / 75 = 3
    16'b11110101_01001100 : OUT <= 3;  //245 / 76 = 3
    16'b11110101_01001101 : OUT <= 3;  //245 / 77 = 3
    16'b11110101_01001110 : OUT <= 3;  //245 / 78 = 3
    16'b11110101_01001111 : OUT <= 3;  //245 / 79 = 3
    16'b11110101_01010000 : OUT <= 3;  //245 / 80 = 3
    16'b11110101_01010001 : OUT <= 3;  //245 / 81 = 3
    16'b11110101_01010010 : OUT <= 2;  //245 / 82 = 2
    16'b11110101_01010011 : OUT <= 2;  //245 / 83 = 2
    16'b11110101_01010100 : OUT <= 2;  //245 / 84 = 2
    16'b11110101_01010101 : OUT <= 2;  //245 / 85 = 2
    16'b11110101_01010110 : OUT <= 2;  //245 / 86 = 2
    16'b11110101_01010111 : OUT <= 2;  //245 / 87 = 2
    16'b11110101_01011000 : OUT <= 2;  //245 / 88 = 2
    16'b11110101_01011001 : OUT <= 2;  //245 / 89 = 2
    16'b11110101_01011010 : OUT <= 2;  //245 / 90 = 2
    16'b11110101_01011011 : OUT <= 2;  //245 / 91 = 2
    16'b11110101_01011100 : OUT <= 2;  //245 / 92 = 2
    16'b11110101_01011101 : OUT <= 2;  //245 / 93 = 2
    16'b11110101_01011110 : OUT <= 2;  //245 / 94 = 2
    16'b11110101_01011111 : OUT <= 2;  //245 / 95 = 2
    16'b11110101_01100000 : OUT <= 2;  //245 / 96 = 2
    16'b11110101_01100001 : OUT <= 2;  //245 / 97 = 2
    16'b11110101_01100010 : OUT <= 2;  //245 / 98 = 2
    16'b11110101_01100011 : OUT <= 2;  //245 / 99 = 2
    16'b11110101_01100100 : OUT <= 2;  //245 / 100 = 2
    16'b11110101_01100101 : OUT <= 2;  //245 / 101 = 2
    16'b11110101_01100110 : OUT <= 2;  //245 / 102 = 2
    16'b11110101_01100111 : OUT <= 2;  //245 / 103 = 2
    16'b11110101_01101000 : OUT <= 2;  //245 / 104 = 2
    16'b11110101_01101001 : OUT <= 2;  //245 / 105 = 2
    16'b11110101_01101010 : OUT <= 2;  //245 / 106 = 2
    16'b11110101_01101011 : OUT <= 2;  //245 / 107 = 2
    16'b11110101_01101100 : OUT <= 2;  //245 / 108 = 2
    16'b11110101_01101101 : OUT <= 2;  //245 / 109 = 2
    16'b11110101_01101110 : OUT <= 2;  //245 / 110 = 2
    16'b11110101_01101111 : OUT <= 2;  //245 / 111 = 2
    16'b11110101_01110000 : OUT <= 2;  //245 / 112 = 2
    16'b11110101_01110001 : OUT <= 2;  //245 / 113 = 2
    16'b11110101_01110010 : OUT <= 2;  //245 / 114 = 2
    16'b11110101_01110011 : OUT <= 2;  //245 / 115 = 2
    16'b11110101_01110100 : OUT <= 2;  //245 / 116 = 2
    16'b11110101_01110101 : OUT <= 2;  //245 / 117 = 2
    16'b11110101_01110110 : OUT <= 2;  //245 / 118 = 2
    16'b11110101_01110111 : OUT <= 2;  //245 / 119 = 2
    16'b11110101_01111000 : OUT <= 2;  //245 / 120 = 2
    16'b11110101_01111001 : OUT <= 2;  //245 / 121 = 2
    16'b11110101_01111010 : OUT <= 2;  //245 / 122 = 2
    16'b11110101_01111011 : OUT <= 1;  //245 / 123 = 1
    16'b11110101_01111100 : OUT <= 1;  //245 / 124 = 1
    16'b11110101_01111101 : OUT <= 1;  //245 / 125 = 1
    16'b11110101_01111110 : OUT <= 1;  //245 / 126 = 1
    16'b11110101_01111111 : OUT <= 1;  //245 / 127 = 1
    16'b11110101_10000000 : OUT <= 1;  //245 / 128 = 1
    16'b11110101_10000001 : OUT <= 1;  //245 / 129 = 1
    16'b11110101_10000010 : OUT <= 1;  //245 / 130 = 1
    16'b11110101_10000011 : OUT <= 1;  //245 / 131 = 1
    16'b11110101_10000100 : OUT <= 1;  //245 / 132 = 1
    16'b11110101_10000101 : OUT <= 1;  //245 / 133 = 1
    16'b11110101_10000110 : OUT <= 1;  //245 / 134 = 1
    16'b11110101_10000111 : OUT <= 1;  //245 / 135 = 1
    16'b11110101_10001000 : OUT <= 1;  //245 / 136 = 1
    16'b11110101_10001001 : OUT <= 1;  //245 / 137 = 1
    16'b11110101_10001010 : OUT <= 1;  //245 / 138 = 1
    16'b11110101_10001011 : OUT <= 1;  //245 / 139 = 1
    16'b11110101_10001100 : OUT <= 1;  //245 / 140 = 1
    16'b11110101_10001101 : OUT <= 1;  //245 / 141 = 1
    16'b11110101_10001110 : OUT <= 1;  //245 / 142 = 1
    16'b11110101_10001111 : OUT <= 1;  //245 / 143 = 1
    16'b11110101_10010000 : OUT <= 1;  //245 / 144 = 1
    16'b11110101_10010001 : OUT <= 1;  //245 / 145 = 1
    16'b11110101_10010010 : OUT <= 1;  //245 / 146 = 1
    16'b11110101_10010011 : OUT <= 1;  //245 / 147 = 1
    16'b11110101_10010100 : OUT <= 1;  //245 / 148 = 1
    16'b11110101_10010101 : OUT <= 1;  //245 / 149 = 1
    16'b11110101_10010110 : OUT <= 1;  //245 / 150 = 1
    16'b11110101_10010111 : OUT <= 1;  //245 / 151 = 1
    16'b11110101_10011000 : OUT <= 1;  //245 / 152 = 1
    16'b11110101_10011001 : OUT <= 1;  //245 / 153 = 1
    16'b11110101_10011010 : OUT <= 1;  //245 / 154 = 1
    16'b11110101_10011011 : OUT <= 1;  //245 / 155 = 1
    16'b11110101_10011100 : OUT <= 1;  //245 / 156 = 1
    16'b11110101_10011101 : OUT <= 1;  //245 / 157 = 1
    16'b11110101_10011110 : OUT <= 1;  //245 / 158 = 1
    16'b11110101_10011111 : OUT <= 1;  //245 / 159 = 1
    16'b11110101_10100000 : OUT <= 1;  //245 / 160 = 1
    16'b11110101_10100001 : OUT <= 1;  //245 / 161 = 1
    16'b11110101_10100010 : OUT <= 1;  //245 / 162 = 1
    16'b11110101_10100011 : OUT <= 1;  //245 / 163 = 1
    16'b11110101_10100100 : OUT <= 1;  //245 / 164 = 1
    16'b11110101_10100101 : OUT <= 1;  //245 / 165 = 1
    16'b11110101_10100110 : OUT <= 1;  //245 / 166 = 1
    16'b11110101_10100111 : OUT <= 1;  //245 / 167 = 1
    16'b11110101_10101000 : OUT <= 1;  //245 / 168 = 1
    16'b11110101_10101001 : OUT <= 1;  //245 / 169 = 1
    16'b11110101_10101010 : OUT <= 1;  //245 / 170 = 1
    16'b11110101_10101011 : OUT <= 1;  //245 / 171 = 1
    16'b11110101_10101100 : OUT <= 1;  //245 / 172 = 1
    16'b11110101_10101101 : OUT <= 1;  //245 / 173 = 1
    16'b11110101_10101110 : OUT <= 1;  //245 / 174 = 1
    16'b11110101_10101111 : OUT <= 1;  //245 / 175 = 1
    16'b11110101_10110000 : OUT <= 1;  //245 / 176 = 1
    16'b11110101_10110001 : OUT <= 1;  //245 / 177 = 1
    16'b11110101_10110010 : OUT <= 1;  //245 / 178 = 1
    16'b11110101_10110011 : OUT <= 1;  //245 / 179 = 1
    16'b11110101_10110100 : OUT <= 1;  //245 / 180 = 1
    16'b11110101_10110101 : OUT <= 1;  //245 / 181 = 1
    16'b11110101_10110110 : OUT <= 1;  //245 / 182 = 1
    16'b11110101_10110111 : OUT <= 1;  //245 / 183 = 1
    16'b11110101_10111000 : OUT <= 1;  //245 / 184 = 1
    16'b11110101_10111001 : OUT <= 1;  //245 / 185 = 1
    16'b11110101_10111010 : OUT <= 1;  //245 / 186 = 1
    16'b11110101_10111011 : OUT <= 1;  //245 / 187 = 1
    16'b11110101_10111100 : OUT <= 1;  //245 / 188 = 1
    16'b11110101_10111101 : OUT <= 1;  //245 / 189 = 1
    16'b11110101_10111110 : OUT <= 1;  //245 / 190 = 1
    16'b11110101_10111111 : OUT <= 1;  //245 / 191 = 1
    16'b11110101_11000000 : OUT <= 1;  //245 / 192 = 1
    16'b11110101_11000001 : OUT <= 1;  //245 / 193 = 1
    16'b11110101_11000010 : OUT <= 1;  //245 / 194 = 1
    16'b11110101_11000011 : OUT <= 1;  //245 / 195 = 1
    16'b11110101_11000100 : OUT <= 1;  //245 / 196 = 1
    16'b11110101_11000101 : OUT <= 1;  //245 / 197 = 1
    16'b11110101_11000110 : OUT <= 1;  //245 / 198 = 1
    16'b11110101_11000111 : OUT <= 1;  //245 / 199 = 1
    16'b11110101_11001000 : OUT <= 1;  //245 / 200 = 1
    16'b11110101_11001001 : OUT <= 1;  //245 / 201 = 1
    16'b11110101_11001010 : OUT <= 1;  //245 / 202 = 1
    16'b11110101_11001011 : OUT <= 1;  //245 / 203 = 1
    16'b11110101_11001100 : OUT <= 1;  //245 / 204 = 1
    16'b11110101_11001101 : OUT <= 1;  //245 / 205 = 1
    16'b11110101_11001110 : OUT <= 1;  //245 / 206 = 1
    16'b11110101_11001111 : OUT <= 1;  //245 / 207 = 1
    16'b11110101_11010000 : OUT <= 1;  //245 / 208 = 1
    16'b11110101_11010001 : OUT <= 1;  //245 / 209 = 1
    16'b11110101_11010010 : OUT <= 1;  //245 / 210 = 1
    16'b11110101_11010011 : OUT <= 1;  //245 / 211 = 1
    16'b11110101_11010100 : OUT <= 1;  //245 / 212 = 1
    16'b11110101_11010101 : OUT <= 1;  //245 / 213 = 1
    16'b11110101_11010110 : OUT <= 1;  //245 / 214 = 1
    16'b11110101_11010111 : OUT <= 1;  //245 / 215 = 1
    16'b11110101_11011000 : OUT <= 1;  //245 / 216 = 1
    16'b11110101_11011001 : OUT <= 1;  //245 / 217 = 1
    16'b11110101_11011010 : OUT <= 1;  //245 / 218 = 1
    16'b11110101_11011011 : OUT <= 1;  //245 / 219 = 1
    16'b11110101_11011100 : OUT <= 1;  //245 / 220 = 1
    16'b11110101_11011101 : OUT <= 1;  //245 / 221 = 1
    16'b11110101_11011110 : OUT <= 1;  //245 / 222 = 1
    16'b11110101_11011111 : OUT <= 1;  //245 / 223 = 1
    16'b11110101_11100000 : OUT <= 1;  //245 / 224 = 1
    16'b11110101_11100001 : OUT <= 1;  //245 / 225 = 1
    16'b11110101_11100010 : OUT <= 1;  //245 / 226 = 1
    16'b11110101_11100011 : OUT <= 1;  //245 / 227 = 1
    16'b11110101_11100100 : OUT <= 1;  //245 / 228 = 1
    16'b11110101_11100101 : OUT <= 1;  //245 / 229 = 1
    16'b11110101_11100110 : OUT <= 1;  //245 / 230 = 1
    16'b11110101_11100111 : OUT <= 1;  //245 / 231 = 1
    16'b11110101_11101000 : OUT <= 1;  //245 / 232 = 1
    16'b11110101_11101001 : OUT <= 1;  //245 / 233 = 1
    16'b11110101_11101010 : OUT <= 1;  //245 / 234 = 1
    16'b11110101_11101011 : OUT <= 1;  //245 / 235 = 1
    16'b11110101_11101100 : OUT <= 1;  //245 / 236 = 1
    16'b11110101_11101101 : OUT <= 1;  //245 / 237 = 1
    16'b11110101_11101110 : OUT <= 1;  //245 / 238 = 1
    16'b11110101_11101111 : OUT <= 1;  //245 / 239 = 1
    16'b11110101_11110000 : OUT <= 1;  //245 / 240 = 1
    16'b11110101_11110001 : OUT <= 1;  //245 / 241 = 1
    16'b11110101_11110010 : OUT <= 1;  //245 / 242 = 1
    16'b11110101_11110011 : OUT <= 1;  //245 / 243 = 1
    16'b11110101_11110100 : OUT <= 1;  //245 / 244 = 1
    16'b11110101_11110101 : OUT <= 1;  //245 / 245 = 1
    16'b11110101_11110110 : OUT <= 0;  //245 / 246 = 0
    16'b11110101_11110111 : OUT <= 0;  //245 / 247 = 0
    16'b11110101_11111000 : OUT <= 0;  //245 / 248 = 0
    16'b11110101_11111001 : OUT <= 0;  //245 / 249 = 0
    16'b11110101_11111010 : OUT <= 0;  //245 / 250 = 0
    16'b11110101_11111011 : OUT <= 0;  //245 / 251 = 0
    16'b11110101_11111100 : OUT <= 0;  //245 / 252 = 0
    16'b11110101_11111101 : OUT <= 0;  //245 / 253 = 0
    16'b11110101_11111110 : OUT <= 0;  //245 / 254 = 0
    16'b11110101_11111111 : OUT <= 0;  //245 / 255 = 0
    16'b11110110_00000000 : OUT <= 0;  //246 / 0 = 0
    16'b11110110_00000001 : OUT <= 246;  //246 / 1 = 246
    16'b11110110_00000010 : OUT <= 123;  //246 / 2 = 123
    16'b11110110_00000011 : OUT <= 82;  //246 / 3 = 82
    16'b11110110_00000100 : OUT <= 61;  //246 / 4 = 61
    16'b11110110_00000101 : OUT <= 49;  //246 / 5 = 49
    16'b11110110_00000110 : OUT <= 41;  //246 / 6 = 41
    16'b11110110_00000111 : OUT <= 35;  //246 / 7 = 35
    16'b11110110_00001000 : OUT <= 30;  //246 / 8 = 30
    16'b11110110_00001001 : OUT <= 27;  //246 / 9 = 27
    16'b11110110_00001010 : OUT <= 24;  //246 / 10 = 24
    16'b11110110_00001011 : OUT <= 22;  //246 / 11 = 22
    16'b11110110_00001100 : OUT <= 20;  //246 / 12 = 20
    16'b11110110_00001101 : OUT <= 18;  //246 / 13 = 18
    16'b11110110_00001110 : OUT <= 17;  //246 / 14 = 17
    16'b11110110_00001111 : OUT <= 16;  //246 / 15 = 16
    16'b11110110_00010000 : OUT <= 15;  //246 / 16 = 15
    16'b11110110_00010001 : OUT <= 14;  //246 / 17 = 14
    16'b11110110_00010010 : OUT <= 13;  //246 / 18 = 13
    16'b11110110_00010011 : OUT <= 12;  //246 / 19 = 12
    16'b11110110_00010100 : OUT <= 12;  //246 / 20 = 12
    16'b11110110_00010101 : OUT <= 11;  //246 / 21 = 11
    16'b11110110_00010110 : OUT <= 11;  //246 / 22 = 11
    16'b11110110_00010111 : OUT <= 10;  //246 / 23 = 10
    16'b11110110_00011000 : OUT <= 10;  //246 / 24 = 10
    16'b11110110_00011001 : OUT <= 9;  //246 / 25 = 9
    16'b11110110_00011010 : OUT <= 9;  //246 / 26 = 9
    16'b11110110_00011011 : OUT <= 9;  //246 / 27 = 9
    16'b11110110_00011100 : OUT <= 8;  //246 / 28 = 8
    16'b11110110_00011101 : OUT <= 8;  //246 / 29 = 8
    16'b11110110_00011110 : OUT <= 8;  //246 / 30 = 8
    16'b11110110_00011111 : OUT <= 7;  //246 / 31 = 7
    16'b11110110_00100000 : OUT <= 7;  //246 / 32 = 7
    16'b11110110_00100001 : OUT <= 7;  //246 / 33 = 7
    16'b11110110_00100010 : OUT <= 7;  //246 / 34 = 7
    16'b11110110_00100011 : OUT <= 7;  //246 / 35 = 7
    16'b11110110_00100100 : OUT <= 6;  //246 / 36 = 6
    16'b11110110_00100101 : OUT <= 6;  //246 / 37 = 6
    16'b11110110_00100110 : OUT <= 6;  //246 / 38 = 6
    16'b11110110_00100111 : OUT <= 6;  //246 / 39 = 6
    16'b11110110_00101000 : OUT <= 6;  //246 / 40 = 6
    16'b11110110_00101001 : OUT <= 6;  //246 / 41 = 6
    16'b11110110_00101010 : OUT <= 5;  //246 / 42 = 5
    16'b11110110_00101011 : OUT <= 5;  //246 / 43 = 5
    16'b11110110_00101100 : OUT <= 5;  //246 / 44 = 5
    16'b11110110_00101101 : OUT <= 5;  //246 / 45 = 5
    16'b11110110_00101110 : OUT <= 5;  //246 / 46 = 5
    16'b11110110_00101111 : OUT <= 5;  //246 / 47 = 5
    16'b11110110_00110000 : OUT <= 5;  //246 / 48 = 5
    16'b11110110_00110001 : OUT <= 5;  //246 / 49 = 5
    16'b11110110_00110010 : OUT <= 4;  //246 / 50 = 4
    16'b11110110_00110011 : OUT <= 4;  //246 / 51 = 4
    16'b11110110_00110100 : OUT <= 4;  //246 / 52 = 4
    16'b11110110_00110101 : OUT <= 4;  //246 / 53 = 4
    16'b11110110_00110110 : OUT <= 4;  //246 / 54 = 4
    16'b11110110_00110111 : OUT <= 4;  //246 / 55 = 4
    16'b11110110_00111000 : OUT <= 4;  //246 / 56 = 4
    16'b11110110_00111001 : OUT <= 4;  //246 / 57 = 4
    16'b11110110_00111010 : OUT <= 4;  //246 / 58 = 4
    16'b11110110_00111011 : OUT <= 4;  //246 / 59 = 4
    16'b11110110_00111100 : OUT <= 4;  //246 / 60 = 4
    16'b11110110_00111101 : OUT <= 4;  //246 / 61 = 4
    16'b11110110_00111110 : OUT <= 3;  //246 / 62 = 3
    16'b11110110_00111111 : OUT <= 3;  //246 / 63 = 3
    16'b11110110_01000000 : OUT <= 3;  //246 / 64 = 3
    16'b11110110_01000001 : OUT <= 3;  //246 / 65 = 3
    16'b11110110_01000010 : OUT <= 3;  //246 / 66 = 3
    16'b11110110_01000011 : OUT <= 3;  //246 / 67 = 3
    16'b11110110_01000100 : OUT <= 3;  //246 / 68 = 3
    16'b11110110_01000101 : OUT <= 3;  //246 / 69 = 3
    16'b11110110_01000110 : OUT <= 3;  //246 / 70 = 3
    16'b11110110_01000111 : OUT <= 3;  //246 / 71 = 3
    16'b11110110_01001000 : OUT <= 3;  //246 / 72 = 3
    16'b11110110_01001001 : OUT <= 3;  //246 / 73 = 3
    16'b11110110_01001010 : OUT <= 3;  //246 / 74 = 3
    16'b11110110_01001011 : OUT <= 3;  //246 / 75 = 3
    16'b11110110_01001100 : OUT <= 3;  //246 / 76 = 3
    16'b11110110_01001101 : OUT <= 3;  //246 / 77 = 3
    16'b11110110_01001110 : OUT <= 3;  //246 / 78 = 3
    16'b11110110_01001111 : OUT <= 3;  //246 / 79 = 3
    16'b11110110_01010000 : OUT <= 3;  //246 / 80 = 3
    16'b11110110_01010001 : OUT <= 3;  //246 / 81 = 3
    16'b11110110_01010010 : OUT <= 3;  //246 / 82 = 3
    16'b11110110_01010011 : OUT <= 2;  //246 / 83 = 2
    16'b11110110_01010100 : OUT <= 2;  //246 / 84 = 2
    16'b11110110_01010101 : OUT <= 2;  //246 / 85 = 2
    16'b11110110_01010110 : OUT <= 2;  //246 / 86 = 2
    16'b11110110_01010111 : OUT <= 2;  //246 / 87 = 2
    16'b11110110_01011000 : OUT <= 2;  //246 / 88 = 2
    16'b11110110_01011001 : OUT <= 2;  //246 / 89 = 2
    16'b11110110_01011010 : OUT <= 2;  //246 / 90 = 2
    16'b11110110_01011011 : OUT <= 2;  //246 / 91 = 2
    16'b11110110_01011100 : OUT <= 2;  //246 / 92 = 2
    16'b11110110_01011101 : OUT <= 2;  //246 / 93 = 2
    16'b11110110_01011110 : OUT <= 2;  //246 / 94 = 2
    16'b11110110_01011111 : OUT <= 2;  //246 / 95 = 2
    16'b11110110_01100000 : OUT <= 2;  //246 / 96 = 2
    16'b11110110_01100001 : OUT <= 2;  //246 / 97 = 2
    16'b11110110_01100010 : OUT <= 2;  //246 / 98 = 2
    16'b11110110_01100011 : OUT <= 2;  //246 / 99 = 2
    16'b11110110_01100100 : OUT <= 2;  //246 / 100 = 2
    16'b11110110_01100101 : OUT <= 2;  //246 / 101 = 2
    16'b11110110_01100110 : OUT <= 2;  //246 / 102 = 2
    16'b11110110_01100111 : OUT <= 2;  //246 / 103 = 2
    16'b11110110_01101000 : OUT <= 2;  //246 / 104 = 2
    16'b11110110_01101001 : OUT <= 2;  //246 / 105 = 2
    16'b11110110_01101010 : OUT <= 2;  //246 / 106 = 2
    16'b11110110_01101011 : OUT <= 2;  //246 / 107 = 2
    16'b11110110_01101100 : OUT <= 2;  //246 / 108 = 2
    16'b11110110_01101101 : OUT <= 2;  //246 / 109 = 2
    16'b11110110_01101110 : OUT <= 2;  //246 / 110 = 2
    16'b11110110_01101111 : OUT <= 2;  //246 / 111 = 2
    16'b11110110_01110000 : OUT <= 2;  //246 / 112 = 2
    16'b11110110_01110001 : OUT <= 2;  //246 / 113 = 2
    16'b11110110_01110010 : OUT <= 2;  //246 / 114 = 2
    16'b11110110_01110011 : OUT <= 2;  //246 / 115 = 2
    16'b11110110_01110100 : OUT <= 2;  //246 / 116 = 2
    16'b11110110_01110101 : OUT <= 2;  //246 / 117 = 2
    16'b11110110_01110110 : OUT <= 2;  //246 / 118 = 2
    16'b11110110_01110111 : OUT <= 2;  //246 / 119 = 2
    16'b11110110_01111000 : OUT <= 2;  //246 / 120 = 2
    16'b11110110_01111001 : OUT <= 2;  //246 / 121 = 2
    16'b11110110_01111010 : OUT <= 2;  //246 / 122 = 2
    16'b11110110_01111011 : OUT <= 2;  //246 / 123 = 2
    16'b11110110_01111100 : OUT <= 1;  //246 / 124 = 1
    16'b11110110_01111101 : OUT <= 1;  //246 / 125 = 1
    16'b11110110_01111110 : OUT <= 1;  //246 / 126 = 1
    16'b11110110_01111111 : OUT <= 1;  //246 / 127 = 1
    16'b11110110_10000000 : OUT <= 1;  //246 / 128 = 1
    16'b11110110_10000001 : OUT <= 1;  //246 / 129 = 1
    16'b11110110_10000010 : OUT <= 1;  //246 / 130 = 1
    16'b11110110_10000011 : OUT <= 1;  //246 / 131 = 1
    16'b11110110_10000100 : OUT <= 1;  //246 / 132 = 1
    16'b11110110_10000101 : OUT <= 1;  //246 / 133 = 1
    16'b11110110_10000110 : OUT <= 1;  //246 / 134 = 1
    16'b11110110_10000111 : OUT <= 1;  //246 / 135 = 1
    16'b11110110_10001000 : OUT <= 1;  //246 / 136 = 1
    16'b11110110_10001001 : OUT <= 1;  //246 / 137 = 1
    16'b11110110_10001010 : OUT <= 1;  //246 / 138 = 1
    16'b11110110_10001011 : OUT <= 1;  //246 / 139 = 1
    16'b11110110_10001100 : OUT <= 1;  //246 / 140 = 1
    16'b11110110_10001101 : OUT <= 1;  //246 / 141 = 1
    16'b11110110_10001110 : OUT <= 1;  //246 / 142 = 1
    16'b11110110_10001111 : OUT <= 1;  //246 / 143 = 1
    16'b11110110_10010000 : OUT <= 1;  //246 / 144 = 1
    16'b11110110_10010001 : OUT <= 1;  //246 / 145 = 1
    16'b11110110_10010010 : OUT <= 1;  //246 / 146 = 1
    16'b11110110_10010011 : OUT <= 1;  //246 / 147 = 1
    16'b11110110_10010100 : OUT <= 1;  //246 / 148 = 1
    16'b11110110_10010101 : OUT <= 1;  //246 / 149 = 1
    16'b11110110_10010110 : OUT <= 1;  //246 / 150 = 1
    16'b11110110_10010111 : OUT <= 1;  //246 / 151 = 1
    16'b11110110_10011000 : OUT <= 1;  //246 / 152 = 1
    16'b11110110_10011001 : OUT <= 1;  //246 / 153 = 1
    16'b11110110_10011010 : OUT <= 1;  //246 / 154 = 1
    16'b11110110_10011011 : OUT <= 1;  //246 / 155 = 1
    16'b11110110_10011100 : OUT <= 1;  //246 / 156 = 1
    16'b11110110_10011101 : OUT <= 1;  //246 / 157 = 1
    16'b11110110_10011110 : OUT <= 1;  //246 / 158 = 1
    16'b11110110_10011111 : OUT <= 1;  //246 / 159 = 1
    16'b11110110_10100000 : OUT <= 1;  //246 / 160 = 1
    16'b11110110_10100001 : OUT <= 1;  //246 / 161 = 1
    16'b11110110_10100010 : OUT <= 1;  //246 / 162 = 1
    16'b11110110_10100011 : OUT <= 1;  //246 / 163 = 1
    16'b11110110_10100100 : OUT <= 1;  //246 / 164 = 1
    16'b11110110_10100101 : OUT <= 1;  //246 / 165 = 1
    16'b11110110_10100110 : OUT <= 1;  //246 / 166 = 1
    16'b11110110_10100111 : OUT <= 1;  //246 / 167 = 1
    16'b11110110_10101000 : OUT <= 1;  //246 / 168 = 1
    16'b11110110_10101001 : OUT <= 1;  //246 / 169 = 1
    16'b11110110_10101010 : OUT <= 1;  //246 / 170 = 1
    16'b11110110_10101011 : OUT <= 1;  //246 / 171 = 1
    16'b11110110_10101100 : OUT <= 1;  //246 / 172 = 1
    16'b11110110_10101101 : OUT <= 1;  //246 / 173 = 1
    16'b11110110_10101110 : OUT <= 1;  //246 / 174 = 1
    16'b11110110_10101111 : OUT <= 1;  //246 / 175 = 1
    16'b11110110_10110000 : OUT <= 1;  //246 / 176 = 1
    16'b11110110_10110001 : OUT <= 1;  //246 / 177 = 1
    16'b11110110_10110010 : OUT <= 1;  //246 / 178 = 1
    16'b11110110_10110011 : OUT <= 1;  //246 / 179 = 1
    16'b11110110_10110100 : OUT <= 1;  //246 / 180 = 1
    16'b11110110_10110101 : OUT <= 1;  //246 / 181 = 1
    16'b11110110_10110110 : OUT <= 1;  //246 / 182 = 1
    16'b11110110_10110111 : OUT <= 1;  //246 / 183 = 1
    16'b11110110_10111000 : OUT <= 1;  //246 / 184 = 1
    16'b11110110_10111001 : OUT <= 1;  //246 / 185 = 1
    16'b11110110_10111010 : OUT <= 1;  //246 / 186 = 1
    16'b11110110_10111011 : OUT <= 1;  //246 / 187 = 1
    16'b11110110_10111100 : OUT <= 1;  //246 / 188 = 1
    16'b11110110_10111101 : OUT <= 1;  //246 / 189 = 1
    16'b11110110_10111110 : OUT <= 1;  //246 / 190 = 1
    16'b11110110_10111111 : OUT <= 1;  //246 / 191 = 1
    16'b11110110_11000000 : OUT <= 1;  //246 / 192 = 1
    16'b11110110_11000001 : OUT <= 1;  //246 / 193 = 1
    16'b11110110_11000010 : OUT <= 1;  //246 / 194 = 1
    16'b11110110_11000011 : OUT <= 1;  //246 / 195 = 1
    16'b11110110_11000100 : OUT <= 1;  //246 / 196 = 1
    16'b11110110_11000101 : OUT <= 1;  //246 / 197 = 1
    16'b11110110_11000110 : OUT <= 1;  //246 / 198 = 1
    16'b11110110_11000111 : OUT <= 1;  //246 / 199 = 1
    16'b11110110_11001000 : OUT <= 1;  //246 / 200 = 1
    16'b11110110_11001001 : OUT <= 1;  //246 / 201 = 1
    16'b11110110_11001010 : OUT <= 1;  //246 / 202 = 1
    16'b11110110_11001011 : OUT <= 1;  //246 / 203 = 1
    16'b11110110_11001100 : OUT <= 1;  //246 / 204 = 1
    16'b11110110_11001101 : OUT <= 1;  //246 / 205 = 1
    16'b11110110_11001110 : OUT <= 1;  //246 / 206 = 1
    16'b11110110_11001111 : OUT <= 1;  //246 / 207 = 1
    16'b11110110_11010000 : OUT <= 1;  //246 / 208 = 1
    16'b11110110_11010001 : OUT <= 1;  //246 / 209 = 1
    16'b11110110_11010010 : OUT <= 1;  //246 / 210 = 1
    16'b11110110_11010011 : OUT <= 1;  //246 / 211 = 1
    16'b11110110_11010100 : OUT <= 1;  //246 / 212 = 1
    16'b11110110_11010101 : OUT <= 1;  //246 / 213 = 1
    16'b11110110_11010110 : OUT <= 1;  //246 / 214 = 1
    16'b11110110_11010111 : OUT <= 1;  //246 / 215 = 1
    16'b11110110_11011000 : OUT <= 1;  //246 / 216 = 1
    16'b11110110_11011001 : OUT <= 1;  //246 / 217 = 1
    16'b11110110_11011010 : OUT <= 1;  //246 / 218 = 1
    16'b11110110_11011011 : OUT <= 1;  //246 / 219 = 1
    16'b11110110_11011100 : OUT <= 1;  //246 / 220 = 1
    16'b11110110_11011101 : OUT <= 1;  //246 / 221 = 1
    16'b11110110_11011110 : OUT <= 1;  //246 / 222 = 1
    16'b11110110_11011111 : OUT <= 1;  //246 / 223 = 1
    16'b11110110_11100000 : OUT <= 1;  //246 / 224 = 1
    16'b11110110_11100001 : OUT <= 1;  //246 / 225 = 1
    16'b11110110_11100010 : OUT <= 1;  //246 / 226 = 1
    16'b11110110_11100011 : OUT <= 1;  //246 / 227 = 1
    16'b11110110_11100100 : OUT <= 1;  //246 / 228 = 1
    16'b11110110_11100101 : OUT <= 1;  //246 / 229 = 1
    16'b11110110_11100110 : OUT <= 1;  //246 / 230 = 1
    16'b11110110_11100111 : OUT <= 1;  //246 / 231 = 1
    16'b11110110_11101000 : OUT <= 1;  //246 / 232 = 1
    16'b11110110_11101001 : OUT <= 1;  //246 / 233 = 1
    16'b11110110_11101010 : OUT <= 1;  //246 / 234 = 1
    16'b11110110_11101011 : OUT <= 1;  //246 / 235 = 1
    16'b11110110_11101100 : OUT <= 1;  //246 / 236 = 1
    16'b11110110_11101101 : OUT <= 1;  //246 / 237 = 1
    16'b11110110_11101110 : OUT <= 1;  //246 / 238 = 1
    16'b11110110_11101111 : OUT <= 1;  //246 / 239 = 1
    16'b11110110_11110000 : OUT <= 1;  //246 / 240 = 1
    16'b11110110_11110001 : OUT <= 1;  //246 / 241 = 1
    16'b11110110_11110010 : OUT <= 1;  //246 / 242 = 1
    16'b11110110_11110011 : OUT <= 1;  //246 / 243 = 1
    16'b11110110_11110100 : OUT <= 1;  //246 / 244 = 1
    16'b11110110_11110101 : OUT <= 1;  //246 / 245 = 1
    16'b11110110_11110110 : OUT <= 1;  //246 / 246 = 1
    16'b11110110_11110111 : OUT <= 0;  //246 / 247 = 0
    16'b11110110_11111000 : OUT <= 0;  //246 / 248 = 0
    16'b11110110_11111001 : OUT <= 0;  //246 / 249 = 0
    16'b11110110_11111010 : OUT <= 0;  //246 / 250 = 0
    16'b11110110_11111011 : OUT <= 0;  //246 / 251 = 0
    16'b11110110_11111100 : OUT <= 0;  //246 / 252 = 0
    16'b11110110_11111101 : OUT <= 0;  //246 / 253 = 0
    16'b11110110_11111110 : OUT <= 0;  //246 / 254 = 0
    16'b11110110_11111111 : OUT <= 0;  //246 / 255 = 0
    16'b11110111_00000000 : OUT <= 0;  //247 / 0 = 0
    16'b11110111_00000001 : OUT <= 247;  //247 / 1 = 247
    16'b11110111_00000010 : OUT <= 123;  //247 / 2 = 123
    16'b11110111_00000011 : OUT <= 82;  //247 / 3 = 82
    16'b11110111_00000100 : OUT <= 61;  //247 / 4 = 61
    16'b11110111_00000101 : OUT <= 49;  //247 / 5 = 49
    16'b11110111_00000110 : OUT <= 41;  //247 / 6 = 41
    16'b11110111_00000111 : OUT <= 35;  //247 / 7 = 35
    16'b11110111_00001000 : OUT <= 30;  //247 / 8 = 30
    16'b11110111_00001001 : OUT <= 27;  //247 / 9 = 27
    16'b11110111_00001010 : OUT <= 24;  //247 / 10 = 24
    16'b11110111_00001011 : OUT <= 22;  //247 / 11 = 22
    16'b11110111_00001100 : OUT <= 20;  //247 / 12 = 20
    16'b11110111_00001101 : OUT <= 19;  //247 / 13 = 19
    16'b11110111_00001110 : OUT <= 17;  //247 / 14 = 17
    16'b11110111_00001111 : OUT <= 16;  //247 / 15 = 16
    16'b11110111_00010000 : OUT <= 15;  //247 / 16 = 15
    16'b11110111_00010001 : OUT <= 14;  //247 / 17 = 14
    16'b11110111_00010010 : OUT <= 13;  //247 / 18 = 13
    16'b11110111_00010011 : OUT <= 13;  //247 / 19 = 13
    16'b11110111_00010100 : OUT <= 12;  //247 / 20 = 12
    16'b11110111_00010101 : OUT <= 11;  //247 / 21 = 11
    16'b11110111_00010110 : OUT <= 11;  //247 / 22 = 11
    16'b11110111_00010111 : OUT <= 10;  //247 / 23 = 10
    16'b11110111_00011000 : OUT <= 10;  //247 / 24 = 10
    16'b11110111_00011001 : OUT <= 9;  //247 / 25 = 9
    16'b11110111_00011010 : OUT <= 9;  //247 / 26 = 9
    16'b11110111_00011011 : OUT <= 9;  //247 / 27 = 9
    16'b11110111_00011100 : OUT <= 8;  //247 / 28 = 8
    16'b11110111_00011101 : OUT <= 8;  //247 / 29 = 8
    16'b11110111_00011110 : OUT <= 8;  //247 / 30 = 8
    16'b11110111_00011111 : OUT <= 7;  //247 / 31 = 7
    16'b11110111_00100000 : OUT <= 7;  //247 / 32 = 7
    16'b11110111_00100001 : OUT <= 7;  //247 / 33 = 7
    16'b11110111_00100010 : OUT <= 7;  //247 / 34 = 7
    16'b11110111_00100011 : OUT <= 7;  //247 / 35 = 7
    16'b11110111_00100100 : OUT <= 6;  //247 / 36 = 6
    16'b11110111_00100101 : OUT <= 6;  //247 / 37 = 6
    16'b11110111_00100110 : OUT <= 6;  //247 / 38 = 6
    16'b11110111_00100111 : OUT <= 6;  //247 / 39 = 6
    16'b11110111_00101000 : OUT <= 6;  //247 / 40 = 6
    16'b11110111_00101001 : OUT <= 6;  //247 / 41 = 6
    16'b11110111_00101010 : OUT <= 5;  //247 / 42 = 5
    16'b11110111_00101011 : OUT <= 5;  //247 / 43 = 5
    16'b11110111_00101100 : OUT <= 5;  //247 / 44 = 5
    16'b11110111_00101101 : OUT <= 5;  //247 / 45 = 5
    16'b11110111_00101110 : OUT <= 5;  //247 / 46 = 5
    16'b11110111_00101111 : OUT <= 5;  //247 / 47 = 5
    16'b11110111_00110000 : OUT <= 5;  //247 / 48 = 5
    16'b11110111_00110001 : OUT <= 5;  //247 / 49 = 5
    16'b11110111_00110010 : OUT <= 4;  //247 / 50 = 4
    16'b11110111_00110011 : OUT <= 4;  //247 / 51 = 4
    16'b11110111_00110100 : OUT <= 4;  //247 / 52 = 4
    16'b11110111_00110101 : OUT <= 4;  //247 / 53 = 4
    16'b11110111_00110110 : OUT <= 4;  //247 / 54 = 4
    16'b11110111_00110111 : OUT <= 4;  //247 / 55 = 4
    16'b11110111_00111000 : OUT <= 4;  //247 / 56 = 4
    16'b11110111_00111001 : OUT <= 4;  //247 / 57 = 4
    16'b11110111_00111010 : OUT <= 4;  //247 / 58 = 4
    16'b11110111_00111011 : OUT <= 4;  //247 / 59 = 4
    16'b11110111_00111100 : OUT <= 4;  //247 / 60 = 4
    16'b11110111_00111101 : OUT <= 4;  //247 / 61 = 4
    16'b11110111_00111110 : OUT <= 3;  //247 / 62 = 3
    16'b11110111_00111111 : OUT <= 3;  //247 / 63 = 3
    16'b11110111_01000000 : OUT <= 3;  //247 / 64 = 3
    16'b11110111_01000001 : OUT <= 3;  //247 / 65 = 3
    16'b11110111_01000010 : OUT <= 3;  //247 / 66 = 3
    16'b11110111_01000011 : OUT <= 3;  //247 / 67 = 3
    16'b11110111_01000100 : OUT <= 3;  //247 / 68 = 3
    16'b11110111_01000101 : OUT <= 3;  //247 / 69 = 3
    16'b11110111_01000110 : OUT <= 3;  //247 / 70 = 3
    16'b11110111_01000111 : OUT <= 3;  //247 / 71 = 3
    16'b11110111_01001000 : OUT <= 3;  //247 / 72 = 3
    16'b11110111_01001001 : OUT <= 3;  //247 / 73 = 3
    16'b11110111_01001010 : OUT <= 3;  //247 / 74 = 3
    16'b11110111_01001011 : OUT <= 3;  //247 / 75 = 3
    16'b11110111_01001100 : OUT <= 3;  //247 / 76 = 3
    16'b11110111_01001101 : OUT <= 3;  //247 / 77 = 3
    16'b11110111_01001110 : OUT <= 3;  //247 / 78 = 3
    16'b11110111_01001111 : OUT <= 3;  //247 / 79 = 3
    16'b11110111_01010000 : OUT <= 3;  //247 / 80 = 3
    16'b11110111_01010001 : OUT <= 3;  //247 / 81 = 3
    16'b11110111_01010010 : OUT <= 3;  //247 / 82 = 3
    16'b11110111_01010011 : OUT <= 2;  //247 / 83 = 2
    16'b11110111_01010100 : OUT <= 2;  //247 / 84 = 2
    16'b11110111_01010101 : OUT <= 2;  //247 / 85 = 2
    16'b11110111_01010110 : OUT <= 2;  //247 / 86 = 2
    16'b11110111_01010111 : OUT <= 2;  //247 / 87 = 2
    16'b11110111_01011000 : OUT <= 2;  //247 / 88 = 2
    16'b11110111_01011001 : OUT <= 2;  //247 / 89 = 2
    16'b11110111_01011010 : OUT <= 2;  //247 / 90 = 2
    16'b11110111_01011011 : OUT <= 2;  //247 / 91 = 2
    16'b11110111_01011100 : OUT <= 2;  //247 / 92 = 2
    16'b11110111_01011101 : OUT <= 2;  //247 / 93 = 2
    16'b11110111_01011110 : OUT <= 2;  //247 / 94 = 2
    16'b11110111_01011111 : OUT <= 2;  //247 / 95 = 2
    16'b11110111_01100000 : OUT <= 2;  //247 / 96 = 2
    16'b11110111_01100001 : OUT <= 2;  //247 / 97 = 2
    16'b11110111_01100010 : OUT <= 2;  //247 / 98 = 2
    16'b11110111_01100011 : OUT <= 2;  //247 / 99 = 2
    16'b11110111_01100100 : OUT <= 2;  //247 / 100 = 2
    16'b11110111_01100101 : OUT <= 2;  //247 / 101 = 2
    16'b11110111_01100110 : OUT <= 2;  //247 / 102 = 2
    16'b11110111_01100111 : OUT <= 2;  //247 / 103 = 2
    16'b11110111_01101000 : OUT <= 2;  //247 / 104 = 2
    16'b11110111_01101001 : OUT <= 2;  //247 / 105 = 2
    16'b11110111_01101010 : OUT <= 2;  //247 / 106 = 2
    16'b11110111_01101011 : OUT <= 2;  //247 / 107 = 2
    16'b11110111_01101100 : OUT <= 2;  //247 / 108 = 2
    16'b11110111_01101101 : OUT <= 2;  //247 / 109 = 2
    16'b11110111_01101110 : OUT <= 2;  //247 / 110 = 2
    16'b11110111_01101111 : OUT <= 2;  //247 / 111 = 2
    16'b11110111_01110000 : OUT <= 2;  //247 / 112 = 2
    16'b11110111_01110001 : OUT <= 2;  //247 / 113 = 2
    16'b11110111_01110010 : OUT <= 2;  //247 / 114 = 2
    16'b11110111_01110011 : OUT <= 2;  //247 / 115 = 2
    16'b11110111_01110100 : OUT <= 2;  //247 / 116 = 2
    16'b11110111_01110101 : OUT <= 2;  //247 / 117 = 2
    16'b11110111_01110110 : OUT <= 2;  //247 / 118 = 2
    16'b11110111_01110111 : OUT <= 2;  //247 / 119 = 2
    16'b11110111_01111000 : OUT <= 2;  //247 / 120 = 2
    16'b11110111_01111001 : OUT <= 2;  //247 / 121 = 2
    16'b11110111_01111010 : OUT <= 2;  //247 / 122 = 2
    16'b11110111_01111011 : OUT <= 2;  //247 / 123 = 2
    16'b11110111_01111100 : OUT <= 1;  //247 / 124 = 1
    16'b11110111_01111101 : OUT <= 1;  //247 / 125 = 1
    16'b11110111_01111110 : OUT <= 1;  //247 / 126 = 1
    16'b11110111_01111111 : OUT <= 1;  //247 / 127 = 1
    16'b11110111_10000000 : OUT <= 1;  //247 / 128 = 1
    16'b11110111_10000001 : OUT <= 1;  //247 / 129 = 1
    16'b11110111_10000010 : OUT <= 1;  //247 / 130 = 1
    16'b11110111_10000011 : OUT <= 1;  //247 / 131 = 1
    16'b11110111_10000100 : OUT <= 1;  //247 / 132 = 1
    16'b11110111_10000101 : OUT <= 1;  //247 / 133 = 1
    16'b11110111_10000110 : OUT <= 1;  //247 / 134 = 1
    16'b11110111_10000111 : OUT <= 1;  //247 / 135 = 1
    16'b11110111_10001000 : OUT <= 1;  //247 / 136 = 1
    16'b11110111_10001001 : OUT <= 1;  //247 / 137 = 1
    16'b11110111_10001010 : OUT <= 1;  //247 / 138 = 1
    16'b11110111_10001011 : OUT <= 1;  //247 / 139 = 1
    16'b11110111_10001100 : OUT <= 1;  //247 / 140 = 1
    16'b11110111_10001101 : OUT <= 1;  //247 / 141 = 1
    16'b11110111_10001110 : OUT <= 1;  //247 / 142 = 1
    16'b11110111_10001111 : OUT <= 1;  //247 / 143 = 1
    16'b11110111_10010000 : OUT <= 1;  //247 / 144 = 1
    16'b11110111_10010001 : OUT <= 1;  //247 / 145 = 1
    16'b11110111_10010010 : OUT <= 1;  //247 / 146 = 1
    16'b11110111_10010011 : OUT <= 1;  //247 / 147 = 1
    16'b11110111_10010100 : OUT <= 1;  //247 / 148 = 1
    16'b11110111_10010101 : OUT <= 1;  //247 / 149 = 1
    16'b11110111_10010110 : OUT <= 1;  //247 / 150 = 1
    16'b11110111_10010111 : OUT <= 1;  //247 / 151 = 1
    16'b11110111_10011000 : OUT <= 1;  //247 / 152 = 1
    16'b11110111_10011001 : OUT <= 1;  //247 / 153 = 1
    16'b11110111_10011010 : OUT <= 1;  //247 / 154 = 1
    16'b11110111_10011011 : OUT <= 1;  //247 / 155 = 1
    16'b11110111_10011100 : OUT <= 1;  //247 / 156 = 1
    16'b11110111_10011101 : OUT <= 1;  //247 / 157 = 1
    16'b11110111_10011110 : OUT <= 1;  //247 / 158 = 1
    16'b11110111_10011111 : OUT <= 1;  //247 / 159 = 1
    16'b11110111_10100000 : OUT <= 1;  //247 / 160 = 1
    16'b11110111_10100001 : OUT <= 1;  //247 / 161 = 1
    16'b11110111_10100010 : OUT <= 1;  //247 / 162 = 1
    16'b11110111_10100011 : OUT <= 1;  //247 / 163 = 1
    16'b11110111_10100100 : OUT <= 1;  //247 / 164 = 1
    16'b11110111_10100101 : OUT <= 1;  //247 / 165 = 1
    16'b11110111_10100110 : OUT <= 1;  //247 / 166 = 1
    16'b11110111_10100111 : OUT <= 1;  //247 / 167 = 1
    16'b11110111_10101000 : OUT <= 1;  //247 / 168 = 1
    16'b11110111_10101001 : OUT <= 1;  //247 / 169 = 1
    16'b11110111_10101010 : OUT <= 1;  //247 / 170 = 1
    16'b11110111_10101011 : OUT <= 1;  //247 / 171 = 1
    16'b11110111_10101100 : OUT <= 1;  //247 / 172 = 1
    16'b11110111_10101101 : OUT <= 1;  //247 / 173 = 1
    16'b11110111_10101110 : OUT <= 1;  //247 / 174 = 1
    16'b11110111_10101111 : OUT <= 1;  //247 / 175 = 1
    16'b11110111_10110000 : OUT <= 1;  //247 / 176 = 1
    16'b11110111_10110001 : OUT <= 1;  //247 / 177 = 1
    16'b11110111_10110010 : OUT <= 1;  //247 / 178 = 1
    16'b11110111_10110011 : OUT <= 1;  //247 / 179 = 1
    16'b11110111_10110100 : OUT <= 1;  //247 / 180 = 1
    16'b11110111_10110101 : OUT <= 1;  //247 / 181 = 1
    16'b11110111_10110110 : OUT <= 1;  //247 / 182 = 1
    16'b11110111_10110111 : OUT <= 1;  //247 / 183 = 1
    16'b11110111_10111000 : OUT <= 1;  //247 / 184 = 1
    16'b11110111_10111001 : OUT <= 1;  //247 / 185 = 1
    16'b11110111_10111010 : OUT <= 1;  //247 / 186 = 1
    16'b11110111_10111011 : OUT <= 1;  //247 / 187 = 1
    16'b11110111_10111100 : OUT <= 1;  //247 / 188 = 1
    16'b11110111_10111101 : OUT <= 1;  //247 / 189 = 1
    16'b11110111_10111110 : OUT <= 1;  //247 / 190 = 1
    16'b11110111_10111111 : OUT <= 1;  //247 / 191 = 1
    16'b11110111_11000000 : OUT <= 1;  //247 / 192 = 1
    16'b11110111_11000001 : OUT <= 1;  //247 / 193 = 1
    16'b11110111_11000010 : OUT <= 1;  //247 / 194 = 1
    16'b11110111_11000011 : OUT <= 1;  //247 / 195 = 1
    16'b11110111_11000100 : OUT <= 1;  //247 / 196 = 1
    16'b11110111_11000101 : OUT <= 1;  //247 / 197 = 1
    16'b11110111_11000110 : OUT <= 1;  //247 / 198 = 1
    16'b11110111_11000111 : OUT <= 1;  //247 / 199 = 1
    16'b11110111_11001000 : OUT <= 1;  //247 / 200 = 1
    16'b11110111_11001001 : OUT <= 1;  //247 / 201 = 1
    16'b11110111_11001010 : OUT <= 1;  //247 / 202 = 1
    16'b11110111_11001011 : OUT <= 1;  //247 / 203 = 1
    16'b11110111_11001100 : OUT <= 1;  //247 / 204 = 1
    16'b11110111_11001101 : OUT <= 1;  //247 / 205 = 1
    16'b11110111_11001110 : OUT <= 1;  //247 / 206 = 1
    16'b11110111_11001111 : OUT <= 1;  //247 / 207 = 1
    16'b11110111_11010000 : OUT <= 1;  //247 / 208 = 1
    16'b11110111_11010001 : OUT <= 1;  //247 / 209 = 1
    16'b11110111_11010010 : OUT <= 1;  //247 / 210 = 1
    16'b11110111_11010011 : OUT <= 1;  //247 / 211 = 1
    16'b11110111_11010100 : OUT <= 1;  //247 / 212 = 1
    16'b11110111_11010101 : OUT <= 1;  //247 / 213 = 1
    16'b11110111_11010110 : OUT <= 1;  //247 / 214 = 1
    16'b11110111_11010111 : OUT <= 1;  //247 / 215 = 1
    16'b11110111_11011000 : OUT <= 1;  //247 / 216 = 1
    16'b11110111_11011001 : OUT <= 1;  //247 / 217 = 1
    16'b11110111_11011010 : OUT <= 1;  //247 / 218 = 1
    16'b11110111_11011011 : OUT <= 1;  //247 / 219 = 1
    16'b11110111_11011100 : OUT <= 1;  //247 / 220 = 1
    16'b11110111_11011101 : OUT <= 1;  //247 / 221 = 1
    16'b11110111_11011110 : OUT <= 1;  //247 / 222 = 1
    16'b11110111_11011111 : OUT <= 1;  //247 / 223 = 1
    16'b11110111_11100000 : OUT <= 1;  //247 / 224 = 1
    16'b11110111_11100001 : OUT <= 1;  //247 / 225 = 1
    16'b11110111_11100010 : OUT <= 1;  //247 / 226 = 1
    16'b11110111_11100011 : OUT <= 1;  //247 / 227 = 1
    16'b11110111_11100100 : OUT <= 1;  //247 / 228 = 1
    16'b11110111_11100101 : OUT <= 1;  //247 / 229 = 1
    16'b11110111_11100110 : OUT <= 1;  //247 / 230 = 1
    16'b11110111_11100111 : OUT <= 1;  //247 / 231 = 1
    16'b11110111_11101000 : OUT <= 1;  //247 / 232 = 1
    16'b11110111_11101001 : OUT <= 1;  //247 / 233 = 1
    16'b11110111_11101010 : OUT <= 1;  //247 / 234 = 1
    16'b11110111_11101011 : OUT <= 1;  //247 / 235 = 1
    16'b11110111_11101100 : OUT <= 1;  //247 / 236 = 1
    16'b11110111_11101101 : OUT <= 1;  //247 / 237 = 1
    16'b11110111_11101110 : OUT <= 1;  //247 / 238 = 1
    16'b11110111_11101111 : OUT <= 1;  //247 / 239 = 1
    16'b11110111_11110000 : OUT <= 1;  //247 / 240 = 1
    16'b11110111_11110001 : OUT <= 1;  //247 / 241 = 1
    16'b11110111_11110010 : OUT <= 1;  //247 / 242 = 1
    16'b11110111_11110011 : OUT <= 1;  //247 / 243 = 1
    16'b11110111_11110100 : OUT <= 1;  //247 / 244 = 1
    16'b11110111_11110101 : OUT <= 1;  //247 / 245 = 1
    16'b11110111_11110110 : OUT <= 1;  //247 / 246 = 1
    16'b11110111_11110111 : OUT <= 1;  //247 / 247 = 1
    16'b11110111_11111000 : OUT <= 0;  //247 / 248 = 0
    16'b11110111_11111001 : OUT <= 0;  //247 / 249 = 0
    16'b11110111_11111010 : OUT <= 0;  //247 / 250 = 0
    16'b11110111_11111011 : OUT <= 0;  //247 / 251 = 0
    16'b11110111_11111100 : OUT <= 0;  //247 / 252 = 0
    16'b11110111_11111101 : OUT <= 0;  //247 / 253 = 0
    16'b11110111_11111110 : OUT <= 0;  //247 / 254 = 0
    16'b11110111_11111111 : OUT <= 0;  //247 / 255 = 0
    16'b11111000_00000000 : OUT <= 0;  //248 / 0 = 0
    16'b11111000_00000001 : OUT <= 248;  //248 / 1 = 248
    16'b11111000_00000010 : OUT <= 124;  //248 / 2 = 124
    16'b11111000_00000011 : OUT <= 82;  //248 / 3 = 82
    16'b11111000_00000100 : OUT <= 62;  //248 / 4 = 62
    16'b11111000_00000101 : OUT <= 49;  //248 / 5 = 49
    16'b11111000_00000110 : OUT <= 41;  //248 / 6 = 41
    16'b11111000_00000111 : OUT <= 35;  //248 / 7 = 35
    16'b11111000_00001000 : OUT <= 31;  //248 / 8 = 31
    16'b11111000_00001001 : OUT <= 27;  //248 / 9 = 27
    16'b11111000_00001010 : OUT <= 24;  //248 / 10 = 24
    16'b11111000_00001011 : OUT <= 22;  //248 / 11 = 22
    16'b11111000_00001100 : OUT <= 20;  //248 / 12 = 20
    16'b11111000_00001101 : OUT <= 19;  //248 / 13 = 19
    16'b11111000_00001110 : OUT <= 17;  //248 / 14 = 17
    16'b11111000_00001111 : OUT <= 16;  //248 / 15 = 16
    16'b11111000_00010000 : OUT <= 15;  //248 / 16 = 15
    16'b11111000_00010001 : OUT <= 14;  //248 / 17 = 14
    16'b11111000_00010010 : OUT <= 13;  //248 / 18 = 13
    16'b11111000_00010011 : OUT <= 13;  //248 / 19 = 13
    16'b11111000_00010100 : OUT <= 12;  //248 / 20 = 12
    16'b11111000_00010101 : OUT <= 11;  //248 / 21 = 11
    16'b11111000_00010110 : OUT <= 11;  //248 / 22 = 11
    16'b11111000_00010111 : OUT <= 10;  //248 / 23 = 10
    16'b11111000_00011000 : OUT <= 10;  //248 / 24 = 10
    16'b11111000_00011001 : OUT <= 9;  //248 / 25 = 9
    16'b11111000_00011010 : OUT <= 9;  //248 / 26 = 9
    16'b11111000_00011011 : OUT <= 9;  //248 / 27 = 9
    16'b11111000_00011100 : OUT <= 8;  //248 / 28 = 8
    16'b11111000_00011101 : OUT <= 8;  //248 / 29 = 8
    16'b11111000_00011110 : OUT <= 8;  //248 / 30 = 8
    16'b11111000_00011111 : OUT <= 8;  //248 / 31 = 8
    16'b11111000_00100000 : OUT <= 7;  //248 / 32 = 7
    16'b11111000_00100001 : OUT <= 7;  //248 / 33 = 7
    16'b11111000_00100010 : OUT <= 7;  //248 / 34 = 7
    16'b11111000_00100011 : OUT <= 7;  //248 / 35 = 7
    16'b11111000_00100100 : OUT <= 6;  //248 / 36 = 6
    16'b11111000_00100101 : OUT <= 6;  //248 / 37 = 6
    16'b11111000_00100110 : OUT <= 6;  //248 / 38 = 6
    16'b11111000_00100111 : OUT <= 6;  //248 / 39 = 6
    16'b11111000_00101000 : OUT <= 6;  //248 / 40 = 6
    16'b11111000_00101001 : OUT <= 6;  //248 / 41 = 6
    16'b11111000_00101010 : OUT <= 5;  //248 / 42 = 5
    16'b11111000_00101011 : OUT <= 5;  //248 / 43 = 5
    16'b11111000_00101100 : OUT <= 5;  //248 / 44 = 5
    16'b11111000_00101101 : OUT <= 5;  //248 / 45 = 5
    16'b11111000_00101110 : OUT <= 5;  //248 / 46 = 5
    16'b11111000_00101111 : OUT <= 5;  //248 / 47 = 5
    16'b11111000_00110000 : OUT <= 5;  //248 / 48 = 5
    16'b11111000_00110001 : OUT <= 5;  //248 / 49 = 5
    16'b11111000_00110010 : OUT <= 4;  //248 / 50 = 4
    16'b11111000_00110011 : OUT <= 4;  //248 / 51 = 4
    16'b11111000_00110100 : OUT <= 4;  //248 / 52 = 4
    16'b11111000_00110101 : OUT <= 4;  //248 / 53 = 4
    16'b11111000_00110110 : OUT <= 4;  //248 / 54 = 4
    16'b11111000_00110111 : OUT <= 4;  //248 / 55 = 4
    16'b11111000_00111000 : OUT <= 4;  //248 / 56 = 4
    16'b11111000_00111001 : OUT <= 4;  //248 / 57 = 4
    16'b11111000_00111010 : OUT <= 4;  //248 / 58 = 4
    16'b11111000_00111011 : OUT <= 4;  //248 / 59 = 4
    16'b11111000_00111100 : OUT <= 4;  //248 / 60 = 4
    16'b11111000_00111101 : OUT <= 4;  //248 / 61 = 4
    16'b11111000_00111110 : OUT <= 4;  //248 / 62 = 4
    16'b11111000_00111111 : OUT <= 3;  //248 / 63 = 3
    16'b11111000_01000000 : OUT <= 3;  //248 / 64 = 3
    16'b11111000_01000001 : OUT <= 3;  //248 / 65 = 3
    16'b11111000_01000010 : OUT <= 3;  //248 / 66 = 3
    16'b11111000_01000011 : OUT <= 3;  //248 / 67 = 3
    16'b11111000_01000100 : OUT <= 3;  //248 / 68 = 3
    16'b11111000_01000101 : OUT <= 3;  //248 / 69 = 3
    16'b11111000_01000110 : OUT <= 3;  //248 / 70 = 3
    16'b11111000_01000111 : OUT <= 3;  //248 / 71 = 3
    16'b11111000_01001000 : OUT <= 3;  //248 / 72 = 3
    16'b11111000_01001001 : OUT <= 3;  //248 / 73 = 3
    16'b11111000_01001010 : OUT <= 3;  //248 / 74 = 3
    16'b11111000_01001011 : OUT <= 3;  //248 / 75 = 3
    16'b11111000_01001100 : OUT <= 3;  //248 / 76 = 3
    16'b11111000_01001101 : OUT <= 3;  //248 / 77 = 3
    16'b11111000_01001110 : OUT <= 3;  //248 / 78 = 3
    16'b11111000_01001111 : OUT <= 3;  //248 / 79 = 3
    16'b11111000_01010000 : OUT <= 3;  //248 / 80 = 3
    16'b11111000_01010001 : OUT <= 3;  //248 / 81 = 3
    16'b11111000_01010010 : OUT <= 3;  //248 / 82 = 3
    16'b11111000_01010011 : OUT <= 2;  //248 / 83 = 2
    16'b11111000_01010100 : OUT <= 2;  //248 / 84 = 2
    16'b11111000_01010101 : OUT <= 2;  //248 / 85 = 2
    16'b11111000_01010110 : OUT <= 2;  //248 / 86 = 2
    16'b11111000_01010111 : OUT <= 2;  //248 / 87 = 2
    16'b11111000_01011000 : OUT <= 2;  //248 / 88 = 2
    16'b11111000_01011001 : OUT <= 2;  //248 / 89 = 2
    16'b11111000_01011010 : OUT <= 2;  //248 / 90 = 2
    16'b11111000_01011011 : OUT <= 2;  //248 / 91 = 2
    16'b11111000_01011100 : OUT <= 2;  //248 / 92 = 2
    16'b11111000_01011101 : OUT <= 2;  //248 / 93 = 2
    16'b11111000_01011110 : OUT <= 2;  //248 / 94 = 2
    16'b11111000_01011111 : OUT <= 2;  //248 / 95 = 2
    16'b11111000_01100000 : OUT <= 2;  //248 / 96 = 2
    16'b11111000_01100001 : OUT <= 2;  //248 / 97 = 2
    16'b11111000_01100010 : OUT <= 2;  //248 / 98 = 2
    16'b11111000_01100011 : OUT <= 2;  //248 / 99 = 2
    16'b11111000_01100100 : OUT <= 2;  //248 / 100 = 2
    16'b11111000_01100101 : OUT <= 2;  //248 / 101 = 2
    16'b11111000_01100110 : OUT <= 2;  //248 / 102 = 2
    16'b11111000_01100111 : OUT <= 2;  //248 / 103 = 2
    16'b11111000_01101000 : OUT <= 2;  //248 / 104 = 2
    16'b11111000_01101001 : OUT <= 2;  //248 / 105 = 2
    16'b11111000_01101010 : OUT <= 2;  //248 / 106 = 2
    16'b11111000_01101011 : OUT <= 2;  //248 / 107 = 2
    16'b11111000_01101100 : OUT <= 2;  //248 / 108 = 2
    16'b11111000_01101101 : OUT <= 2;  //248 / 109 = 2
    16'b11111000_01101110 : OUT <= 2;  //248 / 110 = 2
    16'b11111000_01101111 : OUT <= 2;  //248 / 111 = 2
    16'b11111000_01110000 : OUT <= 2;  //248 / 112 = 2
    16'b11111000_01110001 : OUT <= 2;  //248 / 113 = 2
    16'b11111000_01110010 : OUT <= 2;  //248 / 114 = 2
    16'b11111000_01110011 : OUT <= 2;  //248 / 115 = 2
    16'b11111000_01110100 : OUT <= 2;  //248 / 116 = 2
    16'b11111000_01110101 : OUT <= 2;  //248 / 117 = 2
    16'b11111000_01110110 : OUT <= 2;  //248 / 118 = 2
    16'b11111000_01110111 : OUT <= 2;  //248 / 119 = 2
    16'b11111000_01111000 : OUT <= 2;  //248 / 120 = 2
    16'b11111000_01111001 : OUT <= 2;  //248 / 121 = 2
    16'b11111000_01111010 : OUT <= 2;  //248 / 122 = 2
    16'b11111000_01111011 : OUT <= 2;  //248 / 123 = 2
    16'b11111000_01111100 : OUT <= 2;  //248 / 124 = 2
    16'b11111000_01111101 : OUT <= 1;  //248 / 125 = 1
    16'b11111000_01111110 : OUT <= 1;  //248 / 126 = 1
    16'b11111000_01111111 : OUT <= 1;  //248 / 127 = 1
    16'b11111000_10000000 : OUT <= 1;  //248 / 128 = 1
    16'b11111000_10000001 : OUT <= 1;  //248 / 129 = 1
    16'b11111000_10000010 : OUT <= 1;  //248 / 130 = 1
    16'b11111000_10000011 : OUT <= 1;  //248 / 131 = 1
    16'b11111000_10000100 : OUT <= 1;  //248 / 132 = 1
    16'b11111000_10000101 : OUT <= 1;  //248 / 133 = 1
    16'b11111000_10000110 : OUT <= 1;  //248 / 134 = 1
    16'b11111000_10000111 : OUT <= 1;  //248 / 135 = 1
    16'b11111000_10001000 : OUT <= 1;  //248 / 136 = 1
    16'b11111000_10001001 : OUT <= 1;  //248 / 137 = 1
    16'b11111000_10001010 : OUT <= 1;  //248 / 138 = 1
    16'b11111000_10001011 : OUT <= 1;  //248 / 139 = 1
    16'b11111000_10001100 : OUT <= 1;  //248 / 140 = 1
    16'b11111000_10001101 : OUT <= 1;  //248 / 141 = 1
    16'b11111000_10001110 : OUT <= 1;  //248 / 142 = 1
    16'b11111000_10001111 : OUT <= 1;  //248 / 143 = 1
    16'b11111000_10010000 : OUT <= 1;  //248 / 144 = 1
    16'b11111000_10010001 : OUT <= 1;  //248 / 145 = 1
    16'b11111000_10010010 : OUT <= 1;  //248 / 146 = 1
    16'b11111000_10010011 : OUT <= 1;  //248 / 147 = 1
    16'b11111000_10010100 : OUT <= 1;  //248 / 148 = 1
    16'b11111000_10010101 : OUT <= 1;  //248 / 149 = 1
    16'b11111000_10010110 : OUT <= 1;  //248 / 150 = 1
    16'b11111000_10010111 : OUT <= 1;  //248 / 151 = 1
    16'b11111000_10011000 : OUT <= 1;  //248 / 152 = 1
    16'b11111000_10011001 : OUT <= 1;  //248 / 153 = 1
    16'b11111000_10011010 : OUT <= 1;  //248 / 154 = 1
    16'b11111000_10011011 : OUT <= 1;  //248 / 155 = 1
    16'b11111000_10011100 : OUT <= 1;  //248 / 156 = 1
    16'b11111000_10011101 : OUT <= 1;  //248 / 157 = 1
    16'b11111000_10011110 : OUT <= 1;  //248 / 158 = 1
    16'b11111000_10011111 : OUT <= 1;  //248 / 159 = 1
    16'b11111000_10100000 : OUT <= 1;  //248 / 160 = 1
    16'b11111000_10100001 : OUT <= 1;  //248 / 161 = 1
    16'b11111000_10100010 : OUT <= 1;  //248 / 162 = 1
    16'b11111000_10100011 : OUT <= 1;  //248 / 163 = 1
    16'b11111000_10100100 : OUT <= 1;  //248 / 164 = 1
    16'b11111000_10100101 : OUT <= 1;  //248 / 165 = 1
    16'b11111000_10100110 : OUT <= 1;  //248 / 166 = 1
    16'b11111000_10100111 : OUT <= 1;  //248 / 167 = 1
    16'b11111000_10101000 : OUT <= 1;  //248 / 168 = 1
    16'b11111000_10101001 : OUT <= 1;  //248 / 169 = 1
    16'b11111000_10101010 : OUT <= 1;  //248 / 170 = 1
    16'b11111000_10101011 : OUT <= 1;  //248 / 171 = 1
    16'b11111000_10101100 : OUT <= 1;  //248 / 172 = 1
    16'b11111000_10101101 : OUT <= 1;  //248 / 173 = 1
    16'b11111000_10101110 : OUT <= 1;  //248 / 174 = 1
    16'b11111000_10101111 : OUT <= 1;  //248 / 175 = 1
    16'b11111000_10110000 : OUT <= 1;  //248 / 176 = 1
    16'b11111000_10110001 : OUT <= 1;  //248 / 177 = 1
    16'b11111000_10110010 : OUT <= 1;  //248 / 178 = 1
    16'b11111000_10110011 : OUT <= 1;  //248 / 179 = 1
    16'b11111000_10110100 : OUT <= 1;  //248 / 180 = 1
    16'b11111000_10110101 : OUT <= 1;  //248 / 181 = 1
    16'b11111000_10110110 : OUT <= 1;  //248 / 182 = 1
    16'b11111000_10110111 : OUT <= 1;  //248 / 183 = 1
    16'b11111000_10111000 : OUT <= 1;  //248 / 184 = 1
    16'b11111000_10111001 : OUT <= 1;  //248 / 185 = 1
    16'b11111000_10111010 : OUT <= 1;  //248 / 186 = 1
    16'b11111000_10111011 : OUT <= 1;  //248 / 187 = 1
    16'b11111000_10111100 : OUT <= 1;  //248 / 188 = 1
    16'b11111000_10111101 : OUT <= 1;  //248 / 189 = 1
    16'b11111000_10111110 : OUT <= 1;  //248 / 190 = 1
    16'b11111000_10111111 : OUT <= 1;  //248 / 191 = 1
    16'b11111000_11000000 : OUT <= 1;  //248 / 192 = 1
    16'b11111000_11000001 : OUT <= 1;  //248 / 193 = 1
    16'b11111000_11000010 : OUT <= 1;  //248 / 194 = 1
    16'b11111000_11000011 : OUT <= 1;  //248 / 195 = 1
    16'b11111000_11000100 : OUT <= 1;  //248 / 196 = 1
    16'b11111000_11000101 : OUT <= 1;  //248 / 197 = 1
    16'b11111000_11000110 : OUT <= 1;  //248 / 198 = 1
    16'b11111000_11000111 : OUT <= 1;  //248 / 199 = 1
    16'b11111000_11001000 : OUT <= 1;  //248 / 200 = 1
    16'b11111000_11001001 : OUT <= 1;  //248 / 201 = 1
    16'b11111000_11001010 : OUT <= 1;  //248 / 202 = 1
    16'b11111000_11001011 : OUT <= 1;  //248 / 203 = 1
    16'b11111000_11001100 : OUT <= 1;  //248 / 204 = 1
    16'b11111000_11001101 : OUT <= 1;  //248 / 205 = 1
    16'b11111000_11001110 : OUT <= 1;  //248 / 206 = 1
    16'b11111000_11001111 : OUT <= 1;  //248 / 207 = 1
    16'b11111000_11010000 : OUT <= 1;  //248 / 208 = 1
    16'b11111000_11010001 : OUT <= 1;  //248 / 209 = 1
    16'b11111000_11010010 : OUT <= 1;  //248 / 210 = 1
    16'b11111000_11010011 : OUT <= 1;  //248 / 211 = 1
    16'b11111000_11010100 : OUT <= 1;  //248 / 212 = 1
    16'b11111000_11010101 : OUT <= 1;  //248 / 213 = 1
    16'b11111000_11010110 : OUT <= 1;  //248 / 214 = 1
    16'b11111000_11010111 : OUT <= 1;  //248 / 215 = 1
    16'b11111000_11011000 : OUT <= 1;  //248 / 216 = 1
    16'b11111000_11011001 : OUT <= 1;  //248 / 217 = 1
    16'b11111000_11011010 : OUT <= 1;  //248 / 218 = 1
    16'b11111000_11011011 : OUT <= 1;  //248 / 219 = 1
    16'b11111000_11011100 : OUT <= 1;  //248 / 220 = 1
    16'b11111000_11011101 : OUT <= 1;  //248 / 221 = 1
    16'b11111000_11011110 : OUT <= 1;  //248 / 222 = 1
    16'b11111000_11011111 : OUT <= 1;  //248 / 223 = 1
    16'b11111000_11100000 : OUT <= 1;  //248 / 224 = 1
    16'b11111000_11100001 : OUT <= 1;  //248 / 225 = 1
    16'b11111000_11100010 : OUT <= 1;  //248 / 226 = 1
    16'b11111000_11100011 : OUT <= 1;  //248 / 227 = 1
    16'b11111000_11100100 : OUT <= 1;  //248 / 228 = 1
    16'b11111000_11100101 : OUT <= 1;  //248 / 229 = 1
    16'b11111000_11100110 : OUT <= 1;  //248 / 230 = 1
    16'b11111000_11100111 : OUT <= 1;  //248 / 231 = 1
    16'b11111000_11101000 : OUT <= 1;  //248 / 232 = 1
    16'b11111000_11101001 : OUT <= 1;  //248 / 233 = 1
    16'b11111000_11101010 : OUT <= 1;  //248 / 234 = 1
    16'b11111000_11101011 : OUT <= 1;  //248 / 235 = 1
    16'b11111000_11101100 : OUT <= 1;  //248 / 236 = 1
    16'b11111000_11101101 : OUT <= 1;  //248 / 237 = 1
    16'b11111000_11101110 : OUT <= 1;  //248 / 238 = 1
    16'b11111000_11101111 : OUT <= 1;  //248 / 239 = 1
    16'b11111000_11110000 : OUT <= 1;  //248 / 240 = 1
    16'b11111000_11110001 : OUT <= 1;  //248 / 241 = 1
    16'b11111000_11110010 : OUT <= 1;  //248 / 242 = 1
    16'b11111000_11110011 : OUT <= 1;  //248 / 243 = 1
    16'b11111000_11110100 : OUT <= 1;  //248 / 244 = 1
    16'b11111000_11110101 : OUT <= 1;  //248 / 245 = 1
    16'b11111000_11110110 : OUT <= 1;  //248 / 246 = 1
    16'b11111000_11110111 : OUT <= 1;  //248 / 247 = 1
    16'b11111000_11111000 : OUT <= 1;  //248 / 248 = 1
    16'b11111000_11111001 : OUT <= 0;  //248 / 249 = 0
    16'b11111000_11111010 : OUT <= 0;  //248 / 250 = 0
    16'b11111000_11111011 : OUT <= 0;  //248 / 251 = 0
    16'b11111000_11111100 : OUT <= 0;  //248 / 252 = 0
    16'b11111000_11111101 : OUT <= 0;  //248 / 253 = 0
    16'b11111000_11111110 : OUT <= 0;  //248 / 254 = 0
    16'b11111000_11111111 : OUT <= 0;  //248 / 255 = 0
    16'b11111001_00000000 : OUT <= 0;  //249 / 0 = 0
    16'b11111001_00000001 : OUT <= 249;  //249 / 1 = 249
    16'b11111001_00000010 : OUT <= 124;  //249 / 2 = 124
    16'b11111001_00000011 : OUT <= 83;  //249 / 3 = 83
    16'b11111001_00000100 : OUT <= 62;  //249 / 4 = 62
    16'b11111001_00000101 : OUT <= 49;  //249 / 5 = 49
    16'b11111001_00000110 : OUT <= 41;  //249 / 6 = 41
    16'b11111001_00000111 : OUT <= 35;  //249 / 7 = 35
    16'b11111001_00001000 : OUT <= 31;  //249 / 8 = 31
    16'b11111001_00001001 : OUT <= 27;  //249 / 9 = 27
    16'b11111001_00001010 : OUT <= 24;  //249 / 10 = 24
    16'b11111001_00001011 : OUT <= 22;  //249 / 11 = 22
    16'b11111001_00001100 : OUT <= 20;  //249 / 12 = 20
    16'b11111001_00001101 : OUT <= 19;  //249 / 13 = 19
    16'b11111001_00001110 : OUT <= 17;  //249 / 14 = 17
    16'b11111001_00001111 : OUT <= 16;  //249 / 15 = 16
    16'b11111001_00010000 : OUT <= 15;  //249 / 16 = 15
    16'b11111001_00010001 : OUT <= 14;  //249 / 17 = 14
    16'b11111001_00010010 : OUT <= 13;  //249 / 18 = 13
    16'b11111001_00010011 : OUT <= 13;  //249 / 19 = 13
    16'b11111001_00010100 : OUT <= 12;  //249 / 20 = 12
    16'b11111001_00010101 : OUT <= 11;  //249 / 21 = 11
    16'b11111001_00010110 : OUT <= 11;  //249 / 22 = 11
    16'b11111001_00010111 : OUT <= 10;  //249 / 23 = 10
    16'b11111001_00011000 : OUT <= 10;  //249 / 24 = 10
    16'b11111001_00011001 : OUT <= 9;  //249 / 25 = 9
    16'b11111001_00011010 : OUT <= 9;  //249 / 26 = 9
    16'b11111001_00011011 : OUT <= 9;  //249 / 27 = 9
    16'b11111001_00011100 : OUT <= 8;  //249 / 28 = 8
    16'b11111001_00011101 : OUT <= 8;  //249 / 29 = 8
    16'b11111001_00011110 : OUT <= 8;  //249 / 30 = 8
    16'b11111001_00011111 : OUT <= 8;  //249 / 31 = 8
    16'b11111001_00100000 : OUT <= 7;  //249 / 32 = 7
    16'b11111001_00100001 : OUT <= 7;  //249 / 33 = 7
    16'b11111001_00100010 : OUT <= 7;  //249 / 34 = 7
    16'b11111001_00100011 : OUT <= 7;  //249 / 35 = 7
    16'b11111001_00100100 : OUT <= 6;  //249 / 36 = 6
    16'b11111001_00100101 : OUT <= 6;  //249 / 37 = 6
    16'b11111001_00100110 : OUT <= 6;  //249 / 38 = 6
    16'b11111001_00100111 : OUT <= 6;  //249 / 39 = 6
    16'b11111001_00101000 : OUT <= 6;  //249 / 40 = 6
    16'b11111001_00101001 : OUT <= 6;  //249 / 41 = 6
    16'b11111001_00101010 : OUT <= 5;  //249 / 42 = 5
    16'b11111001_00101011 : OUT <= 5;  //249 / 43 = 5
    16'b11111001_00101100 : OUT <= 5;  //249 / 44 = 5
    16'b11111001_00101101 : OUT <= 5;  //249 / 45 = 5
    16'b11111001_00101110 : OUT <= 5;  //249 / 46 = 5
    16'b11111001_00101111 : OUT <= 5;  //249 / 47 = 5
    16'b11111001_00110000 : OUT <= 5;  //249 / 48 = 5
    16'b11111001_00110001 : OUT <= 5;  //249 / 49 = 5
    16'b11111001_00110010 : OUT <= 4;  //249 / 50 = 4
    16'b11111001_00110011 : OUT <= 4;  //249 / 51 = 4
    16'b11111001_00110100 : OUT <= 4;  //249 / 52 = 4
    16'b11111001_00110101 : OUT <= 4;  //249 / 53 = 4
    16'b11111001_00110110 : OUT <= 4;  //249 / 54 = 4
    16'b11111001_00110111 : OUT <= 4;  //249 / 55 = 4
    16'b11111001_00111000 : OUT <= 4;  //249 / 56 = 4
    16'b11111001_00111001 : OUT <= 4;  //249 / 57 = 4
    16'b11111001_00111010 : OUT <= 4;  //249 / 58 = 4
    16'b11111001_00111011 : OUT <= 4;  //249 / 59 = 4
    16'b11111001_00111100 : OUT <= 4;  //249 / 60 = 4
    16'b11111001_00111101 : OUT <= 4;  //249 / 61 = 4
    16'b11111001_00111110 : OUT <= 4;  //249 / 62 = 4
    16'b11111001_00111111 : OUT <= 3;  //249 / 63 = 3
    16'b11111001_01000000 : OUT <= 3;  //249 / 64 = 3
    16'b11111001_01000001 : OUT <= 3;  //249 / 65 = 3
    16'b11111001_01000010 : OUT <= 3;  //249 / 66 = 3
    16'b11111001_01000011 : OUT <= 3;  //249 / 67 = 3
    16'b11111001_01000100 : OUT <= 3;  //249 / 68 = 3
    16'b11111001_01000101 : OUT <= 3;  //249 / 69 = 3
    16'b11111001_01000110 : OUT <= 3;  //249 / 70 = 3
    16'b11111001_01000111 : OUT <= 3;  //249 / 71 = 3
    16'b11111001_01001000 : OUT <= 3;  //249 / 72 = 3
    16'b11111001_01001001 : OUT <= 3;  //249 / 73 = 3
    16'b11111001_01001010 : OUT <= 3;  //249 / 74 = 3
    16'b11111001_01001011 : OUT <= 3;  //249 / 75 = 3
    16'b11111001_01001100 : OUT <= 3;  //249 / 76 = 3
    16'b11111001_01001101 : OUT <= 3;  //249 / 77 = 3
    16'b11111001_01001110 : OUT <= 3;  //249 / 78 = 3
    16'b11111001_01001111 : OUT <= 3;  //249 / 79 = 3
    16'b11111001_01010000 : OUT <= 3;  //249 / 80 = 3
    16'b11111001_01010001 : OUT <= 3;  //249 / 81 = 3
    16'b11111001_01010010 : OUT <= 3;  //249 / 82 = 3
    16'b11111001_01010011 : OUT <= 3;  //249 / 83 = 3
    16'b11111001_01010100 : OUT <= 2;  //249 / 84 = 2
    16'b11111001_01010101 : OUT <= 2;  //249 / 85 = 2
    16'b11111001_01010110 : OUT <= 2;  //249 / 86 = 2
    16'b11111001_01010111 : OUT <= 2;  //249 / 87 = 2
    16'b11111001_01011000 : OUT <= 2;  //249 / 88 = 2
    16'b11111001_01011001 : OUT <= 2;  //249 / 89 = 2
    16'b11111001_01011010 : OUT <= 2;  //249 / 90 = 2
    16'b11111001_01011011 : OUT <= 2;  //249 / 91 = 2
    16'b11111001_01011100 : OUT <= 2;  //249 / 92 = 2
    16'b11111001_01011101 : OUT <= 2;  //249 / 93 = 2
    16'b11111001_01011110 : OUT <= 2;  //249 / 94 = 2
    16'b11111001_01011111 : OUT <= 2;  //249 / 95 = 2
    16'b11111001_01100000 : OUT <= 2;  //249 / 96 = 2
    16'b11111001_01100001 : OUT <= 2;  //249 / 97 = 2
    16'b11111001_01100010 : OUT <= 2;  //249 / 98 = 2
    16'b11111001_01100011 : OUT <= 2;  //249 / 99 = 2
    16'b11111001_01100100 : OUT <= 2;  //249 / 100 = 2
    16'b11111001_01100101 : OUT <= 2;  //249 / 101 = 2
    16'b11111001_01100110 : OUT <= 2;  //249 / 102 = 2
    16'b11111001_01100111 : OUT <= 2;  //249 / 103 = 2
    16'b11111001_01101000 : OUT <= 2;  //249 / 104 = 2
    16'b11111001_01101001 : OUT <= 2;  //249 / 105 = 2
    16'b11111001_01101010 : OUT <= 2;  //249 / 106 = 2
    16'b11111001_01101011 : OUT <= 2;  //249 / 107 = 2
    16'b11111001_01101100 : OUT <= 2;  //249 / 108 = 2
    16'b11111001_01101101 : OUT <= 2;  //249 / 109 = 2
    16'b11111001_01101110 : OUT <= 2;  //249 / 110 = 2
    16'b11111001_01101111 : OUT <= 2;  //249 / 111 = 2
    16'b11111001_01110000 : OUT <= 2;  //249 / 112 = 2
    16'b11111001_01110001 : OUT <= 2;  //249 / 113 = 2
    16'b11111001_01110010 : OUT <= 2;  //249 / 114 = 2
    16'b11111001_01110011 : OUT <= 2;  //249 / 115 = 2
    16'b11111001_01110100 : OUT <= 2;  //249 / 116 = 2
    16'b11111001_01110101 : OUT <= 2;  //249 / 117 = 2
    16'b11111001_01110110 : OUT <= 2;  //249 / 118 = 2
    16'b11111001_01110111 : OUT <= 2;  //249 / 119 = 2
    16'b11111001_01111000 : OUT <= 2;  //249 / 120 = 2
    16'b11111001_01111001 : OUT <= 2;  //249 / 121 = 2
    16'b11111001_01111010 : OUT <= 2;  //249 / 122 = 2
    16'b11111001_01111011 : OUT <= 2;  //249 / 123 = 2
    16'b11111001_01111100 : OUT <= 2;  //249 / 124 = 2
    16'b11111001_01111101 : OUT <= 1;  //249 / 125 = 1
    16'b11111001_01111110 : OUT <= 1;  //249 / 126 = 1
    16'b11111001_01111111 : OUT <= 1;  //249 / 127 = 1
    16'b11111001_10000000 : OUT <= 1;  //249 / 128 = 1
    16'b11111001_10000001 : OUT <= 1;  //249 / 129 = 1
    16'b11111001_10000010 : OUT <= 1;  //249 / 130 = 1
    16'b11111001_10000011 : OUT <= 1;  //249 / 131 = 1
    16'b11111001_10000100 : OUT <= 1;  //249 / 132 = 1
    16'b11111001_10000101 : OUT <= 1;  //249 / 133 = 1
    16'b11111001_10000110 : OUT <= 1;  //249 / 134 = 1
    16'b11111001_10000111 : OUT <= 1;  //249 / 135 = 1
    16'b11111001_10001000 : OUT <= 1;  //249 / 136 = 1
    16'b11111001_10001001 : OUT <= 1;  //249 / 137 = 1
    16'b11111001_10001010 : OUT <= 1;  //249 / 138 = 1
    16'b11111001_10001011 : OUT <= 1;  //249 / 139 = 1
    16'b11111001_10001100 : OUT <= 1;  //249 / 140 = 1
    16'b11111001_10001101 : OUT <= 1;  //249 / 141 = 1
    16'b11111001_10001110 : OUT <= 1;  //249 / 142 = 1
    16'b11111001_10001111 : OUT <= 1;  //249 / 143 = 1
    16'b11111001_10010000 : OUT <= 1;  //249 / 144 = 1
    16'b11111001_10010001 : OUT <= 1;  //249 / 145 = 1
    16'b11111001_10010010 : OUT <= 1;  //249 / 146 = 1
    16'b11111001_10010011 : OUT <= 1;  //249 / 147 = 1
    16'b11111001_10010100 : OUT <= 1;  //249 / 148 = 1
    16'b11111001_10010101 : OUT <= 1;  //249 / 149 = 1
    16'b11111001_10010110 : OUT <= 1;  //249 / 150 = 1
    16'b11111001_10010111 : OUT <= 1;  //249 / 151 = 1
    16'b11111001_10011000 : OUT <= 1;  //249 / 152 = 1
    16'b11111001_10011001 : OUT <= 1;  //249 / 153 = 1
    16'b11111001_10011010 : OUT <= 1;  //249 / 154 = 1
    16'b11111001_10011011 : OUT <= 1;  //249 / 155 = 1
    16'b11111001_10011100 : OUT <= 1;  //249 / 156 = 1
    16'b11111001_10011101 : OUT <= 1;  //249 / 157 = 1
    16'b11111001_10011110 : OUT <= 1;  //249 / 158 = 1
    16'b11111001_10011111 : OUT <= 1;  //249 / 159 = 1
    16'b11111001_10100000 : OUT <= 1;  //249 / 160 = 1
    16'b11111001_10100001 : OUT <= 1;  //249 / 161 = 1
    16'b11111001_10100010 : OUT <= 1;  //249 / 162 = 1
    16'b11111001_10100011 : OUT <= 1;  //249 / 163 = 1
    16'b11111001_10100100 : OUT <= 1;  //249 / 164 = 1
    16'b11111001_10100101 : OUT <= 1;  //249 / 165 = 1
    16'b11111001_10100110 : OUT <= 1;  //249 / 166 = 1
    16'b11111001_10100111 : OUT <= 1;  //249 / 167 = 1
    16'b11111001_10101000 : OUT <= 1;  //249 / 168 = 1
    16'b11111001_10101001 : OUT <= 1;  //249 / 169 = 1
    16'b11111001_10101010 : OUT <= 1;  //249 / 170 = 1
    16'b11111001_10101011 : OUT <= 1;  //249 / 171 = 1
    16'b11111001_10101100 : OUT <= 1;  //249 / 172 = 1
    16'b11111001_10101101 : OUT <= 1;  //249 / 173 = 1
    16'b11111001_10101110 : OUT <= 1;  //249 / 174 = 1
    16'b11111001_10101111 : OUT <= 1;  //249 / 175 = 1
    16'b11111001_10110000 : OUT <= 1;  //249 / 176 = 1
    16'b11111001_10110001 : OUT <= 1;  //249 / 177 = 1
    16'b11111001_10110010 : OUT <= 1;  //249 / 178 = 1
    16'b11111001_10110011 : OUT <= 1;  //249 / 179 = 1
    16'b11111001_10110100 : OUT <= 1;  //249 / 180 = 1
    16'b11111001_10110101 : OUT <= 1;  //249 / 181 = 1
    16'b11111001_10110110 : OUT <= 1;  //249 / 182 = 1
    16'b11111001_10110111 : OUT <= 1;  //249 / 183 = 1
    16'b11111001_10111000 : OUT <= 1;  //249 / 184 = 1
    16'b11111001_10111001 : OUT <= 1;  //249 / 185 = 1
    16'b11111001_10111010 : OUT <= 1;  //249 / 186 = 1
    16'b11111001_10111011 : OUT <= 1;  //249 / 187 = 1
    16'b11111001_10111100 : OUT <= 1;  //249 / 188 = 1
    16'b11111001_10111101 : OUT <= 1;  //249 / 189 = 1
    16'b11111001_10111110 : OUT <= 1;  //249 / 190 = 1
    16'b11111001_10111111 : OUT <= 1;  //249 / 191 = 1
    16'b11111001_11000000 : OUT <= 1;  //249 / 192 = 1
    16'b11111001_11000001 : OUT <= 1;  //249 / 193 = 1
    16'b11111001_11000010 : OUT <= 1;  //249 / 194 = 1
    16'b11111001_11000011 : OUT <= 1;  //249 / 195 = 1
    16'b11111001_11000100 : OUT <= 1;  //249 / 196 = 1
    16'b11111001_11000101 : OUT <= 1;  //249 / 197 = 1
    16'b11111001_11000110 : OUT <= 1;  //249 / 198 = 1
    16'b11111001_11000111 : OUT <= 1;  //249 / 199 = 1
    16'b11111001_11001000 : OUT <= 1;  //249 / 200 = 1
    16'b11111001_11001001 : OUT <= 1;  //249 / 201 = 1
    16'b11111001_11001010 : OUT <= 1;  //249 / 202 = 1
    16'b11111001_11001011 : OUT <= 1;  //249 / 203 = 1
    16'b11111001_11001100 : OUT <= 1;  //249 / 204 = 1
    16'b11111001_11001101 : OUT <= 1;  //249 / 205 = 1
    16'b11111001_11001110 : OUT <= 1;  //249 / 206 = 1
    16'b11111001_11001111 : OUT <= 1;  //249 / 207 = 1
    16'b11111001_11010000 : OUT <= 1;  //249 / 208 = 1
    16'b11111001_11010001 : OUT <= 1;  //249 / 209 = 1
    16'b11111001_11010010 : OUT <= 1;  //249 / 210 = 1
    16'b11111001_11010011 : OUT <= 1;  //249 / 211 = 1
    16'b11111001_11010100 : OUT <= 1;  //249 / 212 = 1
    16'b11111001_11010101 : OUT <= 1;  //249 / 213 = 1
    16'b11111001_11010110 : OUT <= 1;  //249 / 214 = 1
    16'b11111001_11010111 : OUT <= 1;  //249 / 215 = 1
    16'b11111001_11011000 : OUT <= 1;  //249 / 216 = 1
    16'b11111001_11011001 : OUT <= 1;  //249 / 217 = 1
    16'b11111001_11011010 : OUT <= 1;  //249 / 218 = 1
    16'b11111001_11011011 : OUT <= 1;  //249 / 219 = 1
    16'b11111001_11011100 : OUT <= 1;  //249 / 220 = 1
    16'b11111001_11011101 : OUT <= 1;  //249 / 221 = 1
    16'b11111001_11011110 : OUT <= 1;  //249 / 222 = 1
    16'b11111001_11011111 : OUT <= 1;  //249 / 223 = 1
    16'b11111001_11100000 : OUT <= 1;  //249 / 224 = 1
    16'b11111001_11100001 : OUT <= 1;  //249 / 225 = 1
    16'b11111001_11100010 : OUT <= 1;  //249 / 226 = 1
    16'b11111001_11100011 : OUT <= 1;  //249 / 227 = 1
    16'b11111001_11100100 : OUT <= 1;  //249 / 228 = 1
    16'b11111001_11100101 : OUT <= 1;  //249 / 229 = 1
    16'b11111001_11100110 : OUT <= 1;  //249 / 230 = 1
    16'b11111001_11100111 : OUT <= 1;  //249 / 231 = 1
    16'b11111001_11101000 : OUT <= 1;  //249 / 232 = 1
    16'b11111001_11101001 : OUT <= 1;  //249 / 233 = 1
    16'b11111001_11101010 : OUT <= 1;  //249 / 234 = 1
    16'b11111001_11101011 : OUT <= 1;  //249 / 235 = 1
    16'b11111001_11101100 : OUT <= 1;  //249 / 236 = 1
    16'b11111001_11101101 : OUT <= 1;  //249 / 237 = 1
    16'b11111001_11101110 : OUT <= 1;  //249 / 238 = 1
    16'b11111001_11101111 : OUT <= 1;  //249 / 239 = 1
    16'b11111001_11110000 : OUT <= 1;  //249 / 240 = 1
    16'b11111001_11110001 : OUT <= 1;  //249 / 241 = 1
    16'b11111001_11110010 : OUT <= 1;  //249 / 242 = 1
    16'b11111001_11110011 : OUT <= 1;  //249 / 243 = 1
    16'b11111001_11110100 : OUT <= 1;  //249 / 244 = 1
    16'b11111001_11110101 : OUT <= 1;  //249 / 245 = 1
    16'b11111001_11110110 : OUT <= 1;  //249 / 246 = 1
    16'b11111001_11110111 : OUT <= 1;  //249 / 247 = 1
    16'b11111001_11111000 : OUT <= 1;  //249 / 248 = 1
    16'b11111001_11111001 : OUT <= 1;  //249 / 249 = 1
    16'b11111001_11111010 : OUT <= 0;  //249 / 250 = 0
    16'b11111001_11111011 : OUT <= 0;  //249 / 251 = 0
    16'b11111001_11111100 : OUT <= 0;  //249 / 252 = 0
    16'b11111001_11111101 : OUT <= 0;  //249 / 253 = 0
    16'b11111001_11111110 : OUT <= 0;  //249 / 254 = 0
    16'b11111001_11111111 : OUT <= 0;  //249 / 255 = 0
    16'b11111010_00000000 : OUT <= 0;  //250 / 0 = 0
    16'b11111010_00000001 : OUT <= 250;  //250 / 1 = 250
    16'b11111010_00000010 : OUT <= 125;  //250 / 2 = 125
    16'b11111010_00000011 : OUT <= 83;  //250 / 3 = 83
    16'b11111010_00000100 : OUT <= 62;  //250 / 4 = 62
    16'b11111010_00000101 : OUT <= 50;  //250 / 5 = 50
    16'b11111010_00000110 : OUT <= 41;  //250 / 6 = 41
    16'b11111010_00000111 : OUT <= 35;  //250 / 7 = 35
    16'b11111010_00001000 : OUT <= 31;  //250 / 8 = 31
    16'b11111010_00001001 : OUT <= 27;  //250 / 9 = 27
    16'b11111010_00001010 : OUT <= 25;  //250 / 10 = 25
    16'b11111010_00001011 : OUT <= 22;  //250 / 11 = 22
    16'b11111010_00001100 : OUT <= 20;  //250 / 12 = 20
    16'b11111010_00001101 : OUT <= 19;  //250 / 13 = 19
    16'b11111010_00001110 : OUT <= 17;  //250 / 14 = 17
    16'b11111010_00001111 : OUT <= 16;  //250 / 15 = 16
    16'b11111010_00010000 : OUT <= 15;  //250 / 16 = 15
    16'b11111010_00010001 : OUT <= 14;  //250 / 17 = 14
    16'b11111010_00010010 : OUT <= 13;  //250 / 18 = 13
    16'b11111010_00010011 : OUT <= 13;  //250 / 19 = 13
    16'b11111010_00010100 : OUT <= 12;  //250 / 20 = 12
    16'b11111010_00010101 : OUT <= 11;  //250 / 21 = 11
    16'b11111010_00010110 : OUT <= 11;  //250 / 22 = 11
    16'b11111010_00010111 : OUT <= 10;  //250 / 23 = 10
    16'b11111010_00011000 : OUT <= 10;  //250 / 24 = 10
    16'b11111010_00011001 : OUT <= 10;  //250 / 25 = 10
    16'b11111010_00011010 : OUT <= 9;  //250 / 26 = 9
    16'b11111010_00011011 : OUT <= 9;  //250 / 27 = 9
    16'b11111010_00011100 : OUT <= 8;  //250 / 28 = 8
    16'b11111010_00011101 : OUT <= 8;  //250 / 29 = 8
    16'b11111010_00011110 : OUT <= 8;  //250 / 30 = 8
    16'b11111010_00011111 : OUT <= 8;  //250 / 31 = 8
    16'b11111010_00100000 : OUT <= 7;  //250 / 32 = 7
    16'b11111010_00100001 : OUT <= 7;  //250 / 33 = 7
    16'b11111010_00100010 : OUT <= 7;  //250 / 34 = 7
    16'b11111010_00100011 : OUT <= 7;  //250 / 35 = 7
    16'b11111010_00100100 : OUT <= 6;  //250 / 36 = 6
    16'b11111010_00100101 : OUT <= 6;  //250 / 37 = 6
    16'b11111010_00100110 : OUT <= 6;  //250 / 38 = 6
    16'b11111010_00100111 : OUT <= 6;  //250 / 39 = 6
    16'b11111010_00101000 : OUT <= 6;  //250 / 40 = 6
    16'b11111010_00101001 : OUT <= 6;  //250 / 41 = 6
    16'b11111010_00101010 : OUT <= 5;  //250 / 42 = 5
    16'b11111010_00101011 : OUT <= 5;  //250 / 43 = 5
    16'b11111010_00101100 : OUT <= 5;  //250 / 44 = 5
    16'b11111010_00101101 : OUT <= 5;  //250 / 45 = 5
    16'b11111010_00101110 : OUT <= 5;  //250 / 46 = 5
    16'b11111010_00101111 : OUT <= 5;  //250 / 47 = 5
    16'b11111010_00110000 : OUT <= 5;  //250 / 48 = 5
    16'b11111010_00110001 : OUT <= 5;  //250 / 49 = 5
    16'b11111010_00110010 : OUT <= 5;  //250 / 50 = 5
    16'b11111010_00110011 : OUT <= 4;  //250 / 51 = 4
    16'b11111010_00110100 : OUT <= 4;  //250 / 52 = 4
    16'b11111010_00110101 : OUT <= 4;  //250 / 53 = 4
    16'b11111010_00110110 : OUT <= 4;  //250 / 54 = 4
    16'b11111010_00110111 : OUT <= 4;  //250 / 55 = 4
    16'b11111010_00111000 : OUT <= 4;  //250 / 56 = 4
    16'b11111010_00111001 : OUT <= 4;  //250 / 57 = 4
    16'b11111010_00111010 : OUT <= 4;  //250 / 58 = 4
    16'b11111010_00111011 : OUT <= 4;  //250 / 59 = 4
    16'b11111010_00111100 : OUT <= 4;  //250 / 60 = 4
    16'b11111010_00111101 : OUT <= 4;  //250 / 61 = 4
    16'b11111010_00111110 : OUT <= 4;  //250 / 62 = 4
    16'b11111010_00111111 : OUT <= 3;  //250 / 63 = 3
    16'b11111010_01000000 : OUT <= 3;  //250 / 64 = 3
    16'b11111010_01000001 : OUT <= 3;  //250 / 65 = 3
    16'b11111010_01000010 : OUT <= 3;  //250 / 66 = 3
    16'b11111010_01000011 : OUT <= 3;  //250 / 67 = 3
    16'b11111010_01000100 : OUT <= 3;  //250 / 68 = 3
    16'b11111010_01000101 : OUT <= 3;  //250 / 69 = 3
    16'b11111010_01000110 : OUT <= 3;  //250 / 70 = 3
    16'b11111010_01000111 : OUT <= 3;  //250 / 71 = 3
    16'b11111010_01001000 : OUT <= 3;  //250 / 72 = 3
    16'b11111010_01001001 : OUT <= 3;  //250 / 73 = 3
    16'b11111010_01001010 : OUT <= 3;  //250 / 74 = 3
    16'b11111010_01001011 : OUT <= 3;  //250 / 75 = 3
    16'b11111010_01001100 : OUT <= 3;  //250 / 76 = 3
    16'b11111010_01001101 : OUT <= 3;  //250 / 77 = 3
    16'b11111010_01001110 : OUT <= 3;  //250 / 78 = 3
    16'b11111010_01001111 : OUT <= 3;  //250 / 79 = 3
    16'b11111010_01010000 : OUT <= 3;  //250 / 80 = 3
    16'b11111010_01010001 : OUT <= 3;  //250 / 81 = 3
    16'b11111010_01010010 : OUT <= 3;  //250 / 82 = 3
    16'b11111010_01010011 : OUT <= 3;  //250 / 83 = 3
    16'b11111010_01010100 : OUT <= 2;  //250 / 84 = 2
    16'b11111010_01010101 : OUT <= 2;  //250 / 85 = 2
    16'b11111010_01010110 : OUT <= 2;  //250 / 86 = 2
    16'b11111010_01010111 : OUT <= 2;  //250 / 87 = 2
    16'b11111010_01011000 : OUT <= 2;  //250 / 88 = 2
    16'b11111010_01011001 : OUT <= 2;  //250 / 89 = 2
    16'b11111010_01011010 : OUT <= 2;  //250 / 90 = 2
    16'b11111010_01011011 : OUT <= 2;  //250 / 91 = 2
    16'b11111010_01011100 : OUT <= 2;  //250 / 92 = 2
    16'b11111010_01011101 : OUT <= 2;  //250 / 93 = 2
    16'b11111010_01011110 : OUT <= 2;  //250 / 94 = 2
    16'b11111010_01011111 : OUT <= 2;  //250 / 95 = 2
    16'b11111010_01100000 : OUT <= 2;  //250 / 96 = 2
    16'b11111010_01100001 : OUT <= 2;  //250 / 97 = 2
    16'b11111010_01100010 : OUT <= 2;  //250 / 98 = 2
    16'b11111010_01100011 : OUT <= 2;  //250 / 99 = 2
    16'b11111010_01100100 : OUT <= 2;  //250 / 100 = 2
    16'b11111010_01100101 : OUT <= 2;  //250 / 101 = 2
    16'b11111010_01100110 : OUT <= 2;  //250 / 102 = 2
    16'b11111010_01100111 : OUT <= 2;  //250 / 103 = 2
    16'b11111010_01101000 : OUT <= 2;  //250 / 104 = 2
    16'b11111010_01101001 : OUT <= 2;  //250 / 105 = 2
    16'b11111010_01101010 : OUT <= 2;  //250 / 106 = 2
    16'b11111010_01101011 : OUT <= 2;  //250 / 107 = 2
    16'b11111010_01101100 : OUT <= 2;  //250 / 108 = 2
    16'b11111010_01101101 : OUT <= 2;  //250 / 109 = 2
    16'b11111010_01101110 : OUT <= 2;  //250 / 110 = 2
    16'b11111010_01101111 : OUT <= 2;  //250 / 111 = 2
    16'b11111010_01110000 : OUT <= 2;  //250 / 112 = 2
    16'b11111010_01110001 : OUT <= 2;  //250 / 113 = 2
    16'b11111010_01110010 : OUT <= 2;  //250 / 114 = 2
    16'b11111010_01110011 : OUT <= 2;  //250 / 115 = 2
    16'b11111010_01110100 : OUT <= 2;  //250 / 116 = 2
    16'b11111010_01110101 : OUT <= 2;  //250 / 117 = 2
    16'b11111010_01110110 : OUT <= 2;  //250 / 118 = 2
    16'b11111010_01110111 : OUT <= 2;  //250 / 119 = 2
    16'b11111010_01111000 : OUT <= 2;  //250 / 120 = 2
    16'b11111010_01111001 : OUT <= 2;  //250 / 121 = 2
    16'b11111010_01111010 : OUT <= 2;  //250 / 122 = 2
    16'b11111010_01111011 : OUT <= 2;  //250 / 123 = 2
    16'b11111010_01111100 : OUT <= 2;  //250 / 124 = 2
    16'b11111010_01111101 : OUT <= 2;  //250 / 125 = 2
    16'b11111010_01111110 : OUT <= 1;  //250 / 126 = 1
    16'b11111010_01111111 : OUT <= 1;  //250 / 127 = 1
    16'b11111010_10000000 : OUT <= 1;  //250 / 128 = 1
    16'b11111010_10000001 : OUT <= 1;  //250 / 129 = 1
    16'b11111010_10000010 : OUT <= 1;  //250 / 130 = 1
    16'b11111010_10000011 : OUT <= 1;  //250 / 131 = 1
    16'b11111010_10000100 : OUT <= 1;  //250 / 132 = 1
    16'b11111010_10000101 : OUT <= 1;  //250 / 133 = 1
    16'b11111010_10000110 : OUT <= 1;  //250 / 134 = 1
    16'b11111010_10000111 : OUT <= 1;  //250 / 135 = 1
    16'b11111010_10001000 : OUT <= 1;  //250 / 136 = 1
    16'b11111010_10001001 : OUT <= 1;  //250 / 137 = 1
    16'b11111010_10001010 : OUT <= 1;  //250 / 138 = 1
    16'b11111010_10001011 : OUT <= 1;  //250 / 139 = 1
    16'b11111010_10001100 : OUT <= 1;  //250 / 140 = 1
    16'b11111010_10001101 : OUT <= 1;  //250 / 141 = 1
    16'b11111010_10001110 : OUT <= 1;  //250 / 142 = 1
    16'b11111010_10001111 : OUT <= 1;  //250 / 143 = 1
    16'b11111010_10010000 : OUT <= 1;  //250 / 144 = 1
    16'b11111010_10010001 : OUT <= 1;  //250 / 145 = 1
    16'b11111010_10010010 : OUT <= 1;  //250 / 146 = 1
    16'b11111010_10010011 : OUT <= 1;  //250 / 147 = 1
    16'b11111010_10010100 : OUT <= 1;  //250 / 148 = 1
    16'b11111010_10010101 : OUT <= 1;  //250 / 149 = 1
    16'b11111010_10010110 : OUT <= 1;  //250 / 150 = 1
    16'b11111010_10010111 : OUT <= 1;  //250 / 151 = 1
    16'b11111010_10011000 : OUT <= 1;  //250 / 152 = 1
    16'b11111010_10011001 : OUT <= 1;  //250 / 153 = 1
    16'b11111010_10011010 : OUT <= 1;  //250 / 154 = 1
    16'b11111010_10011011 : OUT <= 1;  //250 / 155 = 1
    16'b11111010_10011100 : OUT <= 1;  //250 / 156 = 1
    16'b11111010_10011101 : OUT <= 1;  //250 / 157 = 1
    16'b11111010_10011110 : OUT <= 1;  //250 / 158 = 1
    16'b11111010_10011111 : OUT <= 1;  //250 / 159 = 1
    16'b11111010_10100000 : OUT <= 1;  //250 / 160 = 1
    16'b11111010_10100001 : OUT <= 1;  //250 / 161 = 1
    16'b11111010_10100010 : OUT <= 1;  //250 / 162 = 1
    16'b11111010_10100011 : OUT <= 1;  //250 / 163 = 1
    16'b11111010_10100100 : OUT <= 1;  //250 / 164 = 1
    16'b11111010_10100101 : OUT <= 1;  //250 / 165 = 1
    16'b11111010_10100110 : OUT <= 1;  //250 / 166 = 1
    16'b11111010_10100111 : OUT <= 1;  //250 / 167 = 1
    16'b11111010_10101000 : OUT <= 1;  //250 / 168 = 1
    16'b11111010_10101001 : OUT <= 1;  //250 / 169 = 1
    16'b11111010_10101010 : OUT <= 1;  //250 / 170 = 1
    16'b11111010_10101011 : OUT <= 1;  //250 / 171 = 1
    16'b11111010_10101100 : OUT <= 1;  //250 / 172 = 1
    16'b11111010_10101101 : OUT <= 1;  //250 / 173 = 1
    16'b11111010_10101110 : OUT <= 1;  //250 / 174 = 1
    16'b11111010_10101111 : OUT <= 1;  //250 / 175 = 1
    16'b11111010_10110000 : OUT <= 1;  //250 / 176 = 1
    16'b11111010_10110001 : OUT <= 1;  //250 / 177 = 1
    16'b11111010_10110010 : OUT <= 1;  //250 / 178 = 1
    16'b11111010_10110011 : OUT <= 1;  //250 / 179 = 1
    16'b11111010_10110100 : OUT <= 1;  //250 / 180 = 1
    16'b11111010_10110101 : OUT <= 1;  //250 / 181 = 1
    16'b11111010_10110110 : OUT <= 1;  //250 / 182 = 1
    16'b11111010_10110111 : OUT <= 1;  //250 / 183 = 1
    16'b11111010_10111000 : OUT <= 1;  //250 / 184 = 1
    16'b11111010_10111001 : OUT <= 1;  //250 / 185 = 1
    16'b11111010_10111010 : OUT <= 1;  //250 / 186 = 1
    16'b11111010_10111011 : OUT <= 1;  //250 / 187 = 1
    16'b11111010_10111100 : OUT <= 1;  //250 / 188 = 1
    16'b11111010_10111101 : OUT <= 1;  //250 / 189 = 1
    16'b11111010_10111110 : OUT <= 1;  //250 / 190 = 1
    16'b11111010_10111111 : OUT <= 1;  //250 / 191 = 1
    16'b11111010_11000000 : OUT <= 1;  //250 / 192 = 1
    16'b11111010_11000001 : OUT <= 1;  //250 / 193 = 1
    16'b11111010_11000010 : OUT <= 1;  //250 / 194 = 1
    16'b11111010_11000011 : OUT <= 1;  //250 / 195 = 1
    16'b11111010_11000100 : OUT <= 1;  //250 / 196 = 1
    16'b11111010_11000101 : OUT <= 1;  //250 / 197 = 1
    16'b11111010_11000110 : OUT <= 1;  //250 / 198 = 1
    16'b11111010_11000111 : OUT <= 1;  //250 / 199 = 1
    16'b11111010_11001000 : OUT <= 1;  //250 / 200 = 1
    16'b11111010_11001001 : OUT <= 1;  //250 / 201 = 1
    16'b11111010_11001010 : OUT <= 1;  //250 / 202 = 1
    16'b11111010_11001011 : OUT <= 1;  //250 / 203 = 1
    16'b11111010_11001100 : OUT <= 1;  //250 / 204 = 1
    16'b11111010_11001101 : OUT <= 1;  //250 / 205 = 1
    16'b11111010_11001110 : OUT <= 1;  //250 / 206 = 1
    16'b11111010_11001111 : OUT <= 1;  //250 / 207 = 1
    16'b11111010_11010000 : OUT <= 1;  //250 / 208 = 1
    16'b11111010_11010001 : OUT <= 1;  //250 / 209 = 1
    16'b11111010_11010010 : OUT <= 1;  //250 / 210 = 1
    16'b11111010_11010011 : OUT <= 1;  //250 / 211 = 1
    16'b11111010_11010100 : OUT <= 1;  //250 / 212 = 1
    16'b11111010_11010101 : OUT <= 1;  //250 / 213 = 1
    16'b11111010_11010110 : OUT <= 1;  //250 / 214 = 1
    16'b11111010_11010111 : OUT <= 1;  //250 / 215 = 1
    16'b11111010_11011000 : OUT <= 1;  //250 / 216 = 1
    16'b11111010_11011001 : OUT <= 1;  //250 / 217 = 1
    16'b11111010_11011010 : OUT <= 1;  //250 / 218 = 1
    16'b11111010_11011011 : OUT <= 1;  //250 / 219 = 1
    16'b11111010_11011100 : OUT <= 1;  //250 / 220 = 1
    16'b11111010_11011101 : OUT <= 1;  //250 / 221 = 1
    16'b11111010_11011110 : OUT <= 1;  //250 / 222 = 1
    16'b11111010_11011111 : OUT <= 1;  //250 / 223 = 1
    16'b11111010_11100000 : OUT <= 1;  //250 / 224 = 1
    16'b11111010_11100001 : OUT <= 1;  //250 / 225 = 1
    16'b11111010_11100010 : OUT <= 1;  //250 / 226 = 1
    16'b11111010_11100011 : OUT <= 1;  //250 / 227 = 1
    16'b11111010_11100100 : OUT <= 1;  //250 / 228 = 1
    16'b11111010_11100101 : OUT <= 1;  //250 / 229 = 1
    16'b11111010_11100110 : OUT <= 1;  //250 / 230 = 1
    16'b11111010_11100111 : OUT <= 1;  //250 / 231 = 1
    16'b11111010_11101000 : OUT <= 1;  //250 / 232 = 1
    16'b11111010_11101001 : OUT <= 1;  //250 / 233 = 1
    16'b11111010_11101010 : OUT <= 1;  //250 / 234 = 1
    16'b11111010_11101011 : OUT <= 1;  //250 / 235 = 1
    16'b11111010_11101100 : OUT <= 1;  //250 / 236 = 1
    16'b11111010_11101101 : OUT <= 1;  //250 / 237 = 1
    16'b11111010_11101110 : OUT <= 1;  //250 / 238 = 1
    16'b11111010_11101111 : OUT <= 1;  //250 / 239 = 1
    16'b11111010_11110000 : OUT <= 1;  //250 / 240 = 1
    16'b11111010_11110001 : OUT <= 1;  //250 / 241 = 1
    16'b11111010_11110010 : OUT <= 1;  //250 / 242 = 1
    16'b11111010_11110011 : OUT <= 1;  //250 / 243 = 1
    16'b11111010_11110100 : OUT <= 1;  //250 / 244 = 1
    16'b11111010_11110101 : OUT <= 1;  //250 / 245 = 1
    16'b11111010_11110110 : OUT <= 1;  //250 / 246 = 1
    16'b11111010_11110111 : OUT <= 1;  //250 / 247 = 1
    16'b11111010_11111000 : OUT <= 1;  //250 / 248 = 1
    16'b11111010_11111001 : OUT <= 1;  //250 / 249 = 1
    16'b11111010_11111010 : OUT <= 1;  //250 / 250 = 1
    16'b11111010_11111011 : OUT <= 0;  //250 / 251 = 0
    16'b11111010_11111100 : OUT <= 0;  //250 / 252 = 0
    16'b11111010_11111101 : OUT <= 0;  //250 / 253 = 0
    16'b11111010_11111110 : OUT <= 0;  //250 / 254 = 0
    16'b11111010_11111111 : OUT <= 0;  //250 / 255 = 0
    16'b11111011_00000000 : OUT <= 0;  //251 / 0 = 0
    16'b11111011_00000001 : OUT <= 251;  //251 / 1 = 251
    16'b11111011_00000010 : OUT <= 125;  //251 / 2 = 125
    16'b11111011_00000011 : OUT <= 83;  //251 / 3 = 83
    16'b11111011_00000100 : OUT <= 62;  //251 / 4 = 62
    16'b11111011_00000101 : OUT <= 50;  //251 / 5 = 50
    16'b11111011_00000110 : OUT <= 41;  //251 / 6 = 41
    16'b11111011_00000111 : OUT <= 35;  //251 / 7 = 35
    16'b11111011_00001000 : OUT <= 31;  //251 / 8 = 31
    16'b11111011_00001001 : OUT <= 27;  //251 / 9 = 27
    16'b11111011_00001010 : OUT <= 25;  //251 / 10 = 25
    16'b11111011_00001011 : OUT <= 22;  //251 / 11 = 22
    16'b11111011_00001100 : OUT <= 20;  //251 / 12 = 20
    16'b11111011_00001101 : OUT <= 19;  //251 / 13 = 19
    16'b11111011_00001110 : OUT <= 17;  //251 / 14 = 17
    16'b11111011_00001111 : OUT <= 16;  //251 / 15 = 16
    16'b11111011_00010000 : OUT <= 15;  //251 / 16 = 15
    16'b11111011_00010001 : OUT <= 14;  //251 / 17 = 14
    16'b11111011_00010010 : OUT <= 13;  //251 / 18 = 13
    16'b11111011_00010011 : OUT <= 13;  //251 / 19 = 13
    16'b11111011_00010100 : OUT <= 12;  //251 / 20 = 12
    16'b11111011_00010101 : OUT <= 11;  //251 / 21 = 11
    16'b11111011_00010110 : OUT <= 11;  //251 / 22 = 11
    16'b11111011_00010111 : OUT <= 10;  //251 / 23 = 10
    16'b11111011_00011000 : OUT <= 10;  //251 / 24 = 10
    16'b11111011_00011001 : OUT <= 10;  //251 / 25 = 10
    16'b11111011_00011010 : OUT <= 9;  //251 / 26 = 9
    16'b11111011_00011011 : OUT <= 9;  //251 / 27 = 9
    16'b11111011_00011100 : OUT <= 8;  //251 / 28 = 8
    16'b11111011_00011101 : OUT <= 8;  //251 / 29 = 8
    16'b11111011_00011110 : OUT <= 8;  //251 / 30 = 8
    16'b11111011_00011111 : OUT <= 8;  //251 / 31 = 8
    16'b11111011_00100000 : OUT <= 7;  //251 / 32 = 7
    16'b11111011_00100001 : OUT <= 7;  //251 / 33 = 7
    16'b11111011_00100010 : OUT <= 7;  //251 / 34 = 7
    16'b11111011_00100011 : OUT <= 7;  //251 / 35 = 7
    16'b11111011_00100100 : OUT <= 6;  //251 / 36 = 6
    16'b11111011_00100101 : OUT <= 6;  //251 / 37 = 6
    16'b11111011_00100110 : OUT <= 6;  //251 / 38 = 6
    16'b11111011_00100111 : OUT <= 6;  //251 / 39 = 6
    16'b11111011_00101000 : OUT <= 6;  //251 / 40 = 6
    16'b11111011_00101001 : OUT <= 6;  //251 / 41 = 6
    16'b11111011_00101010 : OUT <= 5;  //251 / 42 = 5
    16'b11111011_00101011 : OUT <= 5;  //251 / 43 = 5
    16'b11111011_00101100 : OUT <= 5;  //251 / 44 = 5
    16'b11111011_00101101 : OUT <= 5;  //251 / 45 = 5
    16'b11111011_00101110 : OUT <= 5;  //251 / 46 = 5
    16'b11111011_00101111 : OUT <= 5;  //251 / 47 = 5
    16'b11111011_00110000 : OUT <= 5;  //251 / 48 = 5
    16'b11111011_00110001 : OUT <= 5;  //251 / 49 = 5
    16'b11111011_00110010 : OUT <= 5;  //251 / 50 = 5
    16'b11111011_00110011 : OUT <= 4;  //251 / 51 = 4
    16'b11111011_00110100 : OUT <= 4;  //251 / 52 = 4
    16'b11111011_00110101 : OUT <= 4;  //251 / 53 = 4
    16'b11111011_00110110 : OUT <= 4;  //251 / 54 = 4
    16'b11111011_00110111 : OUT <= 4;  //251 / 55 = 4
    16'b11111011_00111000 : OUT <= 4;  //251 / 56 = 4
    16'b11111011_00111001 : OUT <= 4;  //251 / 57 = 4
    16'b11111011_00111010 : OUT <= 4;  //251 / 58 = 4
    16'b11111011_00111011 : OUT <= 4;  //251 / 59 = 4
    16'b11111011_00111100 : OUT <= 4;  //251 / 60 = 4
    16'b11111011_00111101 : OUT <= 4;  //251 / 61 = 4
    16'b11111011_00111110 : OUT <= 4;  //251 / 62 = 4
    16'b11111011_00111111 : OUT <= 3;  //251 / 63 = 3
    16'b11111011_01000000 : OUT <= 3;  //251 / 64 = 3
    16'b11111011_01000001 : OUT <= 3;  //251 / 65 = 3
    16'b11111011_01000010 : OUT <= 3;  //251 / 66 = 3
    16'b11111011_01000011 : OUT <= 3;  //251 / 67 = 3
    16'b11111011_01000100 : OUT <= 3;  //251 / 68 = 3
    16'b11111011_01000101 : OUT <= 3;  //251 / 69 = 3
    16'b11111011_01000110 : OUT <= 3;  //251 / 70 = 3
    16'b11111011_01000111 : OUT <= 3;  //251 / 71 = 3
    16'b11111011_01001000 : OUT <= 3;  //251 / 72 = 3
    16'b11111011_01001001 : OUT <= 3;  //251 / 73 = 3
    16'b11111011_01001010 : OUT <= 3;  //251 / 74 = 3
    16'b11111011_01001011 : OUT <= 3;  //251 / 75 = 3
    16'b11111011_01001100 : OUT <= 3;  //251 / 76 = 3
    16'b11111011_01001101 : OUT <= 3;  //251 / 77 = 3
    16'b11111011_01001110 : OUT <= 3;  //251 / 78 = 3
    16'b11111011_01001111 : OUT <= 3;  //251 / 79 = 3
    16'b11111011_01010000 : OUT <= 3;  //251 / 80 = 3
    16'b11111011_01010001 : OUT <= 3;  //251 / 81 = 3
    16'b11111011_01010010 : OUT <= 3;  //251 / 82 = 3
    16'b11111011_01010011 : OUT <= 3;  //251 / 83 = 3
    16'b11111011_01010100 : OUT <= 2;  //251 / 84 = 2
    16'b11111011_01010101 : OUT <= 2;  //251 / 85 = 2
    16'b11111011_01010110 : OUT <= 2;  //251 / 86 = 2
    16'b11111011_01010111 : OUT <= 2;  //251 / 87 = 2
    16'b11111011_01011000 : OUT <= 2;  //251 / 88 = 2
    16'b11111011_01011001 : OUT <= 2;  //251 / 89 = 2
    16'b11111011_01011010 : OUT <= 2;  //251 / 90 = 2
    16'b11111011_01011011 : OUT <= 2;  //251 / 91 = 2
    16'b11111011_01011100 : OUT <= 2;  //251 / 92 = 2
    16'b11111011_01011101 : OUT <= 2;  //251 / 93 = 2
    16'b11111011_01011110 : OUT <= 2;  //251 / 94 = 2
    16'b11111011_01011111 : OUT <= 2;  //251 / 95 = 2
    16'b11111011_01100000 : OUT <= 2;  //251 / 96 = 2
    16'b11111011_01100001 : OUT <= 2;  //251 / 97 = 2
    16'b11111011_01100010 : OUT <= 2;  //251 / 98 = 2
    16'b11111011_01100011 : OUT <= 2;  //251 / 99 = 2
    16'b11111011_01100100 : OUT <= 2;  //251 / 100 = 2
    16'b11111011_01100101 : OUT <= 2;  //251 / 101 = 2
    16'b11111011_01100110 : OUT <= 2;  //251 / 102 = 2
    16'b11111011_01100111 : OUT <= 2;  //251 / 103 = 2
    16'b11111011_01101000 : OUT <= 2;  //251 / 104 = 2
    16'b11111011_01101001 : OUT <= 2;  //251 / 105 = 2
    16'b11111011_01101010 : OUT <= 2;  //251 / 106 = 2
    16'b11111011_01101011 : OUT <= 2;  //251 / 107 = 2
    16'b11111011_01101100 : OUT <= 2;  //251 / 108 = 2
    16'b11111011_01101101 : OUT <= 2;  //251 / 109 = 2
    16'b11111011_01101110 : OUT <= 2;  //251 / 110 = 2
    16'b11111011_01101111 : OUT <= 2;  //251 / 111 = 2
    16'b11111011_01110000 : OUT <= 2;  //251 / 112 = 2
    16'b11111011_01110001 : OUT <= 2;  //251 / 113 = 2
    16'b11111011_01110010 : OUT <= 2;  //251 / 114 = 2
    16'b11111011_01110011 : OUT <= 2;  //251 / 115 = 2
    16'b11111011_01110100 : OUT <= 2;  //251 / 116 = 2
    16'b11111011_01110101 : OUT <= 2;  //251 / 117 = 2
    16'b11111011_01110110 : OUT <= 2;  //251 / 118 = 2
    16'b11111011_01110111 : OUT <= 2;  //251 / 119 = 2
    16'b11111011_01111000 : OUT <= 2;  //251 / 120 = 2
    16'b11111011_01111001 : OUT <= 2;  //251 / 121 = 2
    16'b11111011_01111010 : OUT <= 2;  //251 / 122 = 2
    16'b11111011_01111011 : OUT <= 2;  //251 / 123 = 2
    16'b11111011_01111100 : OUT <= 2;  //251 / 124 = 2
    16'b11111011_01111101 : OUT <= 2;  //251 / 125 = 2
    16'b11111011_01111110 : OUT <= 1;  //251 / 126 = 1
    16'b11111011_01111111 : OUT <= 1;  //251 / 127 = 1
    16'b11111011_10000000 : OUT <= 1;  //251 / 128 = 1
    16'b11111011_10000001 : OUT <= 1;  //251 / 129 = 1
    16'b11111011_10000010 : OUT <= 1;  //251 / 130 = 1
    16'b11111011_10000011 : OUT <= 1;  //251 / 131 = 1
    16'b11111011_10000100 : OUT <= 1;  //251 / 132 = 1
    16'b11111011_10000101 : OUT <= 1;  //251 / 133 = 1
    16'b11111011_10000110 : OUT <= 1;  //251 / 134 = 1
    16'b11111011_10000111 : OUT <= 1;  //251 / 135 = 1
    16'b11111011_10001000 : OUT <= 1;  //251 / 136 = 1
    16'b11111011_10001001 : OUT <= 1;  //251 / 137 = 1
    16'b11111011_10001010 : OUT <= 1;  //251 / 138 = 1
    16'b11111011_10001011 : OUT <= 1;  //251 / 139 = 1
    16'b11111011_10001100 : OUT <= 1;  //251 / 140 = 1
    16'b11111011_10001101 : OUT <= 1;  //251 / 141 = 1
    16'b11111011_10001110 : OUT <= 1;  //251 / 142 = 1
    16'b11111011_10001111 : OUT <= 1;  //251 / 143 = 1
    16'b11111011_10010000 : OUT <= 1;  //251 / 144 = 1
    16'b11111011_10010001 : OUT <= 1;  //251 / 145 = 1
    16'b11111011_10010010 : OUT <= 1;  //251 / 146 = 1
    16'b11111011_10010011 : OUT <= 1;  //251 / 147 = 1
    16'b11111011_10010100 : OUT <= 1;  //251 / 148 = 1
    16'b11111011_10010101 : OUT <= 1;  //251 / 149 = 1
    16'b11111011_10010110 : OUT <= 1;  //251 / 150 = 1
    16'b11111011_10010111 : OUT <= 1;  //251 / 151 = 1
    16'b11111011_10011000 : OUT <= 1;  //251 / 152 = 1
    16'b11111011_10011001 : OUT <= 1;  //251 / 153 = 1
    16'b11111011_10011010 : OUT <= 1;  //251 / 154 = 1
    16'b11111011_10011011 : OUT <= 1;  //251 / 155 = 1
    16'b11111011_10011100 : OUT <= 1;  //251 / 156 = 1
    16'b11111011_10011101 : OUT <= 1;  //251 / 157 = 1
    16'b11111011_10011110 : OUT <= 1;  //251 / 158 = 1
    16'b11111011_10011111 : OUT <= 1;  //251 / 159 = 1
    16'b11111011_10100000 : OUT <= 1;  //251 / 160 = 1
    16'b11111011_10100001 : OUT <= 1;  //251 / 161 = 1
    16'b11111011_10100010 : OUT <= 1;  //251 / 162 = 1
    16'b11111011_10100011 : OUT <= 1;  //251 / 163 = 1
    16'b11111011_10100100 : OUT <= 1;  //251 / 164 = 1
    16'b11111011_10100101 : OUT <= 1;  //251 / 165 = 1
    16'b11111011_10100110 : OUT <= 1;  //251 / 166 = 1
    16'b11111011_10100111 : OUT <= 1;  //251 / 167 = 1
    16'b11111011_10101000 : OUT <= 1;  //251 / 168 = 1
    16'b11111011_10101001 : OUT <= 1;  //251 / 169 = 1
    16'b11111011_10101010 : OUT <= 1;  //251 / 170 = 1
    16'b11111011_10101011 : OUT <= 1;  //251 / 171 = 1
    16'b11111011_10101100 : OUT <= 1;  //251 / 172 = 1
    16'b11111011_10101101 : OUT <= 1;  //251 / 173 = 1
    16'b11111011_10101110 : OUT <= 1;  //251 / 174 = 1
    16'b11111011_10101111 : OUT <= 1;  //251 / 175 = 1
    16'b11111011_10110000 : OUT <= 1;  //251 / 176 = 1
    16'b11111011_10110001 : OUT <= 1;  //251 / 177 = 1
    16'b11111011_10110010 : OUT <= 1;  //251 / 178 = 1
    16'b11111011_10110011 : OUT <= 1;  //251 / 179 = 1
    16'b11111011_10110100 : OUT <= 1;  //251 / 180 = 1
    16'b11111011_10110101 : OUT <= 1;  //251 / 181 = 1
    16'b11111011_10110110 : OUT <= 1;  //251 / 182 = 1
    16'b11111011_10110111 : OUT <= 1;  //251 / 183 = 1
    16'b11111011_10111000 : OUT <= 1;  //251 / 184 = 1
    16'b11111011_10111001 : OUT <= 1;  //251 / 185 = 1
    16'b11111011_10111010 : OUT <= 1;  //251 / 186 = 1
    16'b11111011_10111011 : OUT <= 1;  //251 / 187 = 1
    16'b11111011_10111100 : OUT <= 1;  //251 / 188 = 1
    16'b11111011_10111101 : OUT <= 1;  //251 / 189 = 1
    16'b11111011_10111110 : OUT <= 1;  //251 / 190 = 1
    16'b11111011_10111111 : OUT <= 1;  //251 / 191 = 1
    16'b11111011_11000000 : OUT <= 1;  //251 / 192 = 1
    16'b11111011_11000001 : OUT <= 1;  //251 / 193 = 1
    16'b11111011_11000010 : OUT <= 1;  //251 / 194 = 1
    16'b11111011_11000011 : OUT <= 1;  //251 / 195 = 1
    16'b11111011_11000100 : OUT <= 1;  //251 / 196 = 1
    16'b11111011_11000101 : OUT <= 1;  //251 / 197 = 1
    16'b11111011_11000110 : OUT <= 1;  //251 / 198 = 1
    16'b11111011_11000111 : OUT <= 1;  //251 / 199 = 1
    16'b11111011_11001000 : OUT <= 1;  //251 / 200 = 1
    16'b11111011_11001001 : OUT <= 1;  //251 / 201 = 1
    16'b11111011_11001010 : OUT <= 1;  //251 / 202 = 1
    16'b11111011_11001011 : OUT <= 1;  //251 / 203 = 1
    16'b11111011_11001100 : OUT <= 1;  //251 / 204 = 1
    16'b11111011_11001101 : OUT <= 1;  //251 / 205 = 1
    16'b11111011_11001110 : OUT <= 1;  //251 / 206 = 1
    16'b11111011_11001111 : OUT <= 1;  //251 / 207 = 1
    16'b11111011_11010000 : OUT <= 1;  //251 / 208 = 1
    16'b11111011_11010001 : OUT <= 1;  //251 / 209 = 1
    16'b11111011_11010010 : OUT <= 1;  //251 / 210 = 1
    16'b11111011_11010011 : OUT <= 1;  //251 / 211 = 1
    16'b11111011_11010100 : OUT <= 1;  //251 / 212 = 1
    16'b11111011_11010101 : OUT <= 1;  //251 / 213 = 1
    16'b11111011_11010110 : OUT <= 1;  //251 / 214 = 1
    16'b11111011_11010111 : OUT <= 1;  //251 / 215 = 1
    16'b11111011_11011000 : OUT <= 1;  //251 / 216 = 1
    16'b11111011_11011001 : OUT <= 1;  //251 / 217 = 1
    16'b11111011_11011010 : OUT <= 1;  //251 / 218 = 1
    16'b11111011_11011011 : OUT <= 1;  //251 / 219 = 1
    16'b11111011_11011100 : OUT <= 1;  //251 / 220 = 1
    16'b11111011_11011101 : OUT <= 1;  //251 / 221 = 1
    16'b11111011_11011110 : OUT <= 1;  //251 / 222 = 1
    16'b11111011_11011111 : OUT <= 1;  //251 / 223 = 1
    16'b11111011_11100000 : OUT <= 1;  //251 / 224 = 1
    16'b11111011_11100001 : OUT <= 1;  //251 / 225 = 1
    16'b11111011_11100010 : OUT <= 1;  //251 / 226 = 1
    16'b11111011_11100011 : OUT <= 1;  //251 / 227 = 1
    16'b11111011_11100100 : OUT <= 1;  //251 / 228 = 1
    16'b11111011_11100101 : OUT <= 1;  //251 / 229 = 1
    16'b11111011_11100110 : OUT <= 1;  //251 / 230 = 1
    16'b11111011_11100111 : OUT <= 1;  //251 / 231 = 1
    16'b11111011_11101000 : OUT <= 1;  //251 / 232 = 1
    16'b11111011_11101001 : OUT <= 1;  //251 / 233 = 1
    16'b11111011_11101010 : OUT <= 1;  //251 / 234 = 1
    16'b11111011_11101011 : OUT <= 1;  //251 / 235 = 1
    16'b11111011_11101100 : OUT <= 1;  //251 / 236 = 1
    16'b11111011_11101101 : OUT <= 1;  //251 / 237 = 1
    16'b11111011_11101110 : OUT <= 1;  //251 / 238 = 1
    16'b11111011_11101111 : OUT <= 1;  //251 / 239 = 1
    16'b11111011_11110000 : OUT <= 1;  //251 / 240 = 1
    16'b11111011_11110001 : OUT <= 1;  //251 / 241 = 1
    16'b11111011_11110010 : OUT <= 1;  //251 / 242 = 1
    16'b11111011_11110011 : OUT <= 1;  //251 / 243 = 1
    16'b11111011_11110100 : OUT <= 1;  //251 / 244 = 1
    16'b11111011_11110101 : OUT <= 1;  //251 / 245 = 1
    16'b11111011_11110110 : OUT <= 1;  //251 / 246 = 1
    16'b11111011_11110111 : OUT <= 1;  //251 / 247 = 1
    16'b11111011_11111000 : OUT <= 1;  //251 / 248 = 1
    16'b11111011_11111001 : OUT <= 1;  //251 / 249 = 1
    16'b11111011_11111010 : OUT <= 1;  //251 / 250 = 1
    16'b11111011_11111011 : OUT <= 1;  //251 / 251 = 1
    16'b11111011_11111100 : OUT <= 0;  //251 / 252 = 0
    16'b11111011_11111101 : OUT <= 0;  //251 / 253 = 0
    16'b11111011_11111110 : OUT <= 0;  //251 / 254 = 0
    16'b11111011_11111111 : OUT <= 0;  //251 / 255 = 0
    16'b11111100_00000000 : OUT <= 0;  //252 / 0 = 0
    16'b11111100_00000001 : OUT <= 252;  //252 / 1 = 252
    16'b11111100_00000010 : OUT <= 126;  //252 / 2 = 126
    16'b11111100_00000011 : OUT <= 84;  //252 / 3 = 84
    16'b11111100_00000100 : OUT <= 63;  //252 / 4 = 63
    16'b11111100_00000101 : OUT <= 50;  //252 / 5 = 50
    16'b11111100_00000110 : OUT <= 42;  //252 / 6 = 42
    16'b11111100_00000111 : OUT <= 36;  //252 / 7 = 36
    16'b11111100_00001000 : OUT <= 31;  //252 / 8 = 31
    16'b11111100_00001001 : OUT <= 28;  //252 / 9 = 28
    16'b11111100_00001010 : OUT <= 25;  //252 / 10 = 25
    16'b11111100_00001011 : OUT <= 22;  //252 / 11 = 22
    16'b11111100_00001100 : OUT <= 21;  //252 / 12 = 21
    16'b11111100_00001101 : OUT <= 19;  //252 / 13 = 19
    16'b11111100_00001110 : OUT <= 18;  //252 / 14 = 18
    16'b11111100_00001111 : OUT <= 16;  //252 / 15 = 16
    16'b11111100_00010000 : OUT <= 15;  //252 / 16 = 15
    16'b11111100_00010001 : OUT <= 14;  //252 / 17 = 14
    16'b11111100_00010010 : OUT <= 14;  //252 / 18 = 14
    16'b11111100_00010011 : OUT <= 13;  //252 / 19 = 13
    16'b11111100_00010100 : OUT <= 12;  //252 / 20 = 12
    16'b11111100_00010101 : OUT <= 12;  //252 / 21 = 12
    16'b11111100_00010110 : OUT <= 11;  //252 / 22 = 11
    16'b11111100_00010111 : OUT <= 10;  //252 / 23 = 10
    16'b11111100_00011000 : OUT <= 10;  //252 / 24 = 10
    16'b11111100_00011001 : OUT <= 10;  //252 / 25 = 10
    16'b11111100_00011010 : OUT <= 9;  //252 / 26 = 9
    16'b11111100_00011011 : OUT <= 9;  //252 / 27 = 9
    16'b11111100_00011100 : OUT <= 9;  //252 / 28 = 9
    16'b11111100_00011101 : OUT <= 8;  //252 / 29 = 8
    16'b11111100_00011110 : OUT <= 8;  //252 / 30 = 8
    16'b11111100_00011111 : OUT <= 8;  //252 / 31 = 8
    16'b11111100_00100000 : OUT <= 7;  //252 / 32 = 7
    16'b11111100_00100001 : OUT <= 7;  //252 / 33 = 7
    16'b11111100_00100010 : OUT <= 7;  //252 / 34 = 7
    16'b11111100_00100011 : OUT <= 7;  //252 / 35 = 7
    16'b11111100_00100100 : OUT <= 7;  //252 / 36 = 7
    16'b11111100_00100101 : OUT <= 6;  //252 / 37 = 6
    16'b11111100_00100110 : OUT <= 6;  //252 / 38 = 6
    16'b11111100_00100111 : OUT <= 6;  //252 / 39 = 6
    16'b11111100_00101000 : OUT <= 6;  //252 / 40 = 6
    16'b11111100_00101001 : OUT <= 6;  //252 / 41 = 6
    16'b11111100_00101010 : OUT <= 6;  //252 / 42 = 6
    16'b11111100_00101011 : OUT <= 5;  //252 / 43 = 5
    16'b11111100_00101100 : OUT <= 5;  //252 / 44 = 5
    16'b11111100_00101101 : OUT <= 5;  //252 / 45 = 5
    16'b11111100_00101110 : OUT <= 5;  //252 / 46 = 5
    16'b11111100_00101111 : OUT <= 5;  //252 / 47 = 5
    16'b11111100_00110000 : OUT <= 5;  //252 / 48 = 5
    16'b11111100_00110001 : OUT <= 5;  //252 / 49 = 5
    16'b11111100_00110010 : OUT <= 5;  //252 / 50 = 5
    16'b11111100_00110011 : OUT <= 4;  //252 / 51 = 4
    16'b11111100_00110100 : OUT <= 4;  //252 / 52 = 4
    16'b11111100_00110101 : OUT <= 4;  //252 / 53 = 4
    16'b11111100_00110110 : OUT <= 4;  //252 / 54 = 4
    16'b11111100_00110111 : OUT <= 4;  //252 / 55 = 4
    16'b11111100_00111000 : OUT <= 4;  //252 / 56 = 4
    16'b11111100_00111001 : OUT <= 4;  //252 / 57 = 4
    16'b11111100_00111010 : OUT <= 4;  //252 / 58 = 4
    16'b11111100_00111011 : OUT <= 4;  //252 / 59 = 4
    16'b11111100_00111100 : OUT <= 4;  //252 / 60 = 4
    16'b11111100_00111101 : OUT <= 4;  //252 / 61 = 4
    16'b11111100_00111110 : OUT <= 4;  //252 / 62 = 4
    16'b11111100_00111111 : OUT <= 4;  //252 / 63 = 4
    16'b11111100_01000000 : OUT <= 3;  //252 / 64 = 3
    16'b11111100_01000001 : OUT <= 3;  //252 / 65 = 3
    16'b11111100_01000010 : OUT <= 3;  //252 / 66 = 3
    16'b11111100_01000011 : OUT <= 3;  //252 / 67 = 3
    16'b11111100_01000100 : OUT <= 3;  //252 / 68 = 3
    16'b11111100_01000101 : OUT <= 3;  //252 / 69 = 3
    16'b11111100_01000110 : OUT <= 3;  //252 / 70 = 3
    16'b11111100_01000111 : OUT <= 3;  //252 / 71 = 3
    16'b11111100_01001000 : OUT <= 3;  //252 / 72 = 3
    16'b11111100_01001001 : OUT <= 3;  //252 / 73 = 3
    16'b11111100_01001010 : OUT <= 3;  //252 / 74 = 3
    16'b11111100_01001011 : OUT <= 3;  //252 / 75 = 3
    16'b11111100_01001100 : OUT <= 3;  //252 / 76 = 3
    16'b11111100_01001101 : OUT <= 3;  //252 / 77 = 3
    16'b11111100_01001110 : OUT <= 3;  //252 / 78 = 3
    16'b11111100_01001111 : OUT <= 3;  //252 / 79 = 3
    16'b11111100_01010000 : OUT <= 3;  //252 / 80 = 3
    16'b11111100_01010001 : OUT <= 3;  //252 / 81 = 3
    16'b11111100_01010010 : OUT <= 3;  //252 / 82 = 3
    16'b11111100_01010011 : OUT <= 3;  //252 / 83 = 3
    16'b11111100_01010100 : OUT <= 3;  //252 / 84 = 3
    16'b11111100_01010101 : OUT <= 2;  //252 / 85 = 2
    16'b11111100_01010110 : OUT <= 2;  //252 / 86 = 2
    16'b11111100_01010111 : OUT <= 2;  //252 / 87 = 2
    16'b11111100_01011000 : OUT <= 2;  //252 / 88 = 2
    16'b11111100_01011001 : OUT <= 2;  //252 / 89 = 2
    16'b11111100_01011010 : OUT <= 2;  //252 / 90 = 2
    16'b11111100_01011011 : OUT <= 2;  //252 / 91 = 2
    16'b11111100_01011100 : OUT <= 2;  //252 / 92 = 2
    16'b11111100_01011101 : OUT <= 2;  //252 / 93 = 2
    16'b11111100_01011110 : OUT <= 2;  //252 / 94 = 2
    16'b11111100_01011111 : OUT <= 2;  //252 / 95 = 2
    16'b11111100_01100000 : OUT <= 2;  //252 / 96 = 2
    16'b11111100_01100001 : OUT <= 2;  //252 / 97 = 2
    16'b11111100_01100010 : OUT <= 2;  //252 / 98 = 2
    16'b11111100_01100011 : OUT <= 2;  //252 / 99 = 2
    16'b11111100_01100100 : OUT <= 2;  //252 / 100 = 2
    16'b11111100_01100101 : OUT <= 2;  //252 / 101 = 2
    16'b11111100_01100110 : OUT <= 2;  //252 / 102 = 2
    16'b11111100_01100111 : OUT <= 2;  //252 / 103 = 2
    16'b11111100_01101000 : OUT <= 2;  //252 / 104 = 2
    16'b11111100_01101001 : OUT <= 2;  //252 / 105 = 2
    16'b11111100_01101010 : OUT <= 2;  //252 / 106 = 2
    16'b11111100_01101011 : OUT <= 2;  //252 / 107 = 2
    16'b11111100_01101100 : OUT <= 2;  //252 / 108 = 2
    16'b11111100_01101101 : OUT <= 2;  //252 / 109 = 2
    16'b11111100_01101110 : OUT <= 2;  //252 / 110 = 2
    16'b11111100_01101111 : OUT <= 2;  //252 / 111 = 2
    16'b11111100_01110000 : OUT <= 2;  //252 / 112 = 2
    16'b11111100_01110001 : OUT <= 2;  //252 / 113 = 2
    16'b11111100_01110010 : OUT <= 2;  //252 / 114 = 2
    16'b11111100_01110011 : OUT <= 2;  //252 / 115 = 2
    16'b11111100_01110100 : OUT <= 2;  //252 / 116 = 2
    16'b11111100_01110101 : OUT <= 2;  //252 / 117 = 2
    16'b11111100_01110110 : OUT <= 2;  //252 / 118 = 2
    16'b11111100_01110111 : OUT <= 2;  //252 / 119 = 2
    16'b11111100_01111000 : OUT <= 2;  //252 / 120 = 2
    16'b11111100_01111001 : OUT <= 2;  //252 / 121 = 2
    16'b11111100_01111010 : OUT <= 2;  //252 / 122 = 2
    16'b11111100_01111011 : OUT <= 2;  //252 / 123 = 2
    16'b11111100_01111100 : OUT <= 2;  //252 / 124 = 2
    16'b11111100_01111101 : OUT <= 2;  //252 / 125 = 2
    16'b11111100_01111110 : OUT <= 2;  //252 / 126 = 2
    16'b11111100_01111111 : OUT <= 1;  //252 / 127 = 1
    16'b11111100_10000000 : OUT <= 1;  //252 / 128 = 1
    16'b11111100_10000001 : OUT <= 1;  //252 / 129 = 1
    16'b11111100_10000010 : OUT <= 1;  //252 / 130 = 1
    16'b11111100_10000011 : OUT <= 1;  //252 / 131 = 1
    16'b11111100_10000100 : OUT <= 1;  //252 / 132 = 1
    16'b11111100_10000101 : OUT <= 1;  //252 / 133 = 1
    16'b11111100_10000110 : OUT <= 1;  //252 / 134 = 1
    16'b11111100_10000111 : OUT <= 1;  //252 / 135 = 1
    16'b11111100_10001000 : OUT <= 1;  //252 / 136 = 1
    16'b11111100_10001001 : OUT <= 1;  //252 / 137 = 1
    16'b11111100_10001010 : OUT <= 1;  //252 / 138 = 1
    16'b11111100_10001011 : OUT <= 1;  //252 / 139 = 1
    16'b11111100_10001100 : OUT <= 1;  //252 / 140 = 1
    16'b11111100_10001101 : OUT <= 1;  //252 / 141 = 1
    16'b11111100_10001110 : OUT <= 1;  //252 / 142 = 1
    16'b11111100_10001111 : OUT <= 1;  //252 / 143 = 1
    16'b11111100_10010000 : OUT <= 1;  //252 / 144 = 1
    16'b11111100_10010001 : OUT <= 1;  //252 / 145 = 1
    16'b11111100_10010010 : OUT <= 1;  //252 / 146 = 1
    16'b11111100_10010011 : OUT <= 1;  //252 / 147 = 1
    16'b11111100_10010100 : OUT <= 1;  //252 / 148 = 1
    16'b11111100_10010101 : OUT <= 1;  //252 / 149 = 1
    16'b11111100_10010110 : OUT <= 1;  //252 / 150 = 1
    16'b11111100_10010111 : OUT <= 1;  //252 / 151 = 1
    16'b11111100_10011000 : OUT <= 1;  //252 / 152 = 1
    16'b11111100_10011001 : OUT <= 1;  //252 / 153 = 1
    16'b11111100_10011010 : OUT <= 1;  //252 / 154 = 1
    16'b11111100_10011011 : OUT <= 1;  //252 / 155 = 1
    16'b11111100_10011100 : OUT <= 1;  //252 / 156 = 1
    16'b11111100_10011101 : OUT <= 1;  //252 / 157 = 1
    16'b11111100_10011110 : OUT <= 1;  //252 / 158 = 1
    16'b11111100_10011111 : OUT <= 1;  //252 / 159 = 1
    16'b11111100_10100000 : OUT <= 1;  //252 / 160 = 1
    16'b11111100_10100001 : OUT <= 1;  //252 / 161 = 1
    16'b11111100_10100010 : OUT <= 1;  //252 / 162 = 1
    16'b11111100_10100011 : OUT <= 1;  //252 / 163 = 1
    16'b11111100_10100100 : OUT <= 1;  //252 / 164 = 1
    16'b11111100_10100101 : OUT <= 1;  //252 / 165 = 1
    16'b11111100_10100110 : OUT <= 1;  //252 / 166 = 1
    16'b11111100_10100111 : OUT <= 1;  //252 / 167 = 1
    16'b11111100_10101000 : OUT <= 1;  //252 / 168 = 1
    16'b11111100_10101001 : OUT <= 1;  //252 / 169 = 1
    16'b11111100_10101010 : OUT <= 1;  //252 / 170 = 1
    16'b11111100_10101011 : OUT <= 1;  //252 / 171 = 1
    16'b11111100_10101100 : OUT <= 1;  //252 / 172 = 1
    16'b11111100_10101101 : OUT <= 1;  //252 / 173 = 1
    16'b11111100_10101110 : OUT <= 1;  //252 / 174 = 1
    16'b11111100_10101111 : OUT <= 1;  //252 / 175 = 1
    16'b11111100_10110000 : OUT <= 1;  //252 / 176 = 1
    16'b11111100_10110001 : OUT <= 1;  //252 / 177 = 1
    16'b11111100_10110010 : OUT <= 1;  //252 / 178 = 1
    16'b11111100_10110011 : OUT <= 1;  //252 / 179 = 1
    16'b11111100_10110100 : OUT <= 1;  //252 / 180 = 1
    16'b11111100_10110101 : OUT <= 1;  //252 / 181 = 1
    16'b11111100_10110110 : OUT <= 1;  //252 / 182 = 1
    16'b11111100_10110111 : OUT <= 1;  //252 / 183 = 1
    16'b11111100_10111000 : OUT <= 1;  //252 / 184 = 1
    16'b11111100_10111001 : OUT <= 1;  //252 / 185 = 1
    16'b11111100_10111010 : OUT <= 1;  //252 / 186 = 1
    16'b11111100_10111011 : OUT <= 1;  //252 / 187 = 1
    16'b11111100_10111100 : OUT <= 1;  //252 / 188 = 1
    16'b11111100_10111101 : OUT <= 1;  //252 / 189 = 1
    16'b11111100_10111110 : OUT <= 1;  //252 / 190 = 1
    16'b11111100_10111111 : OUT <= 1;  //252 / 191 = 1
    16'b11111100_11000000 : OUT <= 1;  //252 / 192 = 1
    16'b11111100_11000001 : OUT <= 1;  //252 / 193 = 1
    16'b11111100_11000010 : OUT <= 1;  //252 / 194 = 1
    16'b11111100_11000011 : OUT <= 1;  //252 / 195 = 1
    16'b11111100_11000100 : OUT <= 1;  //252 / 196 = 1
    16'b11111100_11000101 : OUT <= 1;  //252 / 197 = 1
    16'b11111100_11000110 : OUT <= 1;  //252 / 198 = 1
    16'b11111100_11000111 : OUT <= 1;  //252 / 199 = 1
    16'b11111100_11001000 : OUT <= 1;  //252 / 200 = 1
    16'b11111100_11001001 : OUT <= 1;  //252 / 201 = 1
    16'b11111100_11001010 : OUT <= 1;  //252 / 202 = 1
    16'b11111100_11001011 : OUT <= 1;  //252 / 203 = 1
    16'b11111100_11001100 : OUT <= 1;  //252 / 204 = 1
    16'b11111100_11001101 : OUT <= 1;  //252 / 205 = 1
    16'b11111100_11001110 : OUT <= 1;  //252 / 206 = 1
    16'b11111100_11001111 : OUT <= 1;  //252 / 207 = 1
    16'b11111100_11010000 : OUT <= 1;  //252 / 208 = 1
    16'b11111100_11010001 : OUT <= 1;  //252 / 209 = 1
    16'b11111100_11010010 : OUT <= 1;  //252 / 210 = 1
    16'b11111100_11010011 : OUT <= 1;  //252 / 211 = 1
    16'b11111100_11010100 : OUT <= 1;  //252 / 212 = 1
    16'b11111100_11010101 : OUT <= 1;  //252 / 213 = 1
    16'b11111100_11010110 : OUT <= 1;  //252 / 214 = 1
    16'b11111100_11010111 : OUT <= 1;  //252 / 215 = 1
    16'b11111100_11011000 : OUT <= 1;  //252 / 216 = 1
    16'b11111100_11011001 : OUT <= 1;  //252 / 217 = 1
    16'b11111100_11011010 : OUT <= 1;  //252 / 218 = 1
    16'b11111100_11011011 : OUT <= 1;  //252 / 219 = 1
    16'b11111100_11011100 : OUT <= 1;  //252 / 220 = 1
    16'b11111100_11011101 : OUT <= 1;  //252 / 221 = 1
    16'b11111100_11011110 : OUT <= 1;  //252 / 222 = 1
    16'b11111100_11011111 : OUT <= 1;  //252 / 223 = 1
    16'b11111100_11100000 : OUT <= 1;  //252 / 224 = 1
    16'b11111100_11100001 : OUT <= 1;  //252 / 225 = 1
    16'b11111100_11100010 : OUT <= 1;  //252 / 226 = 1
    16'b11111100_11100011 : OUT <= 1;  //252 / 227 = 1
    16'b11111100_11100100 : OUT <= 1;  //252 / 228 = 1
    16'b11111100_11100101 : OUT <= 1;  //252 / 229 = 1
    16'b11111100_11100110 : OUT <= 1;  //252 / 230 = 1
    16'b11111100_11100111 : OUT <= 1;  //252 / 231 = 1
    16'b11111100_11101000 : OUT <= 1;  //252 / 232 = 1
    16'b11111100_11101001 : OUT <= 1;  //252 / 233 = 1
    16'b11111100_11101010 : OUT <= 1;  //252 / 234 = 1
    16'b11111100_11101011 : OUT <= 1;  //252 / 235 = 1
    16'b11111100_11101100 : OUT <= 1;  //252 / 236 = 1
    16'b11111100_11101101 : OUT <= 1;  //252 / 237 = 1
    16'b11111100_11101110 : OUT <= 1;  //252 / 238 = 1
    16'b11111100_11101111 : OUT <= 1;  //252 / 239 = 1
    16'b11111100_11110000 : OUT <= 1;  //252 / 240 = 1
    16'b11111100_11110001 : OUT <= 1;  //252 / 241 = 1
    16'b11111100_11110010 : OUT <= 1;  //252 / 242 = 1
    16'b11111100_11110011 : OUT <= 1;  //252 / 243 = 1
    16'b11111100_11110100 : OUT <= 1;  //252 / 244 = 1
    16'b11111100_11110101 : OUT <= 1;  //252 / 245 = 1
    16'b11111100_11110110 : OUT <= 1;  //252 / 246 = 1
    16'b11111100_11110111 : OUT <= 1;  //252 / 247 = 1
    16'b11111100_11111000 : OUT <= 1;  //252 / 248 = 1
    16'b11111100_11111001 : OUT <= 1;  //252 / 249 = 1
    16'b11111100_11111010 : OUT <= 1;  //252 / 250 = 1
    16'b11111100_11111011 : OUT <= 1;  //252 / 251 = 1
    16'b11111100_11111100 : OUT <= 1;  //252 / 252 = 1
    16'b11111100_11111101 : OUT <= 0;  //252 / 253 = 0
    16'b11111100_11111110 : OUT <= 0;  //252 / 254 = 0
    16'b11111100_11111111 : OUT <= 0;  //252 / 255 = 0
    16'b11111101_00000000 : OUT <= 0;  //253 / 0 = 0
    16'b11111101_00000001 : OUT <= 253;  //253 / 1 = 253
    16'b11111101_00000010 : OUT <= 126;  //253 / 2 = 126
    16'b11111101_00000011 : OUT <= 84;  //253 / 3 = 84
    16'b11111101_00000100 : OUT <= 63;  //253 / 4 = 63
    16'b11111101_00000101 : OUT <= 50;  //253 / 5 = 50
    16'b11111101_00000110 : OUT <= 42;  //253 / 6 = 42
    16'b11111101_00000111 : OUT <= 36;  //253 / 7 = 36
    16'b11111101_00001000 : OUT <= 31;  //253 / 8 = 31
    16'b11111101_00001001 : OUT <= 28;  //253 / 9 = 28
    16'b11111101_00001010 : OUT <= 25;  //253 / 10 = 25
    16'b11111101_00001011 : OUT <= 23;  //253 / 11 = 23
    16'b11111101_00001100 : OUT <= 21;  //253 / 12 = 21
    16'b11111101_00001101 : OUT <= 19;  //253 / 13 = 19
    16'b11111101_00001110 : OUT <= 18;  //253 / 14 = 18
    16'b11111101_00001111 : OUT <= 16;  //253 / 15 = 16
    16'b11111101_00010000 : OUT <= 15;  //253 / 16 = 15
    16'b11111101_00010001 : OUT <= 14;  //253 / 17 = 14
    16'b11111101_00010010 : OUT <= 14;  //253 / 18 = 14
    16'b11111101_00010011 : OUT <= 13;  //253 / 19 = 13
    16'b11111101_00010100 : OUT <= 12;  //253 / 20 = 12
    16'b11111101_00010101 : OUT <= 12;  //253 / 21 = 12
    16'b11111101_00010110 : OUT <= 11;  //253 / 22 = 11
    16'b11111101_00010111 : OUT <= 11;  //253 / 23 = 11
    16'b11111101_00011000 : OUT <= 10;  //253 / 24 = 10
    16'b11111101_00011001 : OUT <= 10;  //253 / 25 = 10
    16'b11111101_00011010 : OUT <= 9;  //253 / 26 = 9
    16'b11111101_00011011 : OUT <= 9;  //253 / 27 = 9
    16'b11111101_00011100 : OUT <= 9;  //253 / 28 = 9
    16'b11111101_00011101 : OUT <= 8;  //253 / 29 = 8
    16'b11111101_00011110 : OUT <= 8;  //253 / 30 = 8
    16'b11111101_00011111 : OUT <= 8;  //253 / 31 = 8
    16'b11111101_00100000 : OUT <= 7;  //253 / 32 = 7
    16'b11111101_00100001 : OUT <= 7;  //253 / 33 = 7
    16'b11111101_00100010 : OUT <= 7;  //253 / 34 = 7
    16'b11111101_00100011 : OUT <= 7;  //253 / 35 = 7
    16'b11111101_00100100 : OUT <= 7;  //253 / 36 = 7
    16'b11111101_00100101 : OUT <= 6;  //253 / 37 = 6
    16'b11111101_00100110 : OUT <= 6;  //253 / 38 = 6
    16'b11111101_00100111 : OUT <= 6;  //253 / 39 = 6
    16'b11111101_00101000 : OUT <= 6;  //253 / 40 = 6
    16'b11111101_00101001 : OUT <= 6;  //253 / 41 = 6
    16'b11111101_00101010 : OUT <= 6;  //253 / 42 = 6
    16'b11111101_00101011 : OUT <= 5;  //253 / 43 = 5
    16'b11111101_00101100 : OUT <= 5;  //253 / 44 = 5
    16'b11111101_00101101 : OUT <= 5;  //253 / 45 = 5
    16'b11111101_00101110 : OUT <= 5;  //253 / 46 = 5
    16'b11111101_00101111 : OUT <= 5;  //253 / 47 = 5
    16'b11111101_00110000 : OUT <= 5;  //253 / 48 = 5
    16'b11111101_00110001 : OUT <= 5;  //253 / 49 = 5
    16'b11111101_00110010 : OUT <= 5;  //253 / 50 = 5
    16'b11111101_00110011 : OUT <= 4;  //253 / 51 = 4
    16'b11111101_00110100 : OUT <= 4;  //253 / 52 = 4
    16'b11111101_00110101 : OUT <= 4;  //253 / 53 = 4
    16'b11111101_00110110 : OUT <= 4;  //253 / 54 = 4
    16'b11111101_00110111 : OUT <= 4;  //253 / 55 = 4
    16'b11111101_00111000 : OUT <= 4;  //253 / 56 = 4
    16'b11111101_00111001 : OUT <= 4;  //253 / 57 = 4
    16'b11111101_00111010 : OUT <= 4;  //253 / 58 = 4
    16'b11111101_00111011 : OUT <= 4;  //253 / 59 = 4
    16'b11111101_00111100 : OUT <= 4;  //253 / 60 = 4
    16'b11111101_00111101 : OUT <= 4;  //253 / 61 = 4
    16'b11111101_00111110 : OUT <= 4;  //253 / 62 = 4
    16'b11111101_00111111 : OUT <= 4;  //253 / 63 = 4
    16'b11111101_01000000 : OUT <= 3;  //253 / 64 = 3
    16'b11111101_01000001 : OUT <= 3;  //253 / 65 = 3
    16'b11111101_01000010 : OUT <= 3;  //253 / 66 = 3
    16'b11111101_01000011 : OUT <= 3;  //253 / 67 = 3
    16'b11111101_01000100 : OUT <= 3;  //253 / 68 = 3
    16'b11111101_01000101 : OUT <= 3;  //253 / 69 = 3
    16'b11111101_01000110 : OUT <= 3;  //253 / 70 = 3
    16'b11111101_01000111 : OUT <= 3;  //253 / 71 = 3
    16'b11111101_01001000 : OUT <= 3;  //253 / 72 = 3
    16'b11111101_01001001 : OUT <= 3;  //253 / 73 = 3
    16'b11111101_01001010 : OUT <= 3;  //253 / 74 = 3
    16'b11111101_01001011 : OUT <= 3;  //253 / 75 = 3
    16'b11111101_01001100 : OUT <= 3;  //253 / 76 = 3
    16'b11111101_01001101 : OUT <= 3;  //253 / 77 = 3
    16'b11111101_01001110 : OUT <= 3;  //253 / 78 = 3
    16'b11111101_01001111 : OUT <= 3;  //253 / 79 = 3
    16'b11111101_01010000 : OUT <= 3;  //253 / 80 = 3
    16'b11111101_01010001 : OUT <= 3;  //253 / 81 = 3
    16'b11111101_01010010 : OUT <= 3;  //253 / 82 = 3
    16'b11111101_01010011 : OUT <= 3;  //253 / 83 = 3
    16'b11111101_01010100 : OUT <= 3;  //253 / 84 = 3
    16'b11111101_01010101 : OUT <= 2;  //253 / 85 = 2
    16'b11111101_01010110 : OUT <= 2;  //253 / 86 = 2
    16'b11111101_01010111 : OUT <= 2;  //253 / 87 = 2
    16'b11111101_01011000 : OUT <= 2;  //253 / 88 = 2
    16'b11111101_01011001 : OUT <= 2;  //253 / 89 = 2
    16'b11111101_01011010 : OUT <= 2;  //253 / 90 = 2
    16'b11111101_01011011 : OUT <= 2;  //253 / 91 = 2
    16'b11111101_01011100 : OUT <= 2;  //253 / 92 = 2
    16'b11111101_01011101 : OUT <= 2;  //253 / 93 = 2
    16'b11111101_01011110 : OUT <= 2;  //253 / 94 = 2
    16'b11111101_01011111 : OUT <= 2;  //253 / 95 = 2
    16'b11111101_01100000 : OUT <= 2;  //253 / 96 = 2
    16'b11111101_01100001 : OUT <= 2;  //253 / 97 = 2
    16'b11111101_01100010 : OUT <= 2;  //253 / 98 = 2
    16'b11111101_01100011 : OUT <= 2;  //253 / 99 = 2
    16'b11111101_01100100 : OUT <= 2;  //253 / 100 = 2
    16'b11111101_01100101 : OUT <= 2;  //253 / 101 = 2
    16'b11111101_01100110 : OUT <= 2;  //253 / 102 = 2
    16'b11111101_01100111 : OUT <= 2;  //253 / 103 = 2
    16'b11111101_01101000 : OUT <= 2;  //253 / 104 = 2
    16'b11111101_01101001 : OUT <= 2;  //253 / 105 = 2
    16'b11111101_01101010 : OUT <= 2;  //253 / 106 = 2
    16'b11111101_01101011 : OUT <= 2;  //253 / 107 = 2
    16'b11111101_01101100 : OUT <= 2;  //253 / 108 = 2
    16'b11111101_01101101 : OUT <= 2;  //253 / 109 = 2
    16'b11111101_01101110 : OUT <= 2;  //253 / 110 = 2
    16'b11111101_01101111 : OUT <= 2;  //253 / 111 = 2
    16'b11111101_01110000 : OUT <= 2;  //253 / 112 = 2
    16'b11111101_01110001 : OUT <= 2;  //253 / 113 = 2
    16'b11111101_01110010 : OUT <= 2;  //253 / 114 = 2
    16'b11111101_01110011 : OUT <= 2;  //253 / 115 = 2
    16'b11111101_01110100 : OUT <= 2;  //253 / 116 = 2
    16'b11111101_01110101 : OUT <= 2;  //253 / 117 = 2
    16'b11111101_01110110 : OUT <= 2;  //253 / 118 = 2
    16'b11111101_01110111 : OUT <= 2;  //253 / 119 = 2
    16'b11111101_01111000 : OUT <= 2;  //253 / 120 = 2
    16'b11111101_01111001 : OUT <= 2;  //253 / 121 = 2
    16'b11111101_01111010 : OUT <= 2;  //253 / 122 = 2
    16'b11111101_01111011 : OUT <= 2;  //253 / 123 = 2
    16'b11111101_01111100 : OUT <= 2;  //253 / 124 = 2
    16'b11111101_01111101 : OUT <= 2;  //253 / 125 = 2
    16'b11111101_01111110 : OUT <= 2;  //253 / 126 = 2
    16'b11111101_01111111 : OUT <= 1;  //253 / 127 = 1
    16'b11111101_10000000 : OUT <= 1;  //253 / 128 = 1
    16'b11111101_10000001 : OUT <= 1;  //253 / 129 = 1
    16'b11111101_10000010 : OUT <= 1;  //253 / 130 = 1
    16'b11111101_10000011 : OUT <= 1;  //253 / 131 = 1
    16'b11111101_10000100 : OUT <= 1;  //253 / 132 = 1
    16'b11111101_10000101 : OUT <= 1;  //253 / 133 = 1
    16'b11111101_10000110 : OUT <= 1;  //253 / 134 = 1
    16'b11111101_10000111 : OUT <= 1;  //253 / 135 = 1
    16'b11111101_10001000 : OUT <= 1;  //253 / 136 = 1
    16'b11111101_10001001 : OUT <= 1;  //253 / 137 = 1
    16'b11111101_10001010 : OUT <= 1;  //253 / 138 = 1
    16'b11111101_10001011 : OUT <= 1;  //253 / 139 = 1
    16'b11111101_10001100 : OUT <= 1;  //253 / 140 = 1
    16'b11111101_10001101 : OUT <= 1;  //253 / 141 = 1
    16'b11111101_10001110 : OUT <= 1;  //253 / 142 = 1
    16'b11111101_10001111 : OUT <= 1;  //253 / 143 = 1
    16'b11111101_10010000 : OUT <= 1;  //253 / 144 = 1
    16'b11111101_10010001 : OUT <= 1;  //253 / 145 = 1
    16'b11111101_10010010 : OUT <= 1;  //253 / 146 = 1
    16'b11111101_10010011 : OUT <= 1;  //253 / 147 = 1
    16'b11111101_10010100 : OUT <= 1;  //253 / 148 = 1
    16'b11111101_10010101 : OUT <= 1;  //253 / 149 = 1
    16'b11111101_10010110 : OUT <= 1;  //253 / 150 = 1
    16'b11111101_10010111 : OUT <= 1;  //253 / 151 = 1
    16'b11111101_10011000 : OUT <= 1;  //253 / 152 = 1
    16'b11111101_10011001 : OUT <= 1;  //253 / 153 = 1
    16'b11111101_10011010 : OUT <= 1;  //253 / 154 = 1
    16'b11111101_10011011 : OUT <= 1;  //253 / 155 = 1
    16'b11111101_10011100 : OUT <= 1;  //253 / 156 = 1
    16'b11111101_10011101 : OUT <= 1;  //253 / 157 = 1
    16'b11111101_10011110 : OUT <= 1;  //253 / 158 = 1
    16'b11111101_10011111 : OUT <= 1;  //253 / 159 = 1
    16'b11111101_10100000 : OUT <= 1;  //253 / 160 = 1
    16'b11111101_10100001 : OUT <= 1;  //253 / 161 = 1
    16'b11111101_10100010 : OUT <= 1;  //253 / 162 = 1
    16'b11111101_10100011 : OUT <= 1;  //253 / 163 = 1
    16'b11111101_10100100 : OUT <= 1;  //253 / 164 = 1
    16'b11111101_10100101 : OUT <= 1;  //253 / 165 = 1
    16'b11111101_10100110 : OUT <= 1;  //253 / 166 = 1
    16'b11111101_10100111 : OUT <= 1;  //253 / 167 = 1
    16'b11111101_10101000 : OUT <= 1;  //253 / 168 = 1
    16'b11111101_10101001 : OUT <= 1;  //253 / 169 = 1
    16'b11111101_10101010 : OUT <= 1;  //253 / 170 = 1
    16'b11111101_10101011 : OUT <= 1;  //253 / 171 = 1
    16'b11111101_10101100 : OUT <= 1;  //253 / 172 = 1
    16'b11111101_10101101 : OUT <= 1;  //253 / 173 = 1
    16'b11111101_10101110 : OUT <= 1;  //253 / 174 = 1
    16'b11111101_10101111 : OUT <= 1;  //253 / 175 = 1
    16'b11111101_10110000 : OUT <= 1;  //253 / 176 = 1
    16'b11111101_10110001 : OUT <= 1;  //253 / 177 = 1
    16'b11111101_10110010 : OUT <= 1;  //253 / 178 = 1
    16'b11111101_10110011 : OUT <= 1;  //253 / 179 = 1
    16'b11111101_10110100 : OUT <= 1;  //253 / 180 = 1
    16'b11111101_10110101 : OUT <= 1;  //253 / 181 = 1
    16'b11111101_10110110 : OUT <= 1;  //253 / 182 = 1
    16'b11111101_10110111 : OUT <= 1;  //253 / 183 = 1
    16'b11111101_10111000 : OUT <= 1;  //253 / 184 = 1
    16'b11111101_10111001 : OUT <= 1;  //253 / 185 = 1
    16'b11111101_10111010 : OUT <= 1;  //253 / 186 = 1
    16'b11111101_10111011 : OUT <= 1;  //253 / 187 = 1
    16'b11111101_10111100 : OUT <= 1;  //253 / 188 = 1
    16'b11111101_10111101 : OUT <= 1;  //253 / 189 = 1
    16'b11111101_10111110 : OUT <= 1;  //253 / 190 = 1
    16'b11111101_10111111 : OUT <= 1;  //253 / 191 = 1
    16'b11111101_11000000 : OUT <= 1;  //253 / 192 = 1
    16'b11111101_11000001 : OUT <= 1;  //253 / 193 = 1
    16'b11111101_11000010 : OUT <= 1;  //253 / 194 = 1
    16'b11111101_11000011 : OUT <= 1;  //253 / 195 = 1
    16'b11111101_11000100 : OUT <= 1;  //253 / 196 = 1
    16'b11111101_11000101 : OUT <= 1;  //253 / 197 = 1
    16'b11111101_11000110 : OUT <= 1;  //253 / 198 = 1
    16'b11111101_11000111 : OUT <= 1;  //253 / 199 = 1
    16'b11111101_11001000 : OUT <= 1;  //253 / 200 = 1
    16'b11111101_11001001 : OUT <= 1;  //253 / 201 = 1
    16'b11111101_11001010 : OUT <= 1;  //253 / 202 = 1
    16'b11111101_11001011 : OUT <= 1;  //253 / 203 = 1
    16'b11111101_11001100 : OUT <= 1;  //253 / 204 = 1
    16'b11111101_11001101 : OUT <= 1;  //253 / 205 = 1
    16'b11111101_11001110 : OUT <= 1;  //253 / 206 = 1
    16'b11111101_11001111 : OUT <= 1;  //253 / 207 = 1
    16'b11111101_11010000 : OUT <= 1;  //253 / 208 = 1
    16'b11111101_11010001 : OUT <= 1;  //253 / 209 = 1
    16'b11111101_11010010 : OUT <= 1;  //253 / 210 = 1
    16'b11111101_11010011 : OUT <= 1;  //253 / 211 = 1
    16'b11111101_11010100 : OUT <= 1;  //253 / 212 = 1
    16'b11111101_11010101 : OUT <= 1;  //253 / 213 = 1
    16'b11111101_11010110 : OUT <= 1;  //253 / 214 = 1
    16'b11111101_11010111 : OUT <= 1;  //253 / 215 = 1
    16'b11111101_11011000 : OUT <= 1;  //253 / 216 = 1
    16'b11111101_11011001 : OUT <= 1;  //253 / 217 = 1
    16'b11111101_11011010 : OUT <= 1;  //253 / 218 = 1
    16'b11111101_11011011 : OUT <= 1;  //253 / 219 = 1
    16'b11111101_11011100 : OUT <= 1;  //253 / 220 = 1
    16'b11111101_11011101 : OUT <= 1;  //253 / 221 = 1
    16'b11111101_11011110 : OUT <= 1;  //253 / 222 = 1
    16'b11111101_11011111 : OUT <= 1;  //253 / 223 = 1
    16'b11111101_11100000 : OUT <= 1;  //253 / 224 = 1
    16'b11111101_11100001 : OUT <= 1;  //253 / 225 = 1
    16'b11111101_11100010 : OUT <= 1;  //253 / 226 = 1
    16'b11111101_11100011 : OUT <= 1;  //253 / 227 = 1
    16'b11111101_11100100 : OUT <= 1;  //253 / 228 = 1
    16'b11111101_11100101 : OUT <= 1;  //253 / 229 = 1
    16'b11111101_11100110 : OUT <= 1;  //253 / 230 = 1
    16'b11111101_11100111 : OUT <= 1;  //253 / 231 = 1
    16'b11111101_11101000 : OUT <= 1;  //253 / 232 = 1
    16'b11111101_11101001 : OUT <= 1;  //253 / 233 = 1
    16'b11111101_11101010 : OUT <= 1;  //253 / 234 = 1
    16'b11111101_11101011 : OUT <= 1;  //253 / 235 = 1
    16'b11111101_11101100 : OUT <= 1;  //253 / 236 = 1
    16'b11111101_11101101 : OUT <= 1;  //253 / 237 = 1
    16'b11111101_11101110 : OUT <= 1;  //253 / 238 = 1
    16'b11111101_11101111 : OUT <= 1;  //253 / 239 = 1
    16'b11111101_11110000 : OUT <= 1;  //253 / 240 = 1
    16'b11111101_11110001 : OUT <= 1;  //253 / 241 = 1
    16'b11111101_11110010 : OUT <= 1;  //253 / 242 = 1
    16'b11111101_11110011 : OUT <= 1;  //253 / 243 = 1
    16'b11111101_11110100 : OUT <= 1;  //253 / 244 = 1
    16'b11111101_11110101 : OUT <= 1;  //253 / 245 = 1
    16'b11111101_11110110 : OUT <= 1;  //253 / 246 = 1
    16'b11111101_11110111 : OUT <= 1;  //253 / 247 = 1
    16'b11111101_11111000 : OUT <= 1;  //253 / 248 = 1
    16'b11111101_11111001 : OUT <= 1;  //253 / 249 = 1
    16'b11111101_11111010 : OUT <= 1;  //253 / 250 = 1
    16'b11111101_11111011 : OUT <= 1;  //253 / 251 = 1
    16'b11111101_11111100 : OUT <= 1;  //253 / 252 = 1
    16'b11111101_11111101 : OUT <= 1;  //253 / 253 = 1
    16'b11111101_11111110 : OUT <= 0;  //253 / 254 = 0
    16'b11111101_11111111 : OUT <= 0;  //253 / 255 = 0
    16'b11111110_00000000 : OUT <= 0;  //254 / 0 = 0
    16'b11111110_00000001 : OUT <= 254;  //254 / 1 = 254
    16'b11111110_00000010 : OUT <= 127;  //254 / 2 = 127
    16'b11111110_00000011 : OUT <= 84;  //254 / 3 = 84
    16'b11111110_00000100 : OUT <= 63;  //254 / 4 = 63
    16'b11111110_00000101 : OUT <= 50;  //254 / 5 = 50
    16'b11111110_00000110 : OUT <= 42;  //254 / 6 = 42
    16'b11111110_00000111 : OUT <= 36;  //254 / 7 = 36
    16'b11111110_00001000 : OUT <= 31;  //254 / 8 = 31
    16'b11111110_00001001 : OUT <= 28;  //254 / 9 = 28
    16'b11111110_00001010 : OUT <= 25;  //254 / 10 = 25
    16'b11111110_00001011 : OUT <= 23;  //254 / 11 = 23
    16'b11111110_00001100 : OUT <= 21;  //254 / 12 = 21
    16'b11111110_00001101 : OUT <= 19;  //254 / 13 = 19
    16'b11111110_00001110 : OUT <= 18;  //254 / 14 = 18
    16'b11111110_00001111 : OUT <= 16;  //254 / 15 = 16
    16'b11111110_00010000 : OUT <= 15;  //254 / 16 = 15
    16'b11111110_00010001 : OUT <= 14;  //254 / 17 = 14
    16'b11111110_00010010 : OUT <= 14;  //254 / 18 = 14
    16'b11111110_00010011 : OUT <= 13;  //254 / 19 = 13
    16'b11111110_00010100 : OUT <= 12;  //254 / 20 = 12
    16'b11111110_00010101 : OUT <= 12;  //254 / 21 = 12
    16'b11111110_00010110 : OUT <= 11;  //254 / 22 = 11
    16'b11111110_00010111 : OUT <= 11;  //254 / 23 = 11
    16'b11111110_00011000 : OUT <= 10;  //254 / 24 = 10
    16'b11111110_00011001 : OUT <= 10;  //254 / 25 = 10
    16'b11111110_00011010 : OUT <= 9;  //254 / 26 = 9
    16'b11111110_00011011 : OUT <= 9;  //254 / 27 = 9
    16'b11111110_00011100 : OUT <= 9;  //254 / 28 = 9
    16'b11111110_00011101 : OUT <= 8;  //254 / 29 = 8
    16'b11111110_00011110 : OUT <= 8;  //254 / 30 = 8
    16'b11111110_00011111 : OUT <= 8;  //254 / 31 = 8
    16'b11111110_00100000 : OUT <= 7;  //254 / 32 = 7
    16'b11111110_00100001 : OUT <= 7;  //254 / 33 = 7
    16'b11111110_00100010 : OUT <= 7;  //254 / 34 = 7
    16'b11111110_00100011 : OUT <= 7;  //254 / 35 = 7
    16'b11111110_00100100 : OUT <= 7;  //254 / 36 = 7
    16'b11111110_00100101 : OUT <= 6;  //254 / 37 = 6
    16'b11111110_00100110 : OUT <= 6;  //254 / 38 = 6
    16'b11111110_00100111 : OUT <= 6;  //254 / 39 = 6
    16'b11111110_00101000 : OUT <= 6;  //254 / 40 = 6
    16'b11111110_00101001 : OUT <= 6;  //254 / 41 = 6
    16'b11111110_00101010 : OUT <= 6;  //254 / 42 = 6
    16'b11111110_00101011 : OUT <= 5;  //254 / 43 = 5
    16'b11111110_00101100 : OUT <= 5;  //254 / 44 = 5
    16'b11111110_00101101 : OUT <= 5;  //254 / 45 = 5
    16'b11111110_00101110 : OUT <= 5;  //254 / 46 = 5
    16'b11111110_00101111 : OUT <= 5;  //254 / 47 = 5
    16'b11111110_00110000 : OUT <= 5;  //254 / 48 = 5
    16'b11111110_00110001 : OUT <= 5;  //254 / 49 = 5
    16'b11111110_00110010 : OUT <= 5;  //254 / 50 = 5
    16'b11111110_00110011 : OUT <= 4;  //254 / 51 = 4
    16'b11111110_00110100 : OUT <= 4;  //254 / 52 = 4
    16'b11111110_00110101 : OUT <= 4;  //254 / 53 = 4
    16'b11111110_00110110 : OUT <= 4;  //254 / 54 = 4
    16'b11111110_00110111 : OUT <= 4;  //254 / 55 = 4
    16'b11111110_00111000 : OUT <= 4;  //254 / 56 = 4
    16'b11111110_00111001 : OUT <= 4;  //254 / 57 = 4
    16'b11111110_00111010 : OUT <= 4;  //254 / 58 = 4
    16'b11111110_00111011 : OUT <= 4;  //254 / 59 = 4
    16'b11111110_00111100 : OUT <= 4;  //254 / 60 = 4
    16'b11111110_00111101 : OUT <= 4;  //254 / 61 = 4
    16'b11111110_00111110 : OUT <= 4;  //254 / 62 = 4
    16'b11111110_00111111 : OUT <= 4;  //254 / 63 = 4
    16'b11111110_01000000 : OUT <= 3;  //254 / 64 = 3
    16'b11111110_01000001 : OUT <= 3;  //254 / 65 = 3
    16'b11111110_01000010 : OUT <= 3;  //254 / 66 = 3
    16'b11111110_01000011 : OUT <= 3;  //254 / 67 = 3
    16'b11111110_01000100 : OUT <= 3;  //254 / 68 = 3
    16'b11111110_01000101 : OUT <= 3;  //254 / 69 = 3
    16'b11111110_01000110 : OUT <= 3;  //254 / 70 = 3
    16'b11111110_01000111 : OUT <= 3;  //254 / 71 = 3
    16'b11111110_01001000 : OUT <= 3;  //254 / 72 = 3
    16'b11111110_01001001 : OUT <= 3;  //254 / 73 = 3
    16'b11111110_01001010 : OUT <= 3;  //254 / 74 = 3
    16'b11111110_01001011 : OUT <= 3;  //254 / 75 = 3
    16'b11111110_01001100 : OUT <= 3;  //254 / 76 = 3
    16'b11111110_01001101 : OUT <= 3;  //254 / 77 = 3
    16'b11111110_01001110 : OUT <= 3;  //254 / 78 = 3
    16'b11111110_01001111 : OUT <= 3;  //254 / 79 = 3
    16'b11111110_01010000 : OUT <= 3;  //254 / 80 = 3
    16'b11111110_01010001 : OUT <= 3;  //254 / 81 = 3
    16'b11111110_01010010 : OUT <= 3;  //254 / 82 = 3
    16'b11111110_01010011 : OUT <= 3;  //254 / 83 = 3
    16'b11111110_01010100 : OUT <= 3;  //254 / 84 = 3
    16'b11111110_01010101 : OUT <= 2;  //254 / 85 = 2
    16'b11111110_01010110 : OUT <= 2;  //254 / 86 = 2
    16'b11111110_01010111 : OUT <= 2;  //254 / 87 = 2
    16'b11111110_01011000 : OUT <= 2;  //254 / 88 = 2
    16'b11111110_01011001 : OUT <= 2;  //254 / 89 = 2
    16'b11111110_01011010 : OUT <= 2;  //254 / 90 = 2
    16'b11111110_01011011 : OUT <= 2;  //254 / 91 = 2
    16'b11111110_01011100 : OUT <= 2;  //254 / 92 = 2
    16'b11111110_01011101 : OUT <= 2;  //254 / 93 = 2
    16'b11111110_01011110 : OUT <= 2;  //254 / 94 = 2
    16'b11111110_01011111 : OUT <= 2;  //254 / 95 = 2
    16'b11111110_01100000 : OUT <= 2;  //254 / 96 = 2
    16'b11111110_01100001 : OUT <= 2;  //254 / 97 = 2
    16'b11111110_01100010 : OUT <= 2;  //254 / 98 = 2
    16'b11111110_01100011 : OUT <= 2;  //254 / 99 = 2
    16'b11111110_01100100 : OUT <= 2;  //254 / 100 = 2
    16'b11111110_01100101 : OUT <= 2;  //254 / 101 = 2
    16'b11111110_01100110 : OUT <= 2;  //254 / 102 = 2
    16'b11111110_01100111 : OUT <= 2;  //254 / 103 = 2
    16'b11111110_01101000 : OUT <= 2;  //254 / 104 = 2
    16'b11111110_01101001 : OUT <= 2;  //254 / 105 = 2
    16'b11111110_01101010 : OUT <= 2;  //254 / 106 = 2
    16'b11111110_01101011 : OUT <= 2;  //254 / 107 = 2
    16'b11111110_01101100 : OUT <= 2;  //254 / 108 = 2
    16'b11111110_01101101 : OUT <= 2;  //254 / 109 = 2
    16'b11111110_01101110 : OUT <= 2;  //254 / 110 = 2
    16'b11111110_01101111 : OUT <= 2;  //254 / 111 = 2
    16'b11111110_01110000 : OUT <= 2;  //254 / 112 = 2
    16'b11111110_01110001 : OUT <= 2;  //254 / 113 = 2
    16'b11111110_01110010 : OUT <= 2;  //254 / 114 = 2
    16'b11111110_01110011 : OUT <= 2;  //254 / 115 = 2
    16'b11111110_01110100 : OUT <= 2;  //254 / 116 = 2
    16'b11111110_01110101 : OUT <= 2;  //254 / 117 = 2
    16'b11111110_01110110 : OUT <= 2;  //254 / 118 = 2
    16'b11111110_01110111 : OUT <= 2;  //254 / 119 = 2
    16'b11111110_01111000 : OUT <= 2;  //254 / 120 = 2
    16'b11111110_01111001 : OUT <= 2;  //254 / 121 = 2
    16'b11111110_01111010 : OUT <= 2;  //254 / 122 = 2
    16'b11111110_01111011 : OUT <= 2;  //254 / 123 = 2
    16'b11111110_01111100 : OUT <= 2;  //254 / 124 = 2
    16'b11111110_01111101 : OUT <= 2;  //254 / 125 = 2
    16'b11111110_01111110 : OUT <= 2;  //254 / 126 = 2
    16'b11111110_01111111 : OUT <= 2;  //254 / 127 = 2
    16'b11111110_10000000 : OUT <= 1;  //254 / 128 = 1
    16'b11111110_10000001 : OUT <= 1;  //254 / 129 = 1
    16'b11111110_10000010 : OUT <= 1;  //254 / 130 = 1
    16'b11111110_10000011 : OUT <= 1;  //254 / 131 = 1
    16'b11111110_10000100 : OUT <= 1;  //254 / 132 = 1
    16'b11111110_10000101 : OUT <= 1;  //254 / 133 = 1
    16'b11111110_10000110 : OUT <= 1;  //254 / 134 = 1
    16'b11111110_10000111 : OUT <= 1;  //254 / 135 = 1
    16'b11111110_10001000 : OUT <= 1;  //254 / 136 = 1
    16'b11111110_10001001 : OUT <= 1;  //254 / 137 = 1
    16'b11111110_10001010 : OUT <= 1;  //254 / 138 = 1
    16'b11111110_10001011 : OUT <= 1;  //254 / 139 = 1
    16'b11111110_10001100 : OUT <= 1;  //254 / 140 = 1
    16'b11111110_10001101 : OUT <= 1;  //254 / 141 = 1
    16'b11111110_10001110 : OUT <= 1;  //254 / 142 = 1
    16'b11111110_10001111 : OUT <= 1;  //254 / 143 = 1
    16'b11111110_10010000 : OUT <= 1;  //254 / 144 = 1
    16'b11111110_10010001 : OUT <= 1;  //254 / 145 = 1
    16'b11111110_10010010 : OUT <= 1;  //254 / 146 = 1
    16'b11111110_10010011 : OUT <= 1;  //254 / 147 = 1
    16'b11111110_10010100 : OUT <= 1;  //254 / 148 = 1
    16'b11111110_10010101 : OUT <= 1;  //254 / 149 = 1
    16'b11111110_10010110 : OUT <= 1;  //254 / 150 = 1
    16'b11111110_10010111 : OUT <= 1;  //254 / 151 = 1
    16'b11111110_10011000 : OUT <= 1;  //254 / 152 = 1
    16'b11111110_10011001 : OUT <= 1;  //254 / 153 = 1
    16'b11111110_10011010 : OUT <= 1;  //254 / 154 = 1
    16'b11111110_10011011 : OUT <= 1;  //254 / 155 = 1
    16'b11111110_10011100 : OUT <= 1;  //254 / 156 = 1
    16'b11111110_10011101 : OUT <= 1;  //254 / 157 = 1
    16'b11111110_10011110 : OUT <= 1;  //254 / 158 = 1
    16'b11111110_10011111 : OUT <= 1;  //254 / 159 = 1
    16'b11111110_10100000 : OUT <= 1;  //254 / 160 = 1
    16'b11111110_10100001 : OUT <= 1;  //254 / 161 = 1
    16'b11111110_10100010 : OUT <= 1;  //254 / 162 = 1
    16'b11111110_10100011 : OUT <= 1;  //254 / 163 = 1
    16'b11111110_10100100 : OUT <= 1;  //254 / 164 = 1
    16'b11111110_10100101 : OUT <= 1;  //254 / 165 = 1
    16'b11111110_10100110 : OUT <= 1;  //254 / 166 = 1
    16'b11111110_10100111 : OUT <= 1;  //254 / 167 = 1
    16'b11111110_10101000 : OUT <= 1;  //254 / 168 = 1
    16'b11111110_10101001 : OUT <= 1;  //254 / 169 = 1
    16'b11111110_10101010 : OUT <= 1;  //254 / 170 = 1
    16'b11111110_10101011 : OUT <= 1;  //254 / 171 = 1
    16'b11111110_10101100 : OUT <= 1;  //254 / 172 = 1
    16'b11111110_10101101 : OUT <= 1;  //254 / 173 = 1
    16'b11111110_10101110 : OUT <= 1;  //254 / 174 = 1
    16'b11111110_10101111 : OUT <= 1;  //254 / 175 = 1
    16'b11111110_10110000 : OUT <= 1;  //254 / 176 = 1
    16'b11111110_10110001 : OUT <= 1;  //254 / 177 = 1
    16'b11111110_10110010 : OUT <= 1;  //254 / 178 = 1
    16'b11111110_10110011 : OUT <= 1;  //254 / 179 = 1
    16'b11111110_10110100 : OUT <= 1;  //254 / 180 = 1
    16'b11111110_10110101 : OUT <= 1;  //254 / 181 = 1
    16'b11111110_10110110 : OUT <= 1;  //254 / 182 = 1
    16'b11111110_10110111 : OUT <= 1;  //254 / 183 = 1
    16'b11111110_10111000 : OUT <= 1;  //254 / 184 = 1
    16'b11111110_10111001 : OUT <= 1;  //254 / 185 = 1
    16'b11111110_10111010 : OUT <= 1;  //254 / 186 = 1
    16'b11111110_10111011 : OUT <= 1;  //254 / 187 = 1
    16'b11111110_10111100 : OUT <= 1;  //254 / 188 = 1
    16'b11111110_10111101 : OUT <= 1;  //254 / 189 = 1
    16'b11111110_10111110 : OUT <= 1;  //254 / 190 = 1
    16'b11111110_10111111 : OUT <= 1;  //254 / 191 = 1
    16'b11111110_11000000 : OUT <= 1;  //254 / 192 = 1
    16'b11111110_11000001 : OUT <= 1;  //254 / 193 = 1
    16'b11111110_11000010 : OUT <= 1;  //254 / 194 = 1
    16'b11111110_11000011 : OUT <= 1;  //254 / 195 = 1
    16'b11111110_11000100 : OUT <= 1;  //254 / 196 = 1
    16'b11111110_11000101 : OUT <= 1;  //254 / 197 = 1
    16'b11111110_11000110 : OUT <= 1;  //254 / 198 = 1
    16'b11111110_11000111 : OUT <= 1;  //254 / 199 = 1
    16'b11111110_11001000 : OUT <= 1;  //254 / 200 = 1
    16'b11111110_11001001 : OUT <= 1;  //254 / 201 = 1
    16'b11111110_11001010 : OUT <= 1;  //254 / 202 = 1
    16'b11111110_11001011 : OUT <= 1;  //254 / 203 = 1
    16'b11111110_11001100 : OUT <= 1;  //254 / 204 = 1
    16'b11111110_11001101 : OUT <= 1;  //254 / 205 = 1
    16'b11111110_11001110 : OUT <= 1;  //254 / 206 = 1
    16'b11111110_11001111 : OUT <= 1;  //254 / 207 = 1
    16'b11111110_11010000 : OUT <= 1;  //254 / 208 = 1
    16'b11111110_11010001 : OUT <= 1;  //254 / 209 = 1
    16'b11111110_11010010 : OUT <= 1;  //254 / 210 = 1
    16'b11111110_11010011 : OUT <= 1;  //254 / 211 = 1
    16'b11111110_11010100 : OUT <= 1;  //254 / 212 = 1
    16'b11111110_11010101 : OUT <= 1;  //254 / 213 = 1
    16'b11111110_11010110 : OUT <= 1;  //254 / 214 = 1
    16'b11111110_11010111 : OUT <= 1;  //254 / 215 = 1
    16'b11111110_11011000 : OUT <= 1;  //254 / 216 = 1
    16'b11111110_11011001 : OUT <= 1;  //254 / 217 = 1
    16'b11111110_11011010 : OUT <= 1;  //254 / 218 = 1
    16'b11111110_11011011 : OUT <= 1;  //254 / 219 = 1
    16'b11111110_11011100 : OUT <= 1;  //254 / 220 = 1
    16'b11111110_11011101 : OUT <= 1;  //254 / 221 = 1
    16'b11111110_11011110 : OUT <= 1;  //254 / 222 = 1
    16'b11111110_11011111 : OUT <= 1;  //254 / 223 = 1
    16'b11111110_11100000 : OUT <= 1;  //254 / 224 = 1
    16'b11111110_11100001 : OUT <= 1;  //254 / 225 = 1
    16'b11111110_11100010 : OUT <= 1;  //254 / 226 = 1
    16'b11111110_11100011 : OUT <= 1;  //254 / 227 = 1
    16'b11111110_11100100 : OUT <= 1;  //254 / 228 = 1
    16'b11111110_11100101 : OUT <= 1;  //254 / 229 = 1
    16'b11111110_11100110 : OUT <= 1;  //254 / 230 = 1
    16'b11111110_11100111 : OUT <= 1;  //254 / 231 = 1
    16'b11111110_11101000 : OUT <= 1;  //254 / 232 = 1
    16'b11111110_11101001 : OUT <= 1;  //254 / 233 = 1
    16'b11111110_11101010 : OUT <= 1;  //254 / 234 = 1
    16'b11111110_11101011 : OUT <= 1;  //254 / 235 = 1
    16'b11111110_11101100 : OUT <= 1;  //254 / 236 = 1
    16'b11111110_11101101 : OUT <= 1;  //254 / 237 = 1
    16'b11111110_11101110 : OUT <= 1;  //254 / 238 = 1
    16'b11111110_11101111 : OUT <= 1;  //254 / 239 = 1
    16'b11111110_11110000 : OUT <= 1;  //254 / 240 = 1
    16'b11111110_11110001 : OUT <= 1;  //254 / 241 = 1
    16'b11111110_11110010 : OUT <= 1;  //254 / 242 = 1
    16'b11111110_11110011 : OUT <= 1;  //254 / 243 = 1
    16'b11111110_11110100 : OUT <= 1;  //254 / 244 = 1
    16'b11111110_11110101 : OUT <= 1;  //254 / 245 = 1
    16'b11111110_11110110 : OUT <= 1;  //254 / 246 = 1
    16'b11111110_11110111 : OUT <= 1;  //254 / 247 = 1
    16'b11111110_11111000 : OUT <= 1;  //254 / 248 = 1
    16'b11111110_11111001 : OUT <= 1;  //254 / 249 = 1
    16'b11111110_11111010 : OUT <= 1;  //254 / 250 = 1
    16'b11111110_11111011 : OUT <= 1;  //254 / 251 = 1
    16'b11111110_11111100 : OUT <= 1;  //254 / 252 = 1
    16'b11111110_11111101 : OUT <= 1;  //254 / 253 = 1
    16'b11111110_11111110 : OUT <= 1;  //254 / 254 = 1
    16'b11111110_11111111 : OUT <= 0;  //254 / 255 = 0
    16'b11111111_00000000 : OUT <= 0;  //255 / 0 = 0
    16'b11111111_00000001 : OUT <= 255;  //255 / 1 = 255
    16'b11111111_00000010 : OUT <= 127;  //255 / 2 = 127
    16'b11111111_00000011 : OUT <= 85;  //255 / 3 = 85
    16'b11111111_00000100 : OUT <= 63;  //255 / 4 = 63
    16'b11111111_00000101 : OUT <= 51;  //255 / 5 = 51
    16'b11111111_00000110 : OUT <= 42;  //255 / 6 = 42
    16'b11111111_00000111 : OUT <= 36;  //255 / 7 = 36
    16'b11111111_00001000 : OUT <= 31;  //255 / 8 = 31
    16'b11111111_00001001 : OUT <= 28;  //255 / 9 = 28
    16'b11111111_00001010 : OUT <= 25;  //255 / 10 = 25
    16'b11111111_00001011 : OUT <= 23;  //255 / 11 = 23
    16'b11111111_00001100 : OUT <= 21;  //255 / 12 = 21
    16'b11111111_00001101 : OUT <= 19;  //255 / 13 = 19
    16'b11111111_00001110 : OUT <= 18;  //255 / 14 = 18
    16'b11111111_00001111 : OUT <= 17;  //255 / 15 = 17
    16'b11111111_00010000 : OUT <= 15;  //255 / 16 = 15
    16'b11111111_00010001 : OUT <= 15;  //255 / 17 = 15
    16'b11111111_00010010 : OUT <= 14;  //255 / 18 = 14
    16'b11111111_00010011 : OUT <= 13;  //255 / 19 = 13
    16'b11111111_00010100 : OUT <= 12;  //255 / 20 = 12
    16'b11111111_00010101 : OUT <= 12;  //255 / 21 = 12
    16'b11111111_00010110 : OUT <= 11;  //255 / 22 = 11
    16'b11111111_00010111 : OUT <= 11;  //255 / 23 = 11
    16'b11111111_00011000 : OUT <= 10;  //255 / 24 = 10
    16'b11111111_00011001 : OUT <= 10;  //255 / 25 = 10
    16'b11111111_00011010 : OUT <= 9;  //255 / 26 = 9
    16'b11111111_00011011 : OUT <= 9;  //255 / 27 = 9
    16'b11111111_00011100 : OUT <= 9;  //255 / 28 = 9
    16'b11111111_00011101 : OUT <= 8;  //255 / 29 = 8
    16'b11111111_00011110 : OUT <= 8;  //255 / 30 = 8
    16'b11111111_00011111 : OUT <= 8;  //255 / 31 = 8
    16'b11111111_00100000 : OUT <= 7;  //255 / 32 = 7
    16'b11111111_00100001 : OUT <= 7;  //255 / 33 = 7
    16'b11111111_00100010 : OUT <= 7;  //255 / 34 = 7
    16'b11111111_00100011 : OUT <= 7;  //255 / 35 = 7
    16'b11111111_00100100 : OUT <= 7;  //255 / 36 = 7
    16'b11111111_00100101 : OUT <= 6;  //255 / 37 = 6
    16'b11111111_00100110 : OUT <= 6;  //255 / 38 = 6
    16'b11111111_00100111 : OUT <= 6;  //255 / 39 = 6
    16'b11111111_00101000 : OUT <= 6;  //255 / 40 = 6
    16'b11111111_00101001 : OUT <= 6;  //255 / 41 = 6
    16'b11111111_00101010 : OUT <= 6;  //255 / 42 = 6
    16'b11111111_00101011 : OUT <= 5;  //255 / 43 = 5
    16'b11111111_00101100 : OUT <= 5;  //255 / 44 = 5
    16'b11111111_00101101 : OUT <= 5;  //255 / 45 = 5
    16'b11111111_00101110 : OUT <= 5;  //255 / 46 = 5
    16'b11111111_00101111 : OUT <= 5;  //255 / 47 = 5
    16'b11111111_00110000 : OUT <= 5;  //255 / 48 = 5
    16'b11111111_00110001 : OUT <= 5;  //255 / 49 = 5
    16'b11111111_00110010 : OUT <= 5;  //255 / 50 = 5
    16'b11111111_00110011 : OUT <= 5;  //255 / 51 = 5
    16'b11111111_00110100 : OUT <= 4;  //255 / 52 = 4
    16'b11111111_00110101 : OUT <= 4;  //255 / 53 = 4
    16'b11111111_00110110 : OUT <= 4;  //255 / 54 = 4
    16'b11111111_00110111 : OUT <= 4;  //255 / 55 = 4
    16'b11111111_00111000 : OUT <= 4;  //255 / 56 = 4
    16'b11111111_00111001 : OUT <= 4;  //255 / 57 = 4
    16'b11111111_00111010 : OUT <= 4;  //255 / 58 = 4
    16'b11111111_00111011 : OUT <= 4;  //255 / 59 = 4
    16'b11111111_00111100 : OUT <= 4;  //255 / 60 = 4
    16'b11111111_00111101 : OUT <= 4;  //255 / 61 = 4
    16'b11111111_00111110 : OUT <= 4;  //255 / 62 = 4
    16'b11111111_00111111 : OUT <= 4;  //255 / 63 = 4
    16'b11111111_01000000 : OUT <= 3;  //255 / 64 = 3
    16'b11111111_01000001 : OUT <= 3;  //255 / 65 = 3
    16'b11111111_01000010 : OUT <= 3;  //255 / 66 = 3
    16'b11111111_01000011 : OUT <= 3;  //255 / 67 = 3
    16'b11111111_01000100 : OUT <= 3;  //255 / 68 = 3
    16'b11111111_01000101 : OUT <= 3;  //255 / 69 = 3
    16'b11111111_01000110 : OUT <= 3;  //255 / 70 = 3
    16'b11111111_01000111 : OUT <= 3;  //255 / 71 = 3
    16'b11111111_01001000 : OUT <= 3;  //255 / 72 = 3
    16'b11111111_01001001 : OUT <= 3;  //255 / 73 = 3
    16'b11111111_01001010 : OUT <= 3;  //255 / 74 = 3
    16'b11111111_01001011 : OUT <= 3;  //255 / 75 = 3
    16'b11111111_01001100 : OUT <= 3;  //255 / 76 = 3
    16'b11111111_01001101 : OUT <= 3;  //255 / 77 = 3
    16'b11111111_01001110 : OUT <= 3;  //255 / 78 = 3
    16'b11111111_01001111 : OUT <= 3;  //255 / 79 = 3
    16'b11111111_01010000 : OUT <= 3;  //255 / 80 = 3
    16'b11111111_01010001 : OUT <= 3;  //255 / 81 = 3
    16'b11111111_01010010 : OUT <= 3;  //255 / 82 = 3
    16'b11111111_01010011 : OUT <= 3;  //255 / 83 = 3
    16'b11111111_01010100 : OUT <= 3;  //255 / 84 = 3
    16'b11111111_01010101 : OUT <= 3;  //255 / 85 = 3
    16'b11111111_01010110 : OUT <= 2;  //255 / 86 = 2
    16'b11111111_01010111 : OUT <= 2;  //255 / 87 = 2
    16'b11111111_01011000 : OUT <= 2;  //255 / 88 = 2
    16'b11111111_01011001 : OUT <= 2;  //255 / 89 = 2
    16'b11111111_01011010 : OUT <= 2;  //255 / 90 = 2
    16'b11111111_01011011 : OUT <= 2;  //255 / 91 = 2
    16'b11111111_01011100 : OUT <= 2;  //255 / 92 = 2
    16'b11111111_01011101 : OUT <= 2;  //255 / 93 = 2
    16'b11111111_01011110 : OUT <= 2;  //255 / 94 = 2
    16'b11111111_01011111 : OUT <= 2;  //255 / 95 = 2
    16'b11111111_01100000 : OUT <= 2;  //255 / 96 = 2
    16'b11111111_01100001 : OUT <= 2;  //255 / 97 = 2
    16'b11111111_01100010 : OUT <= 2;  //255 / 98 = 2
    16'b11111111_01100011 : OUT <= 2;  //255 / 99 = 2
    16'b11111111_01100100 : OUT <= 2;  //255 / 100 = 2
    16'b11111111_01100101 : OUT <= 2;  //255 / 101 = 2
    16'b11111111_01100110 : OUT <= 2;  //255 / 102 = 2
    16'b11111111_01100111 : OUT <= 2;  //255 / 103 = 2
    16'b11111111_01101000 : OUT <= 2;  //255 / 104 = 2
    16'b11111111_01101001 : OUT <= 2;  //255 / 105 = 2
    16'b11111111_01101010 : OUT <= 2;  //255 / 106 = 2
    16'b11111111_01101011 : OUT <= 2;  //255 / 107 = 2
    16'b11111111_01101100 : OUT <= 2;  //255 / 108 = 2
    16'b11111111_01101101 : OUT <= 2;  //255 / 109 = 2
    16'b11111111_01101110 : OUT <= 2;  //255 / 110 = 2
    16'b11111111_01101111 : OUT <= 2;  //255 / 111 = 2
    16'b11111111_01110000 : OUT <= 2;  //255 / 112 = 2
    16'b11111111_01110001 : OUT <= 2;  //255 / 113 = 2
    16'b11111111_01110010 : OUT <= 2;  //255 / 114 = 2
    16'b11111111_01110011 : OUT <= 2;  //255 / 115 = 2
    16'b11111111_01110100 : OUT <= 2;  //255 / 116 = 2
    16'b11111111_01110101 : OUT <= 2;  //255 / 117 = 2
    16'b11111111_01110110 : OUT <= 2;  //255 / 118 = 2
    16'b11111111_01110111 : OUT <= 2;  //255 / 119 = 2
    16'b11111111_01111000 : OUT <= 2;  //255 / 120 = 2
    16'b11111111_01111001 : OUT <= 2;  //255 / 121 = 2
    16'b11111111_01111010 : OUT <= 2;  //255 / 122 = 2
    16'b11111111_01111011 : OUT <= 2;  //255 / 123 = 2
    16'b11111111_01111100 : OUT <= 2;  //255 / 124 = 2
    16'b11111111_01111101 : OUT <= 2;  //255 / 125 = 2
    16'b11111111_01111110 : OUT <= 2;  //255 / 126 = 2
    16'b11111111_01111111 : OUT <= 2;  //255 / 127 = 2
    16'b11111111_10000000 : OUT <= 1;  //255 / 128 = 1
    16'b11111111_10000001 : OUT <= 1;  //255 / 129 = 1
    16'b11111111_10000010 : OUT <= 1;  //255 / 130 = 1
    16'b11111111_10000011 : OUT <= 1;  //255 / 131 = 1
    16'b11111111_10000100 : OUT <= 1;  //255 / 132 = 1
    16'b11111111_10000101 : OUT <= 1;  //255 / 133 = 1
    16'b11111111_10000110 : OUT <= 1;  //255 / 134 = 1
    16'b11111111_10000111 : OUT <= 1;  //255 / 135 = 1
    16'b11111111_10001000 : OUT <= 1;  //255 / 136 = 1
    16'b11111111_10001001 : OUT <= 1;  //255 / 137 = 1
    16'b11111111_10001010 : OUT <= 1;  //255 / 138 = 1
    16'b11111111_10001011 : OUT <= 1;  //255 / 139 = 1
    16'b11111111_10001100 : OUT <= 1;  //255 / 140 = 1
    16'b11111111_10001101 : OUT <= 1;  //255 / 141 = 1
    16'b11111111_10001110 : OUT <= 1;  //255 / 142 = 1
    16'b11111111_10001111 : OUT <= 1;  //255 / 143 = 1
    16'b11111111_10010000 : OUT <= 1;  //255 / 144 = 1
    16'b11111111_10010001 : OUT <= 1;  //255 / 145 = 1
    16'b11111111_10010010 : OUT <= 1;  //255 / 146 = 1
    16'b11111111_10010011 : OUT <= 1;  //255 / 147 = 1
    16'b11111111_10010100 : OUT <= 1;  //255 / 148 = 1
    16'b11111111_10010101 : OUT <= 1;  //255 / 149 = 1
    16'b11111111_10010110 : OUT <= 1;  //255 / 150 = 1
    16'b11111111_10010111 : OUT <= 1;  //255 / 151 = 1
    16'b11111111_10011000 : OUT <= 1;  //255 / 152 = 1
    16'b11111111_10011001 : OUT <= 1;  //255 / 153 = 1
    16'b11111111_10011010 : OUT <= 1;  //255 / 154 = 1
    16'b11111111_10011011 : OUT <= 1;  //255 / 155 = 1
    16'b11111111_10011100 : OUT <= 1;  //255 / 156 = 1
    16'b11111111_10011101 : OUT <= 1;  //255 / 157 = 1
    16'b11111111_10011110 : OUT <= 1;  //255 / 158 = 1
    16'b11111111_10011111 : OUT <= 1;  //255 / 159 = 1
    16'b11111111_10100000 : OUT <= 1;  //255 / 160 = 1
    16'b11111111_10100001 : OUT <= 1;  //255 / 161 = 1
    16'b11111111_10100010 : OUT <= 1;  //255 / 162 = 1
    16'b11111111_10100011 : OUT <= 1;  //255 / 163 = 1
    16'b11111111_10100100 : OUT <= 1;  //255 / 164 = 1
    16'b11111111_10100101 : OUT <= 1;  //255 / 165 = 1
    16'b11111111_10100110 : OUT <= 1;  //255 / 166 = 1
    16'b11111111_10100111 : OUT <= 1;  //255 / 167 = 1
    16'b11111111_10101000 : OUT <= 1;  //255 / 168 = 1
    16'b11111111_10101001 : OUT <= 1;  //255 / 169 = 1
    16'b11111111_10101010 : OUT <= 1;  //255 / 170 = 1
    16'b11111111_10101011 : OUT <= 1;  //255 / 171 = 1
    16'b11111111_10101100 : OUT <= 1;  //255 / 172 = 1
    16'b11111111_10101101 : OUT <= 1;  //255 / 173 = 1
    16'b11111111_10101110 : OUT <= 1;  //255 / 174 = 1
    16'b11111111_10101111 : OUT <= 1;  //255 / 175 = 1
    16'b11111111_10110000 : OUT <= 1;  //255 / 176 = 1
    16'b11111111_10110001 : OUT <= 1;  //255 / 177 = 1
    16'b11111111_10110010 : OUT <= 1;  //255 / 178 = 1
    16'b11111111_10110011 : OUT <= 1;  //255 / 179 = 1
    16'b11111111_10110100 : OUT <= 1;  //255 / 180 = 1
    16'b11111111_10110101 : OUT <= 1;  //255 / 181 = 1
    16'b11111111_10110110 : OUT <= 1;  //255 / 182 = 1
    16'b11111111_10110111 : OUT <= 1;  //255 / 183 = 1
    16'b11111111_10111000 : OUT <= 1;  //255 / 184 = 1
    16'b11111111_10111001 : OUT <= 1;  //255 / 185 = 1
    16'b11111111_10111010 : OUT <= 1;  //255 / 186 = 1
    16'b11111111_10111011 : OUT <= 1;  //255 / 187 = 1
    16'b11111111_10111100 : OUT <= 1;  //255 / 188 = 1
    16'b11111111_10111101 : OUT <= 1;  //255 / 189 = 1
    16'b11111111_10111110 : OUT <= 1;  //255 / 190 = 1
    16'b11111111_10111111 : OUT <= 1;  //255 / 191 = 1
    16'b11111111_11000000 : OUT <= 1;  //255 / 192 = 1
    16'b11111111_11000001 : OUT <= 1;  //255 / 193 = 1
    16'b11111111_11000010 : OUT <= 1;  //255 / 194 = 1
    16'b11111111_11000011 : OUT <= 1;  //255 / 195 = 1
    16'b11111111_11000100 : OUT <= 1;  //255 / 196 = 1
    16'b11111111_11000101 : OUT <= 1;  //255 / 197 = 1
    16'b11111111_11000110 : OUT <= 1;  //255 / 198 = 1
    16'b11111111_11000111 : OUT <= 1;  //255 / 199 = 1
    16'b11111111_11001000 : OUT <= 1;  //255 / 200 = 1
    16'b11111111_11001001 : OUT <= 1;  //255 / 201 = 1
    16'b11111111_11001010 : OUT <= 1;  //255 / 202 = 1
    16'b11111111_11001011 : OUT <= 1;  //255 / 203 = 1
    16'b11111111_11001100 : OUT <= 1;  //255 / 204 = 1
    16'b11111111_11001101 : OUT <= 1;  //255 / 205 = 1
    16'b11111111_11001110 : OUT <= 1;  //255 / 206 = 1
    16'b11111111_11001111 : OUT <= 1;  //255 / 207 = 1
    16'b11111111_11010000 : OUT <= 1;  //255 / 208 = 1
    16'b11111111_11010001 : OUT <= 1;  //255 / 209 = 1
    16'b11111111_11010010 : OUT <= 1;  //255 / 210 = 1
    16'b11111111_11010011 : OUT <= 1;  //255 / 211 = 1
    16'b11111111_11010100 : OUT <= 1;  //255 / 212 = 1
    16'b11111111_11010101 : OUT <= 1;  //255 / 213 = 1
    16'b11111111_11010110 : OUT <= 1;  //255 / 214 = 1
    16'b11111111_11010111 : OUT <= 1;  //255 / 215 = 1
    16'b11111111_11011000 : OUT <= 1;  //255 / 216 = 1
    16'b11111111_11011001 : OUT <= 1;  //255 / 217 = 1
    16'b11111111_11011010 : OUT <= 1;  //255 / 218 = 1
    16'b11111111_11011011 : OUT <= 1;  //255 / 219 = 1
    16'b11111111_11011100 : OUT <= 1;  //255 / 220 = 1
    16'b11111111_11011101 : OUT <= 1;  //255 / 221 = 1
    16'b11111111_11011110 : OUT <= 1;  //255 / 222 = 1
    16'b11111111_11011111 : OUT <= 1;  //255 / 223 = 1
    16'b11111111_11100000 : OUT <= 1;  //255 / 224 = 1
    16'b11111111_11100001 : OUT <= 1;  //255 / 225 = 1
    16'b11111111_11100010 : OUT <= 1;  //255 / 226 = 1
    16'b11111111_11100011 : OUT <= 1;  //255 / 227 = 1
    16'b11111111_11100100 : OUT <= 1;  //255 / 228 = 1
    16'b11111111_11100101 : OUT <= 1;  //255 / 229 = 1
    16'b11111111_11100110 : OUT <= 1;  //255 / 230 = 1
    16'b11111111_11100111 : OUT <= 1;  //255 / 231 = 1
    16'b11111111_11101000 : OUT <= 1;  //255 / 232 = 1
    16'b11111111_11101001 : OUT <= 1;  //255 / 233 = 1
    16'b11111111_11101010 : OUT <= 1;  //255 / 234 = 1
    16'b11111111_11101011 : OUT <= 1;  //255 / 235 = 1
    16'b11111111_11101100 : OUT <= 1;  //255 / 236 = 1
    16'b11111111_11101101 : OUT <= 1;  //255 / 237 = 1
    16'b11111111_11101110 : OUT <= 1;  //255 / 238 = 1
    16'b11111111_11101111 : OUT <= 1;  //255 / 239 = 1
    16'b11111111_11110000 : OUT <= 1;  //255 / 240 = 1
    16'b11111111_11110001 : OUT <= 1;  //255 / 241 = 1
    16'b11111111_11110010 : OUT <= 1;  //255 / 242 = 1
    16'b11111111_11110011 : OUT <= 1;  //255 / 243 = 1
    16'b11111111_11110100 : OUT <= 1;  //255 / 244 = 1
    16'b11111111_11110101 : OUT <= 1;  //255 / 245 = 1
    16'b11111111_11110110 : OUT <= 1;  //255 / 246 = 1
    16'b11111111_11110111 : OUT <= 1;  //255 / 247 = 1
    16'b11111111_11111000 : OUT <= 1;  //255 / 248 = 1
    16'b11111111_11111001 : OUT <= 1;  //255 / 249 = 1
    16'b11111111_11111010 : OUT <= 1;  //255 / 250 = 1
    16'b11111111_11111011 : OUT <= 1;  //255 / 251 = 1
    16'b11111111_11111100 : OUT <= 1;  //255 / 252 = 1
    16'b11111111_11111101 : OUT <= 1;  //255 / 253 = 1
    16'b11111111_11111110 : OUT <= 1;  //255 / 254 = 1
    16'b11111111_11111111 : OUT <= 1;  //255 / 255 = 1
endcase

endmodule
