`timescale 1ns / 1ps

/*
	Name: Hai Dang Hoang
	Email: danghai@pdx.edu
	Module multiplication 8x8 bit (A^2)
*/

module multi_8x8(clk, operand, OUT);
input clk;
input [7:0] operand;
output reg [15:0] OUT;

always @(posedge clk)
case ({operand,operand}) 

16'b00000000_00000000 : OUT <= 0; //0 * 0 = 0
16'b00000001_00000001 : OUT <= 1; //1 * 1 = 1
16'b00000010_00000010 : OUT <= 4; //2 * 2 = 4
16'b00000011_00000011 : OUT <= 9; //3 * 3 = 9
16'b00000100_00000100 : OUT <= 16; //4 * 4 = 16
16'b00000101_00000101 : OUT <= 25; //5 * 5 = 25
16'b00000110_00000110 : OUT <= 36; //6 * 6 = 36
16'b00000111_00000111 : OUT <= 49; //7 * 7 = 49
16'b00001000_00001000 : OUT <= 64; //8 * 8 = 64
16'b00001001_00001001 : OUT <= 81; //9 * 9 = 81
16'b00001010_00001010 : OUT <= 100; //10 * 10 = 100
16'b00001011_00001011 : OUT <= 121; //11 * 11 = 121
16'b00001100_00001100 : OUT <= 144; //12 * 12 = 144
16'b00001101_00001101 : OUT <= 169; //13 * 13 = 169
16'b00001110_00001110 : OUT <= 196; //14 * 14 = 196
16'b00001111_00001111 : OUT <= 225; //15 * 15 = 225
16'b00010000_00010000 : OUT <= 256; //16 * 16 = 256
16'b00010001_00010001 : OUT <= 289; //17 * 17 = 289
16'b00010010_00010010 : OUT <= 324; //18 * 18 = 324
16'b00010011_00010011 : OUT <= 361; //19 * 19 = 361
16'b00010100_00010100 : OUT <= 400; //20 * 20 = 400
16'b00010101_00010101 : OUT <= 441; //21 * 21 = 441
16'b00010110_00010110 : OUT <= 484; //22 * 22 = 484
16'b00010111_00010111 : OUT <= 529; //23 * 23 = 529
16'b00011000_00011000 : OUT <= 576; //24 * 24 = 576
16'b00011001_00011001 : OUT <= 625; //25 * 25 = 625
16'b00011010_00011010 : OUT <= 676; //26 * 26 = 676
16'b00011011_00011011 : OUT <= 729; //27 * 27 = 729
16'b00011100_00011100 : OUT <= 784; //28 * 28 = 784
16'b00011101_00011101 : OUT <= 841; //29 * 29 = 841
16'b00011110_00011110 : OUT <= 900; //30 * 30 = 900
16'b00011111_00011111 : OUT <= 961; //31 * 31 = 961
16'b00100000_00100000 : OUT <= 1024; //32 * 32 = 1024
16'b00100001_00100001 : OUT <= 1089; //33 * 33 = 1089
16'b00100010_00100010 : OUT <= 1156; //34 * 34 = 1156
16'b00100011_00100011 : OUT <= 1225; //35 * 35 = 1225
16'b00100100_00100100 : OUT <= 1296; //36 * 36 = 1296
16'b00100101_00100101 : OUT <= 1369; //37 * 37 = 1369
16'b00100110_00100110 : OUT <= 1444; //38 * 38 = 1444
16'b00100111_00100111 : OUT <= 1521; //39 * 39 = 1521
16'b00101000_00101000 : OUT <= 1600; //40 * 40 = 1600
16'b00101001_00101001 : OUT <= 1681; //41 * 41 = 1681
16'b00101010_00101010 : OUT <= 1764; //42 * 42 = 1764
16'b00101011_00101011 : OUT <= 1849; //43 * 43 = 1849
16'b00101100_00101100 : OUT <= 1936; //44 * 44 = 1936
16'b00101101_00101101 : OUT <= 2025; //45 * 45 = 2025
16'b00101110_00101110 : OUT <= 2116; //46 * 46 = 2116
16'b00101111_00101111 : OUT <= 2209; //47 * 47 = 2209
16'b00110000_00110000 : OUT <= 2304; //48 * 48 = 2304
16'b00110001_00110001 : OUT <= 2401; //49 * 49 = 2401
16'b00110010_00110010 : OUT <= 2500; //50 * 50 = 2500
16'b00110011_00110011 : OUT <= 2601; //51 * 51 = 2601
16'b00110100_00110100 : OUT <= 2704; //52 * 52 = 2704
16'b00110101_00110101 : OUT <= 2809; //53 * 53 = 2809
16'b00110110_00110110 : OUT <= 2916; //54 * 54 = 2916
16'b00110111_00110111 : OUT <= 3025; //55 * 55 = 3025
16'b00111000_00111000 : OUT <= 3136; //56 * 56 = 3136
16'b00111001_00111001 : OUT <= 3249; //57 * 57 = 3249
16'b00111010_00111010 : OUT <= 3364; //58 * 58 = 3364
16'b00111011_00111011 : OUT <= 3481; //59 * 59 = 3481
16'b00111100_00111100 : OUT <= 3600; //60 * 60 = 3600
16'b00111101_00111101 : OUT <= 3721; //61 * 61 = 3721
16'b00111110_00111110 : OUT <= 3844; //62 * 62 = 3844
16'b00111111_00111111 : OUT <= 3969; //63 * 63 = 3969
16'b01000000_01000000 : OUT <= 4096; //64 * 64 = 4096
16'b01000001_01000001 : OUT <= 4225; //65 * 65 = 4225
16'b01000010_01000010 : OUT <= 4356; //66 * 66 = 4356
16'b01000011_01000011 : OUT <= 4489; //67 * 67 = 4489
16'b01000100_01000100 : OUT <= 4624; //68 * 68 = 4624
16'b01000101_01000101 : OUT <= 4761; //69 * 69 = 4761
16'b01000110_01000110 : OUT <= 4900; //70 * 70 = 4900
16'b01000111_01000111 : OUT <= 5041; //71 * 71 = 5041
16'b01001000_01001000 : OUT <= 5184; //72 * 72 = 5184
16'b01001001_01001001 : OUT <= 5329; //73 * 73 = 5329
16'b01001010_01001010 : OUT <= 5476; //74 * 74 = 5476
16'b01001011_01001011 : OUT <= 5625; //75 * 75 = 5625
16'b01001100_01001100 : OUT <= 5776; //76 * 76 = 5776
16'b01001101_01001101 : OUT <= 5929; //77 * 77 = 5929
16'b01001110_01001110 : OUT <= 6084; //78 * 78 = 6084
16'b01001111_01001111 : OUT <= 6241; //79 * 79 = 6241
16'b01010000_01010000 : OUT <= 6400; //80 * 80 = 6400
16'b01010001_01010001 : OUT <= 6561; //81 * 81 = 6561
16'b01010010_01010010 : OUT <= 6724; //82 * 82 = 6724
16'b01010011_01010011 : OUT <= 6889; //83 * 83 = 6889
16'b01010100_01010100 : OUT <= 7056; //84 * 84 = 7056
16'b01010101_01010101 : OUT <= 7225; //85 * 85 = 7225
16'b01010110_01010110 : OUT <= 7396; //86 * 86 = 7396
16'b01010111_01010111 : OUT <= 7569; //87 * 87 = 7569
16'b01011000_01011000 : OUT <= 7744; //88 * 88 = 7744
16'b01011001_01011001 : OUT <= 7921; //89 * 89 = 7921
16'b01011010_01011010 : OUT <= 8100; //90 * 90 = 8100
16'b01011011_01011011 : OUT <= 8281; //91 * 91 = 8281
16'b01011100_01011100 : OUT <= 8464; //92 * 92 = 8464
16'b01011101_01011101 : OUT <= 8649; //93 * 93 = 8649
16'b01011110_01011110 : OUT <= 8836; //94 * 94 = 8836
16'b01011111_01011111 : OUT <= 9025; //95 * 95 = 9025
16'b01100000_01100000 : OUT <= 9216; //96 * 96 = 9216
16'b01100001_01100001 : OUT <= 9409; //97 * 97 = 9409
16'b01100010_01100010 : OUT <= 9604; //98 * 98 = 9604
16'b01100011_01100011 : OUT <= 9801; //99 * 99 = 9801
16'b01100100_01100100 : OUT <= 10000; //100 * 100 = 10000
16'b01100101_01100101 : OUT <= 10201; //101 * 101 = 10201
16'b01100110_01100110 : OUT <= 10404; //102 * 102 = 10404
16'b01100111_01100111 : OUT <= 10609; //103 * 103 = 10609
16'b01101000_01101000 : OUT <= 10816; //104 * 104 = 10816
16'b01101001_01101001 : OUT <= 11025; //105 * 105 = 11025
16'b01101010_01101010 : OUT <= 11236; //106 * 106 = 11236
16'b01101011_01101011 : OUT <= 11449; //107 * 107 = 11449
16'b01101100_01101100 : OUT <= 11664; //108 * 108 = 11664
16'b01101101_01101101 : OUT <= 11881; //109 * 109 = 11881
16'b01101110_01101110 : OUT <= 12100; //110 * 110 = 12100
16'b01101111_01101111 : OUT <= 12321; //111 * 111 = 12321
16'b01110000_01110000 : OUT <= 12544; //112 * 112 = 12544
16'b01110001_01110001 : OUT <= 12769; //113 * 113 = 12769
16'b01110010_01110010 : OUT <= 12996; //114 * 114 = 12996
16'b01110011_01110011 : OUT <= 13225; //115 * 115 = 13225
16'b01110100_01110100 : OUT <= 13456; //116 * 116 = 13456
16'b01110101_01110101 : OUT <= 13689; //117 * 117 = 13689
16'b01110110_01110110 : OUT <= 13924; //118 * 118 = 13924
16'b01110111_01110111 : OUT <= 14161; //119 * 119 = 14161
16'b01111000_01111000 : OUT <= 14400; //120 * 120 = 14400
16'b01111001_01111001 : OUT <= 14641; //121 * 121 = 14641
16'b01111010_01111010 : OUT <= 14884; //122 * 122 = 14884
16'b01111011_01111011 : OUT <= 15129; //123 * 123 = 15129
16'b01111100_01111100 : OUT <= 15376; //124 * 124 = 15376
16'b01111101_01111101 : OUT <= 15625; //125 * 125 = 15625
16'b01111110_01111110 : OUT <= 15876; //126 * 126 = 15876
16'b01111111_01111111 : OUT <= 16129; //127 * 127 = 16129
16'b10000000_10000000 : OUT <= 16384; //128 * 128 = 16384
16'b10000001_10000001 : OUT <= 16641; //129 * 129 = 16641
16'b10000010_10000010 : OUT <= 16900; //130 * 130 = 16900
16'b10000011_10000011 : OUT <= 17161; //131 * 131 = 17161
16'b10000100_10000100 : OUT <= 17424; //132 * 132 = 17424
16'b10000101_10000101 : OUT <= 17689; //133 * 133 = 17689
16'b10000110_10000110 : OUT <= 17956; //134 * 134 = 17956
16'b10000111_10000111 : OUT <= 18225; //135 * 135 = 18225
16'b10001000_10001000 : OUT <= 18496; //136 * 136 = 18496
16'b10001001_10001001 : OUT <= 18769; //137 * 137 = 18769
16'b10001010_10001010 : OUT <= 19044; //138 * 138 = 19044
16'b10001011_10001011 : OUT <= 19321; //139 * 139 = 19321
16'b10001100_10001100 : OUT <= 19600; //140 * 140 = 19600
16'b10001101_10001101 : OUT <= 19881; //141 * 141 = 19881
16'b10001110_10001110 : OUT <= 20164; //142 * 142 = 20164
16'b10001111_10001111 : OUT <= 20449; //143 * 143 = 20449
16'b10010000_10010000 : OUT <= 20736; //144 * 144 = 20736
16'b10010001_10010001 : OUT <= 21025; //145 * 145 = 21025
16'b10010010_10010010 : OUT <= 21316; //146 * 146 = 21316
16'b10010011_10010011 : OUT <= 21609; //147 * 147 = 21609
16'b10010100_10010100 : OUT <= 21904; //148 * 148 = 21904
16'b10010101_10010101 : OUT <= 22201; //149 * 149 = 22201
16'b10010110_10010110 : OUT <= 22500; //150 * 150 = 22500
16'b10010111_10010111 : OUT <= 22801; //151 * 151 = 22801
16'b10011000_10011000 : OUT <= 23104; //152 * 152 = 23104
16'b10011001_10011001 : OUT <= 23409; //153 * 153 = 23409
16'b10011010_10011010 : OUT <= 23716; //154 * 154 = 23716
16'b10011011_10011011 : OUT <= 24025; //155 * 155 = 24025
16'b10011100_10011100 : OUT <= 24336; //156 * 156 = 24336
16'b10011101_10011101 : OUT <= 24649; //157 * 157 = 24649
16'b10011110_10011110 : OUT <= 24964; //158 * 158 = 24964
16'b10011111_10011111 : OUT <= 25281; //159 * 159 = 25281
16'b10100000_10100000 : OUT <= 25600; //160 * 160 = 25600
16'b10100001_10100001 : OUT <= 25921; //161 * 161 = 25921
16'b10100010_10100010 : OUT <= 26244; //162 * 162 = 26244
16'b10100011_10100011 : OUT <= 26569; //163 * 163 = 26569
16'b10100100_10100100 : OUT <= 26896; //164 * 164 = 26896
16'b10100101_10100101 : OUT <= 27225; //165 * 165 = 27225
16'b10100110_10100110 : OUT <= 27556; //166 * 166 = 27556
16'b10100111_10100111 : OUT <= 27889; //167 * 167 = 27889
16'b10101000_10101000 : OUT <= 28224; //168 * 168 = 28224
16'b10101001_10101001 : OUT <= 28561; //169 * 169 = 28561
16'b10101010_10101010 : OUT <= 28900; //170 * 170 = 28900
16'b10101011_10101011 : OUT <= 29241; //171 * 171 = 29241
16'b10101100_10101100 : OUT <= 29584; //172 * 172 = 29584
16'b10101101_10101101 : OUT <= 29929; //173 * 173 = 29929
16'b10101110_10101110 : OUT <= 30276; //174 * 174 = 30276
16'b10101111_10101111 : OUT <= 30625; //175 * 175 = 30625
16'b10110000_10110000 : OUT <= 30976; //176 * 176 = 30976
16'b10110001_10110001 : OUT <= 31329; //177 * 177 = 31329
16'b10110010_10110010 : OUT <= 31684; //178 * 178 = 31684
16'b10110011_10110011 : OUT <= 32041; //179 * 179 = 32041
16'b10110100_10110100 : OUT <= 32400; //180 * 180 = 32400
16'b10110101_10110101 : OUT <= 32761; //181 * 181 = 32761
16'b10110110_10110110 : OUT <= 33124; //182 * 182 = 33124
16'b10110111_10110111 : OUT <= 33489; //183 * 183 = 33489
16'b10111000_10111000 : OUT <= 33856; //184 * 184 = 33856
16'b10111001_10111001 : OUT <= 34225; //185 * 185 = 34225
16'b10111010_10111010 : OUT <= 34596; //186 * 186 = 34596
16'b10111011_10111011 : OUT <= 34969; //187 * 187 = 34969
16'b10111100_10111100 : OUT <= 35344; //188 * 188 = 35344
16'b10111101_10111101 : OUT <= 35721; //189 * 189 = 35721
16'b10111110_10111110 : OUT <= 36100; //190 * 190 = 36100
16'b10111111_10111111 : OUT <= 36481; //191 * 191 = 36481
16'b11000000_11000000 : OUT <= 36864; //192 * 192 = 36864
16'b11000001_11000001 : OUT <= 37249; //193 * 193 = 37249
16'b11000010_11000010 : OUT <= 37636; //194 * 194 = 37636
16'b11000011_11000011 : OUT <= 38025; //195 * 195 = 38025
16'b11000100_11000100 : OUT <= 38416; //196 * 196 = 38416
16'b11000101_11000101 : OUT <= 38809; //197 * 197 = 38809
16'b11000110_11000110 : OUT <= 39204; //198 * 198 = 39204
16'b11000111_11000111 : OUT <= 39601; //199 * 199 = 39601
16'b11001000_11001000 : OUT <= 40000; //200 * 200 = 40000
16'b11001001_11001001 : OUT <= 40401; //201 * 201 = 40401
16'b11001010_11001010 : OUT <= 40804; //202 * 202 = 40804
16'b11001011_11001011 : OUT <= 41209; //203 * 203 = 41209
16'b11001100_11001100 : OUT <= 41616; //204 * 204 = 41616
16'b11001101_11001101 : OUT <= 42025; //205 * 205 = 42025
16'b11001110_11001110 : OUT <= 42436; //206 * 206 = 42436
16'b11001111_11001111 : OUT <= 42849; //207 * 207 = 42849
16'b11010000_11010000 : OUT <= 43264; //208 * 208 = 43264
16'b11010001_11010001 : OUT <= 43681; //209 * 209 = 43681
16'b11010010_11010010 : OUT <= 44100; //210 * 210 = 44100
16'b11010011_11010011 : OUT <= 44521; //211 * 211 = 44521
16'b11010100_11010100 : OUT <= 44944; //212 * 212 = 44944
16'b11010101_11010101 : OUT <= 45369; //213 * 213 = 45369
16'b11010110_11010110 : OUT <= 45796; //214 * 214 = 45796
16'b11010111_11010111 : OUT <= 46225; //215 * 215 = 46225
16'b11011000_11011000 : OUT <= 46656; //216 * 216 = 46656
16'b11011001_11011001 : OUT <= 47089; //217 * 217 = 47089
16'b11011010_11011010 : OUT <= 47524; //218 * 218 = 47524
16'b11011011_11011011 : OUT <= 47961; //219 * 219 = 47961
16'b11011100_11011100 : OUT <= 48400; //220 * 220 = 48400
16'b11011101_11011101 : OUT <= 48841; //221 * 221 = 48841
16'b11011110_11011110 : OUT <= 49284; //222 * 222 = 49284
16'b11011111_11011111 : OUT <= 49729; //223 * 223 = 49729
16'b11100000_11100000 : OUT <= 50176; //224 * 224 = 50176
16'b11100001_11100001 : OUT <= 50625; //225 * 225 = 50625
16'b11100010_11100010 : OUT <= 51076; //226 * 226 = 51076
16'b11100011_11100011 : OUT <= 51529; //227 * 227 = 51529
16'b11100100_11100100 : OUT <= 51984; //228 * 228 = 51984
16'b11100101_11100101 : OUT <= 52441; //229 * 229 = 52441
16'b11100110_11100110 : OUT <= 52900; //230 * 230 = 52900
16'b11100111_11100111 : OUT <= 53361; //231 * 231 = 53361
16'b11101000_11101000 : OUT <= 53824; //232 * 232 = 53824
16'b11101001_11101001 : OUT <= 54289; //233 * 233 = 54289
16'b11101010_11101010 : OUT <= 54756; //234 * 234 = 54756
16'b11101011_11101011 : OUT <= 55225; //235 * 235 = 55225
16'b11101100_11101100 : OUT <= 55696; //236 * 236 = 55696
16'b11101101_11101101 : OUT <= 56169; //237 * 237 = 56169
16'b11101110_11101110 : OUT <= 56644; //238 * 238 = 56644
16'b11101111_11101111 : OUT <= 57121; //239 * 239 = 57121
16'b11110000_11110000 : OUT <= 57600; //240 * 240 = 57600
16'b11110001_11110001 : OUT <= 58081; //241 * 241 = 58081
16'b11110010_11110010 : OUT <= 58564; //242 * 242 = 58564
16'b11110011_11110011 : OUT <= 59049; //243 * 243 = 59049
16'b11110100_11110100 : OUT <= 59536; //244 * 244 = 59536
16'b11110101_11110101 : OUT <= 60025; //245 * 245 = 60025
16'b11110110_11110110 : OUT <= 60516; //246 * 246 = 60516
16'b11110111_11110111 : OUT <= 61009; //247 * 247 = 61009
16'b11111000_11111000 : OUT <= 61504; //248 * 248 = 61504
16'b11111001_11111001 : OUT <= 62001; //249 * 249 = 62001
16'b11111010_11111010 : OUT <= 62500; //250 * 250 = 62500
16'b11111011_11111011 : OUT <= 63001; //251 * 251 = 63001
16'b11111100_11111100 : OUT <= 63504; //252 * 252 = 63504
16'b11111101_11111101 : OUT <= 64009; //253 * 253 = 64009
16'b11111110_11111110 : OUT <= 64516; //254 * 254 = 64516
16'b11111111_11111111 : OUT <= 65025; //255 * 255 = 65025

default: OUT <= 0;
endcase
endmodule
